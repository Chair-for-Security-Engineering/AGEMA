module Reg1(x, y);
 input [133:0] x;
 output [132:0] y;

  assign y[0] = x[133];
  assign y[5] = x[0];
  assign y[6] = x[11];
  assign y[7] = x[22];
  assign y[8] = x[33];
  assign y[9] = x[44];
  assign y[10] = x[55];
  assign y[11] = x[60];
  assign y[12] = x[61];
  assign y[13] = x[62];
  assign y[14] = x[63];
  assign y[15] = x[1];
  assign y[16] = x[2];
  assign y[17] = x[3];
  assign y[18] = x[4];
  assign y[19] = x[5];
  assign y[20] = x[6];
  assign y[21] = x[7];
  assign y[22] = x[8];
  assign y[23] = x[9];
  assign y[24] = x[10];
  assign y[25] = x[12];
  assign y[26] = x[13];
  assign y[27] = x[14];
  assign y[28] = x[15];
  assign y[29] = x[16];
  assign y[30] = x[17];
  assign y[31] = x[18];
  assign y[32] = x[19];
  assign y[33] = x[20];
  assign y[34] = x[21];
  assign y[35] = x[23];
  assign y[36] = x[24];
  assign y[37] = x[25];
  assign y[38] = x[26];
  assign y[39] = x[27];
  assign y[40] = x[28];
  assign y[41] = x[29];
  assign y[42] = x[30];
  assign y[43] = x[31];
  assign y[44] = x[32];
  assign y[45] = x[34];
  assign y[46] = x[35];
  assign y[47] = x[36];
  assign y[48] = x[37];
  assign y[49] = x[38];
  assign y[50] = x[39];
  assign y[51] = x[40];
  assign y[52] = x[41];
  assign y[53] = x[42];
  assign y[54] = x[43];
  assign y[55] = x[45];
  assign y[56] = x[46];
  assign y[57] = x[47];
  assign y[58] = x[48];
  assign y[59] = x[49];
  assign y[60] = x[50];
  assign y[61] = x[51];
  assign y[62] = x[52];
  assign y[63] = x[53];
  assign y[64] = x[54];
  assign y[65] = x[56];
  assign y[66] = x[57];
  assign y[67] = x[58];
  assign y[68] = x[59];
  register_stage #(.WIDTH(68)) inst_0(.clk(x[128]), .D({x[129],x[130],x[131],x[132],x[64],x[75],x[86],x[97],x[108],x[119],x[124],x[125],x[126],x[127],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[120],x[121],x[122],x[123]}), .Q({y[1],y[2],y[3],y[4],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132]}));
endmodule

module Reg2(x, y);
 input [266:0] x;
 output [265:0] y;

  assign y[0] = x[265];
  assign y[1] = x[266];
  assign y[10] = x[0];
  assign y[11] = x[1];
  assign y[12] = x[22];
  assign y[13] = x[23];
  assign y[14] = x[44];
  assign y[15] = x[45];
  assign y[16] = x[66];
  assign y[17] = x[67];
  assign y[18] = x[88];
  assign y[19] = x[89];
  assign y[20] = x[110];
  assign y[21] = x[111];
  assign y[22] = x[120];
  assign y[23] = x[121];
  assign y[24] = x[122];
  assign y[25] = x[123];
  assign y[26] = x[124];
  assign y[27] = x[125];
  assign y[28] = x[126];
  assign y[29] = x[127];
  assign y[30] = x[2];
  assign y[31] = x[3];
  assign y[32] = x[4];
  assign y[33] = x[5];
  assign y[34] = x[6];
  assign y[35] = x[7];
  assign y[36] = x[8];
  assign y[37] = x[9];
  assign y[38] = x[10];
  assign y[39] = x[11];
  assign y[40] = x[12];
  assign y[41] = x[13];
  assign y[42] = x[14];
  assign y[43] = x[15];
  assign y[44] = x[16];
  assign y[45] = x[17];
  assign y[46] = x[18];
  assign y[47] = x[19];
  assign y[48] = x[20];
  assign y[49] = x[21];
  assign y[50] = x[24];
  assign y[51] = x[25];
  assign y[52] = x[26];
  assign y[53] = x[27];
  assign y[54] = x[28];
  assign y[55] = x[29];
  assign y[56] = x[30];
  assign y[57] = x[31];
  assign y[58] = x[32];
  assign y[59] = x[33];
  assign y[60] = x[34];
  assign y[61] = x[35];
  assign y[62] = x[36];
  assign y[63] = x[37];
  assign y[64] = x[38];
  assign y[65] = x[39];
  assign y[66] = x[40];
  assign y[67] = x[41];
  assign y[68] = x[42];
  assign y[69] = x[43];
  assign y[70] = x[46];
  assign y[71] = x[47];
  assign y[72] = x[48];
  assign y[73] = x[49];
  assign y[74] = x[50];
  assign y[75] = x[51];
  assign y[76] = x[52];
  assign y[77] = x[53];
  assign y[78] = x[54];
  assign y[79] = x[55];
  assign y[80] = x[56];
  assign y[81] = x[57];
  assign y[82] = x[58];
  assign y[83] = x[59];
  assign y[84] = x[60];
  assign y[85] = x[61];
  assign y[86] = x[62];
  assign y[87] = x[63];
  assign y[88] = x[64];
  assign y[89] = x[65];
  assign y[90] = x[68];
  assign y[91] = x[69];
  assign y[92] = x[70];
  assign y[93] = x[71];
  assign y[94] = x[72];
  assign y[95] = x[73];
  assign y[96] = x[74];
  assign y[97] = x[75];
  assign y[98] = x[76];
  assign y[99] = x[77];
  assign y[100] = x[78];
  assign y[101] = x[79];
  assign y[102] = x[80];
  assign y[103] = x[81];
  assign y[104] = x[82];
  assign y[105] = x[83];
  assign y[106] = x[84];
  assign y[107] = x[85];
  assign y[108] = x[86];
  assign y[109] = x[87];
  assign y[110] = x[90];
  assign y[111] = x[91];
  assign y[112] = x[92];
  assign y[113] = x[93];
  assign y[114] = x[94];
  assign y[115] = x[95];
  assign y[116] = x[96];
  assign y[117] = x[97];
  assign y[118] = x[98];
  assign y[119] = x[99];
  assign y[120] = x[100];
  assign y[121] = x[101];
  assign y[122] = x[102];
  assign y[123] = x[103];
  assign y[124] = x[104];
  assign y[125] = x[105];
  assign y[126] = x[106];
  assign y[127] = x[107];
  assign y[128] = x[108];
  assign y[129] = x[109];
  assign y[130] = x[112];
  assign y[131] = x[113];
  assign y[132] = x[114];
  assign y[133] = x[115];
  assign y[134] = x[116];
  assign y[135] = x[117];
  assign y[136] = x[118];
  assign y[137] = x[119];
  register_stage #(.WIDTH(136)) inst_0(.clk(x[256]), .D({x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[128],x[129],x[150],x[151],x[172],x[173],x[194],x[195],x[216],x[217],x[238],x[239],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247]}), .Q({y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [398:0] x;
 output [265:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[223], x[222]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[224], x[222]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[226], x[225]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[227], x[225]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[229], x[228]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[230], x[228]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[232], x[231]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[233], x[231]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[235], x[234]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[236], x[234]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[238], x[237]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[239], x[237]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[241], x[240]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[242], x[240]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[244], x[243]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[245], x[243]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[247], x[246]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[248], x[246]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[250], x[249]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[251], x[249]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[253], x[252]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[254], x[252]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[256], x[255]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[257], x[255]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[259], x[258]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[260], x[258]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[262], x[261]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[263], x[261]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[265], x[264]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[266], x[264]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[268], x[267]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[269], x[267]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[271], x[270]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[272], x[270]}), .y(y[181]));
  Fx182 Fx182_inst(.x({x[274], x[273]}), .y(y[182]));
  Fx183 Fx183_inst(.x({x[275], x[273]}), .y(y[183]));
  Fx184 Fx184_inst(.x({x[277], x[276]}), .y(y[184]));
  Fx185 Fx185_inst(.x({x[278], x[276]}), .y(y[185]));
  Fx186 Fx186_inst(.x({x[280], x[279]}), .y(y[186]));
  Fx187 Fx187_inst(.x({x[281], x[279]}), .y(y[187]));
  Fx188 Fx188_inst(.x({x[283], x[282]}), .y(y[188]));
  Fx189 Fx189_inst(.x({x[284], x[282]}), .y(y[189]));
  Fx190 Fx190_inst(.x({x[286], x[285]}), .y(y[190]));
  Fx191 Fx191_inst(.x({x[287], x[285]}), .y(y[191]));
  Fx192 Fx192_inst(.x({x[289], x[288]}), .y(y[192]));
  Fx193 Fx193_inst(.x({x[290], x[288]}), .y(y[193]));
  Fx194 Fx194_inst(.x({x[292], x[291]}), .y(y[194]));
  Fx195 Fx195_inst(.x({x[293], x[291]}), .y(y[195]));
  Fx196 Fx196_inst(.x({x[295], x[294]}), .y(y[196]));
  Fx197 Fx197_inst(.x({x[296], x[294]}), .y(y[197]));
  Fx198 Fx198_inst(.x({x[298], x[297]}), .y(y[198]));
  Fx199 Fx199_inst(.x({x[299], x[297]}), .y(y[199]));
  Fx200 Fx200_inst(.x({x[301], x[300]}), .y(y[200]));
  Fx201 Fx201_inst(.x({x[302], x[300]}), .y(y[201]));
  Fx202 Fx202_inst(.x({x[304], x[303]}), .y(y[202]));
  Fx203 Fx203_inst(.x({x[305], x[303]}), .y(y[203]));
  Fx204 Fx204_inst(.x({x[307], x[306]}), .y(y[204]));
  Fx205 Fx205_inst(.x({x[308], x[306]}), .y(y[205]));
  Fx206 Fx206_inst(.x({x[310], x[309]}), .y(y[206]));
  Fx207 Fx207_inst(.x({x[311], x[309]}), .y(y[207]));
  Fx208 Fx208_inst(.x({x[313], x[312]}), .y(y[208]));
  Fx209 Fx209_inst(.x({x[314], x[312]}), .y(y[209]));
  Fx210 Fx210_inst(.x({x[316], x[315]}), .y(y[210]));
  Fx211 Fx211_inst(.x({x[317], x[315]}), .y(y[211]));
  Fx212 Fx212_inst(.x({x[319], x[318]}), .y(y[212]));
  Fx213 Fx213_inst(.x({x[320], x[318]}), .y(y[213]));
  Fx214 Fx214_inst(.x({x[322], x[321]}), .y(y[214]));
  Fx215 Fx215_inst(.x({x[323], x[321]}), .y(y[215]));
  Fx216 Fx216_inst(.x({x[325], x[324]}), .y(y[216]));
  Fx217 Fx217_inst(.x({x[326], x[324]}), .y(y[217]));
  Fx218 Fx218_inst(.x({x[328], x[327]}), .y(y[218]));
  Fx219 Fx219_inst(.x({x[329], x[327]}), .y(y[219]));
  Fx220 Fx220_inst(.x({x[331], x[330]}), .y(y[220]));
  Fx221 Fx221_inst(.x({x[332], x[330]}), .y(y[221]));
  Fx222 Fx222_inst(.x({x[334], x[333]}), .y(y[222]));
  Fx223 Fx223_inst(.x({x[335], x[333]}), .y(y[223]));
  Fx224 Fx224_inst(.x({x[337], x[336]}), .y(y[224]));
  Fx225 Fx225_inst(.x({x[338], x[336]}), .y(y[225]));
  Fx226 Fx226_inst(.x({x[340], x[339]}), .y(y[226]));
  Fx227 Fx227_inst(.x({x[341], x[339]}), .y(y[227]));
  Fx228 Fx228_inst(.x({x[343], x[342]}), .y(y[228]));
  Fx229 Fx229_inst(.x({x[344], x[342]}), .y(y[229]));
  Fx230 Fx230_inst(.x({x[346], x[345]}), .y(y[230]));
  Fx231 Fx231_inst(.x({x[347], x[345]}), .y(y[231]));
  Fx232 Fx232_inst(.x({x[349], x[348]}), .y(y[232]));
  Fx233 Fx233_inst(.x({x[350], x[348]}), .y(y[233]));
  Fx234 Fx234_inst(.x({x[352], x[351]}), .y(y[234]));
  Fx235 Fx235_inst(.x({x[353], x[351]}), .y(y[235]));
  Fx236 Fx236_inst(.x({x[355], x[354]}), .y(y[236]));
  Fx237 Fx237_inst(.x({x[356], x[354]}), .y(y[237]));
  Fx238 Fx238_inst(.x({x[358], x[357]}), .y(y[238]));
  Fx239 Fx239_inst(.x({x[359], x[357]}), .y(y[239]));
  Fx240 Fx240_inst(.x({x[361], x[360]}), .y(y[240]));
  Fx241 Fx241_inst(.x({x[362], x[360]}), .y(y[241]));
  Fx242 Fx242_inst(.x({x[364], x[363]}), .y(y[242]));
  Fx243 Fx243_inst(.x({x[365], x[363]}), .y(y[243]));
  Fx244 Fx244_inst(.x({x[367], x[366]}), .y(y[244]));
  Fx245 Fx245_inst(.x({x[368], x[366]}), .y(y[245]));
  Fx246 Fx246_inst(.x({x[370], x[369]}), .y(y[246]));
  Fx247 Fx247_inst(.x({x[371], x[369]}), .y(y[247]));
  Fx248 Fx248_inst(.x({x[373], x[372]}), .y(y[248]));
  Fx249 Fx249_inst(.x({x[374], x[372]}), .y(y[249]));
  Fx250 Fx250_inst(.x({x[376], x[375]}), .y(y[250]));
  Fx251 Fx251_inst(.x({x[377], x[375]}), .y(y[251]));
  Fx252 Fx252_inst(.x({x[379], x[378]}), .y(y[252]));
  Fx253 Fx253_inst(.x({x[380], x[378]}), .y(y[253]));
  Fx254 Fx254_inst(.x({x[382], x[381]}), .y(y[254]));
  Fx255 Fx255_inst(.x({x[383], x[381]}), .y(y[255]));
  Fx256 Fx256_inst(.x({x[385], x[384]}), .y(y[256]));
  Fx257 Fx257_inst(.x({x[386], x[384]}), .y(y[257]));
  Fx258 Fx258_inst(.x({x[388], x[387]}), .y(y[258]));
  Fx259 Fx259_inst(.x({x[389], x[387]}), .y(y[259]));
  Fx260 Fx260_inst(.x({x[391], x[390]}), .y(y[260]));
  Fx261 Fx261_inst(.x({x[392], x[390]}), .y(y[261]));
  Fx262 Fx262_inst(.x({x[394], x[393]}), .y(y[262]));
  Fx263 Fx263_inst(.x({x[395], x[393]}), .y(y[263]));
  Fx264 Fx264_inst(.x({x[397], x[396]}), .y(y[264]));
  Fx265 Fx265_inst(.x({x[398], x[396]}), .y(y[265]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind66(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind67(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind68(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind69(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind70(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind72(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind73(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind74(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind76(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind77(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind78(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind79(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind80(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind81(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind82(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind83(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind84(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind85(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind86(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind87(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind88(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind89(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind90(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind91(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind92(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind93(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind94(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind95(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind96(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind97(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind98(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind99(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind100(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind101(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind102(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind103(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind104(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind105(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind106(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind107(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind108(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind109(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind110(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind111(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind112(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind113(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind114(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind115(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind116(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind117(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind118(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind119(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind120(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind121(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind122(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind123(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind124(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind125(x, y);
 input [13:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[13];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[8] & x[9]);
  assign t[15] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = t[0] ^ t[1];
endmodule

module R1ind126(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind127(x, y);
 input [10:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[5] & x[6]);
  assign t[12] = (x[8] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[7];
  assign t[9] = t[12] ^ x[10];
  assign y = t[0] ^ t[1];
endmodule

module R1ind128(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = t[16] ^ x[13];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[5] & x[6]);
  assign t[15] = (x[8] & x[9]);
  assign t[16] = (x[11] & x[12]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind129(x, y);
 input [11:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[2] = t[6] ^ x[2];
  assign t[3] = t[7] ^ x[5];
  assign t[4] = t[8] ^ x[8];
  assign t[5] = t[9] ^ x[11];
  assign t[6] = (x[0] & x[1]);
  assign t[7] = (x[3] & x[4]);
  assign t[8] = (x[6] & x[7]);
  assign t[9] = (x[9] & x[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind130(x, y);
 input [97:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[11] & x[12]);
  assign t[101] = (x[14] & x[15]);
  assign t[102] = (x[17] & x[18]);
  assign t[103] = (x[20] & x[21]);
  assign t[104] = (x[25] & x[26]);
  assign t[105] = (x[28] & x[29]);
  assign t[106] = (x[31] & x[32]);
  assign t[107] = (x[34] & x[35]);
  assign t[108] = (x[39] & x[40]);
  assign t[109] = (x[44] & x[45]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[47] & x[48]);
  assign t[111] = (x[50] & x[51]);
  assign t[112] = (x[53] & x[54]);
  assign t[113] = (x[56] & x[57]);
  assign t[114] = (x[59] & x[60]);
  assign t[115] = (x[62] & x[63]);
  assign t[116] = (x[65] & x[66]);
  assign t[117] = (x[68] & x[69]);
  assign t[118] = (x[71] & x[72]);
  assign t[119] = (x[74] & x[75]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[120] = (x[77] & x[78]);
  assign t[121] = (x[80] & x[81]);
  assign t[122] = (x[83] & x[84]);
  assign t[123] = (x[86] & x[87]);
  assign t[124] = (x[89] & x[90]);
  assign t[125] = (x[92] & x[93]);
  assign t[126] = (x[95] & x[96]);
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[70] & t[71]);
  assign t[15] = ~(t[72] & t[73]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[72]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] | t[74];
  assign t[24] = t[16] ? x[24] : x[23];
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = ~(t[35] & t[36]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[75]);
  assign t[31] = ~(t[76]);
  assign t[32] = ~(t[43] | t[30]);
  assign t[33] = ~(t[44] & t[45]);
  assign t[34] = t[46] | t[77];
  assign t[35] = ~(t[47] & t[48]);
  assign t[36] = t[49] | t[78];
  assign t[37] = t[50] ? x[38] : x[37];
  assign t[38] = ~(t[51] & t[52]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[79];
  assign t[41] = t[16] ? x[43] : x[42];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[80]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[58] | t[44]);
  assign t[47] = ~(t[83]);
  assign t[48] = ~(t[84]);
  assign t[49] = ~(t[59] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[21]);
  assign t[51] = ~(t[60] & t[61]);
  assign t[52] = t[62] | t[85];
  assign t[53] = ~(t[86]);
  assign t[54] = ~(t[87]);
  assign t[55] = ~(t[63] | t[53]);
  assign t[56] = ~(t[64] & t[65]);
  assign t[57] = t[66] | t[88];
  assign t[58] = ~(t[89]);
  assign t[59] = ~(t[90]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[92]);
  assign t[62] = ~(t[67] | t[60]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[94]);
  assign t[65] = ~(t[95]);
  assign t[66] = ~(t[68] | t[64]);
  assign t[67] = ~(t[96]);
  assign t[68] = ~(t[97]);
  assign t[69] = t[98] ^ x[2];
  assign t[6] = t[11] ^ t[7];
  assign t[70] = t[99] ^ x[10];
  assign t[71] = t[100] ^ x[13];
  assign t[72] = t[101] ^ x[16];
  assign t[73] = t[102] ^ x[19];
  assign t[74] = t[103] ^ x[22];
  assign t[75] = t[104] ^ x[27];
  assign t[76] = t[105] ^ x[30];
  assign t[77] = t[106] ^ x[33];
  assign t[78] = t[107] ^ x[36];
  assign t[79] = t[108] ^ x[41];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[109] ^ x[46];
  assign t[81] = t[110] ^ x[49];
  assign t[82] = t[111] ^ x[52];
  assign t[83] = t[112] ^ x[55];
  assign t[84] = t[113] ^ x[58];
  assign t[85] = t[114] ^ x[61];
  assign t[86] = t[115] ^ x[64];
  assign t[87] = t[116] ^ x[67];
  assign t[88] = t[117] ^ x[70];
  assign t[89] = t[118] ^ x[73];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[119] ^ x[76];
  assign t[91] = t[120] ^ x[79];
  assign t[92] = t[121] ^ x[82];
  assign t[93] = t[122] ^ x[85];
  assign t[94] = t[123] ^ x[88];
  assign t[95] = t[124] ^ x[91];
  assign t[96] = t[125] ^ x[94];
  assign t[97] = t[126] ^ x[97];
  assign t[98] = (x[0] & x[1]);
  assign t[99] = (x[8] & x[9]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[69];
endmodule

module R1ind131(x, y);
 input [97:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[129] ^ x[88];
  assign t[101] = t[130] ^ x[91];
  assign t[102] = t[131] ^ x[94];
  assign t[103] = t[132] ^ x[97];
  assign t[104] = (x[0] & x[1]);
  assign t[105] = (x[8] & x[9]);
  assign t[106] = (x[11] & x[12]);
  assign t[107] = (x[14] & x[15]);
  assign t[108] = (x[17] & x[18]);
  assign t[109] = (x[20] & x[21]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[25] & x[26]);
  assign t[111] = (x[28] & x[29]);
  assign t[112] = (x[31] & x[32]);
  assign t[113] = (x[34] & x[35]);
  assign t[114] = (x[39] & x[40]);
  assign t[115] = (x[44] & x[45]);
  assign t[116] = (x[47] & x[48]);
  assign t[117] = (x[50] & x[51]);
  assign t[118] = (x[53] & x[54]);
  assign t[119] = (x[56] & x[57]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[120] = (x[59] & x[60]);
  assign t[121] = (x[62] & x[63]);
  assign t[122] = (x[65] & x[66]);
  assign t[123] = (x[68] & x[69]);
  assign t[124] = (x[71] & x[72]);
  assign t[125] = (x[74] & x[75]);
  assign t[126] = (x[77] & x[78]);
  assign t[127] = (x[80] & x[81]);
  assign t[128] = (x[83] & x[84]);
  assign t[129] = (x[86] & x[87]);
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[130] = (x[89] & x[90]);
  assign t[131] = (x[92] & x[93]);
  assign t[132] = (x[95] & x[96]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[76] & t[77]);
  assign t[15] = ~(t[78] & t[79]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[78]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] & t[80]);
  assign t[24] = t[16] ? x[24] : x[23];
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = ~(t[35] & t[36]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[81]);
  assign t[31] = ~(t[82]);
  assign t[32] = ~(t[43] & t[44]);
  assign t[33] = ~(t[45] & t[46]);
  assign t[34] = ~(t[47] & t[83]);
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[50] & t[84]);
  assign t[37] = t[51] ? x[38] : x[37];
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[85]);
  assign t[41] = t[16] ? x[43] : x[42];
  assign t[42] = ~(t[57] & t[58]);
  assign t[43] = ~(t[82] & t[81]);
  assign t[44] = ~(t[86]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[59] & t[60]);
  assign t[48] = ~(t[89]);
  assign t[49] = ~(t[90]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[61] & t[62]);
  assign t[51] = ~(t[21]);
  assign t[52] = ~(t[63] & t[64]);
  assign t[53] = ~(t[65] & t[91]);
  assign t[54] = ~(t[92]);
  assign t[55] = ~(t[93]);
  assign t[56] = ~(t[66] & t[67]);
  assign t[57] = ~(t[68] & t[69]);
  assign t[58] = ~(t[70] & t[94]);
  assign t[59] = ~(t[88] & t[87]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[90] & t[89]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[71] & t[72]);
  assign t[66] = ~(t[93] & t[92]);
  assign t[67] = ~(t[99]);
  assign t[68] = ~(t[100]);
  assign t[69] = ~(t[101]);
  assign t[6] = t[11] ^ t[7];
  assign t[70] = ~(t[73] & t[74]);
  assign t[71] = ~(t[98] & t[97]);
  assign t[72] = ~(t[102]);
  assign t[73] = ~(t[101] & t[100]);
  assign t[74] = ~(t[103]);
  assign t[75] = t[104] ^ x[2];
  assign t[76] = t[105] ^ x[10];
  assign t[77] = t[106] ^ x[13];
  assign t[78] = t[107] ^ x[16];
  assign t[79] = t[108] ^ x[19];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[109] ^ x[22];
  assign t[81] = t[110] ^ x[27];
  assign t[82] = t[111] ^ x[30];
  assign t[83] = t[112] ^ x[33];
  assign t[84] = t[113] ^ x[36];
  assign t[85] = t[114] ^ x[41];
  assign t[86] = t[115] ^ x[46];
  assign t[87] = t[116] ^ x[49];
  assign t[88] = t[117] ^ x[52];
  assign t[89] = t[118] ^ x[55];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[119] ^ x[58];
  assign t[91] = t[120] ^ x[61];
  assign t[92] = t[121] ^ x[64];
  assign t[93] = t[122] ^ x[67];
  assign t[94] = t[123] ^ x[70];
  assign t[95] = t[124] ^ x[73];
  assign t[96] = t[125] ^ x[76];
  assign t[97] = t[126] ^ x[79];
  assign t[98] = t[127] ^ x[82];
  assign t[99] = t[128] ^ x[85];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[75];
endmodule

module R1ind132(x, y);
 input [79:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[53] & x[54]);
  assign t[101] = (x[56] & x[57]);
  assign t[102] = (x[59] & x[60]);
  assign t[103] = (x[62] & x[63]);
  assign t[104] = (x[65] & x[66]);
  assign t[105] = (x[68] & x[69]);
  assign t[106] = (x[71] & x[72]);
  assign t[107] = (x[74] & x[75]);
  assign t[108] = (x[77] & x[78]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[64] & t[65]);
  assign t[15] = ~(t[66] & t[67]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[66]);
  assign t[22] = ~(t[68] & t[30]);
  assign t[23] = ~(t[69] & t[31]);
  assign t[24] = t[16] ? x[27] : x[26];
  assign t[25] = ~(t[32] & t[33]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[70]);
  assign t[31] = ~(t[70] & t[42]);
  assign t[32] = ~(t[71] & t[43]);
  assign t[33] = ~(t[72] & t[44]);
  assign t[34] = ~(t[73] & t[45]);
  assign t[35] = ~(t[74] & t[46]);
  assign t[36] = t[47] ? x[44] : x[43];
  assign t[37] = ~(t[48] & t[49]);
  assign t[38] = ~(t[75] & t[50]);
  assign t[39] = ~(t[76] & t[51]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[16] ? x[52] : x[51];
  assign t[41] = ~(t[52] & t[53]);
  assign t[42] = ~(t[68]);
  assign t[43] = ~(t[77]);
  assign t[44] = ~(t[77] & t[54]);
  assign t[45] = ~(t[78]);
  assign t[46] = ~(t[78] & t[55]);
  assign t[47] = ~(t[21]);
  assign t[48] = ~(t[79] & t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81]);
  assign t[51] = ~(t[81] & t[58]);
  assign t[52] = ~(t[82] & t[59]);
  assign t[53] = ~(t[83] & t[60]);
  assign t[54] = ~(t[71]);
  assign t[55] = ~(t[73]);
  assign t[56] = ~(t[84]);
  assign t[57] = ~(t[84] & t[61]);
  assign t[58] = ~(t[75]);
  assign t[59] = ~(t[85]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[85] & t[62]);
  assign t[61] = ~(t[79]);
  assign t[62] = ~(t[82]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[10];
  assign t[65] = t[88] ^ x[13];
  assign t[66] = t[89] ^ x[16];
  assign t[67] = t[90] ^ x[19];
  assign t[68] = t[91] ^ x[22];
  assign t[69] = t[92] ^ x[25];
  assign t[6] = t[11] ^ t[7];
  assign t[70] = t[93] ^ x[30];
  assign t[71] = t[94] ^ x[33];
  assign t[72] = t[95] ^ x[36];
  assign t[73] = t[96] ^ x[39];
  assign t[74] = t[97] ^ x[42];
  assign t[75] = t[98] ^ x[47];
  assign t[76] = t[99] ^ x[50];
  assign t[77] = t[100] ^ x[55];
  assign t[78] = t[101] ^ x[58];
  assign t[79] = t[102] ^ x[61];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[103] ^ x[64];
  assign t[81] = t[104] ^ x[67];
  assign t[82] = t[105] ^ x[70];
  assign t[83] = t[106] ^ x[73];
  assign t[84] = t[107] ^ x[76];
  assign t[85] = t[108] ^ x[79];
  assign t[86] = (x[0] & x[1]);
  assign t[87] = (x[8] & x[9]);
  assign t[88] = (x[11] & x[12]);
  assign t[89] = (x[14] & x[15]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = (x[17] & x[18]);
  assign t[91] = (x[20] & x[21]);
  assign t[92] = (x[23] & x[24]);
  assign t[93] = (x[28] & x[29]);
  assign t[94] = (x[31] & x[32]);
  assign t[95] = (x[34] & x[35]);
  assign t[96] = (x[37] & x[38]);
  assign t[97] = (x[40] & x[41]);
  assign t[98] = (x[45] & x[46]);
  assign t[99] = (x[48] & x[49]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[63];
endmodule

module R1ind133(x, y);
 input [97:0] x;
 output y;

 wire [201:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[161] | t[162]);
  assign t[101] = ~(t[169]);
  assign t[102] = ~(t[170]);
  assign t[103] = ~(t[124] | t[125]);
  assign t[104] = ~(t[33]);
  assign t[105] = ~(t[84] | t[126]);
  assign t[106] = ~(t[127]);
  assign t[107] = x[4] & t[146];
  assign t[108] = ~(t[148]);
  assign t[109] = ~(x[4] | t[146]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[146] | t[148]);
  assign t[111] = ~(x[4] | t[128]);
  assign t[112] = t[145] ? t[129] : t[83];
  assign t[113] = t[145] ? t[80] : t[130];
  assign t[114] = t[145] ? t[80] : t[81];
  assign t[115] = ~(t[34] | t[131]);
  assign t[116] = ~(t[53] & t[132]);
  assign t[117] = ~(t[122] & t[133]);
  assign t[118] = t[53] | t[134];
  assign t[119] = ~(t[171]);
  assign t[11] = ~(t[16] ^ t[17]);
  assign t[120] = ~(t[166] | t[167]);
  assign t[121] = ~(t[57] | t[135]);
  assign t[122] = t[148] & t[136];
  assign t[123] = ~(t[64]);
  assign t[124] = ~(t[172]);
  assign t[125] = ~(t[169] | t[170]);
  assign t[126] = ~(t[137] & t[64]);
  assign t[127] = ~(t[57] | t[138]);
  assign t[128] = ~(t[146]);
  assign t[129] = ~(x[4] & t[139]);
  assign t[12] = x[4] ? t[19] : t[18];
  assign t[130] = ~(t[109] & t[148]);
  assign t[131] = ~(t[57] | t[140]);
  assign t[132] = ~(t[82] & t[86]);
  assign t[133] = t[109] | t[107];
  assign t[134] = t[145] ? t[82] : t[83];
  assign t[135] = t[145] ? t[82] : t[86];
  assign t[136] = ~(t[53] | t[145]);
  assign t[137] = ~(t[141] | t[90]);
  assign t[138] = t[145] ? t[81] : t[142];
  assign t[139] = ~(t[146] | t[108]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[145] ? t[83] : t[129];
  assign t[141] = ~(t[57] | t[143]);
  assign t[142] = ~(t[107] & t[148]);
  assign t[143] = t[145] ? t[142] : t[81];
  assign t[144] = t[173] ^ x[2];
  assign t[145] = t[174] ^ x[10];
  assign t[146] = t[175] ^ x[13];
  assign t[147] = t[176] ^ x[16];
  assign t[148] = t[177] ^ x[19];
  assign t[149] = t[178] ^ x[22];
  assign t[14] = ~(t[145] & t[146]);
  assign t[150] = t[179] ^ x[25];
  assign t[151] = t[180] ^ x[28];
  assign t[152] = t[181] ^ x[31];
  assign t[153] = t[182] ^ x[36];
  assign t[154] = t[183] ^ x[39];
  assign t[155] = t[184] ^ x[42];
  assign t[156] = t[185] ^ x[45];
  assign t[157] = t[186] ^ x[48];
  assign t[158] = t[187] ^ x[51];
  assign t[159] = t[188] ^ x[54];
  assign t[15] = ~(t[147] & t[148]);
  assign t[160] = t[189] ^ x[57];
  assign t[161] = t[190] ^ x[62];
  assign t[162] = t[191] ^ x[65];
  assign t[163] = t[192] ^ x[68];
  assign t[164] = t[193] ^ x[73];
  assign t[165] = t[194] ^ x[76];
  assign t[166] = t[195] ^ x[79];
  assign t[167] = t[196] ^ x[82];
  assign t[168] = t[197] ^ x[85];
  assign t[169] = t[198] ^ x[88];
  assign t[16] = t[22] ? x[7] : x[6];
  assign t[170] = t[199] ^ x[91];
  assign t[171] = t[200] ^ x[94];
  assign t[172] = t[201] ^ x[97];
  assign t[173] = (x[0] & x[1]);
  assign t[174] = (x[8] & x[9]);
  assign t[175] = (x[11] & x[12]);
  assign t[176] = (x[14] & x[15]);
  assign t[177] = (x[17] & x[18]);
  assign t[178] = (x[20] & x[21]);
  assign t[179] = (x[23] & x[24]);
  assign t[17] = ~(t[23] & t[24]);
  assign t[180] = (x[26] & x[27]);
  assign t[181] = (x[29] & x[30]);
  assign t[182] = (x[34] & x[35]);
  assign t[183] = (x[37] & x[38]);
  assign t[184] = (x[40] & x[41]);
  assign t[185] = (x[43] & x[44]);
  assign t[186] = (x[46] & x[47]);
  assign t[187] = (x[49] & x[50]);
  assign t[188] = (x[52] & x[53]);
  assign t[189] = (x[55] & x[56]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[60] & x[61]);
  assign t[191] = (x[63] & x[64]);
  assign t[192] = (x[66] & x[67]);
  assign t[193] = (x[71] & x[72]);
  assign t[194] = (x[74] & x[75]);
  assign t[195] = (x[77] & x[78]);
  assign t[196] = (x[80] & x[81]);
  assign t[197] = (x[83] & x[84]);
  assign t[198] = (x[86] & x[87]);
  assign t[199] = (x[89] & x[90]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[92] & x[93]);
  assign t[201] = (x[95] & x[96]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[34] | t[35]);
  assign t[24] = ~(t[36] | t[37]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[26] = ~(t[149] | t[40]);
  assign t[27] = ~(t[41] | t[42]);
  assign t[28] = ~(t[43] ^ t[44]);
  assign t[29] = ~(t[45] | t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] ^ t[48]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[52]);
  assign t[33] = ~(t[147]);
  assign t[34] = ~(t[53] | t[54]);
  assign t[35] = ~(t[53] | t[55]);
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[150]);
  assign t[39] = ~(t[151]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] | t[60]);
  assign t[41] = ~(t[61] | t[62]);
  assign t[42] = ~(t[152] | t[63]);
  assign t[43] = t[22] ? x[33] : x[32];
  assign t[44] = ~(t[64] & t[65]);
  assign t[45] = ~(t[66] | t[67]);
  assign t[46] = ~(t[153] | t[68]);
  assign t[47] = ~(t[69] | t[70]);
  assign t[48] = ~(t[71] ^ t[72]);
  assign t[49] = ~(t[73] | t[74]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[154] | t[75]);
  assign t[51] = ~(t[76] | t[77]);
  assign t[52] = ~(t[78] ^ t[79]);
  assign t[53] = ~(t[147]);
  assign t[54] = t[145] ? t[81] : t[80];
  assign t[55] = t[145] ? t[83] : t[82];
  assign t[56] = ~(t[84] | t[85]);
  assign t[57] = ~(t[53]);
  assign t[58] = t[145] ? t[86] : t[82];
  assign t[59] = ~(t[155]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[150] | t[151]);
  assign t[61] = ~(t[156]);
  assign t[62] = ~(t[157]);
  assign t[63] = ~(t[87] | t[88]);
  assign t[64] = ~(t[89] | t[35]);
  assign t[65] = ~(t[90] | t[91]);
  assign t[66] = ~(t[158]);
  assign t[67] = ~(t[159]);
  assign t[68] = ~(t[92] | t[93]);
  assign t[69] = ~(t[94] | t[95]);
  assign t[6] = ~(t[7] ^ t[11]);
  assign t[70] = ~(t[160] | t[96]);
  assign t[71] = t[22] ? x[59] : x[58];
  assign t[72] = ~(t[97] & t[98]);
  assign t[73] = ~(t[161]);
  assign t[74] = ~(t[162]);
  assign t[75] = ~(t[99] | t[100]);
  assign t[76] = ~(t[101] | t[102]);
  assign t[77] = ~(t[163] | t[103]);
  assign t[78] = t[104] ? x[70] : x[69];
  assign t[79] = ~(t[105] & t[106]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[107] & t[108]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(x[4] & t[110]);
  assign t[83] = ~(t[111] & t[108]);
  assign t[84] = ~(t[57] | t[112]);
  assign t[85] = ~(t[57] | t[113]);
  assign t[86] = ~(t[148] & t[111]);
  assign t[87] = ~(t[164]);
  assign t[88] = ~(t[156] | t[157]);
  assign t[89] = ~(t[53] | t[114]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[115] & t[116]);
  assign t[91] = ~(t[117] & t[118]);
  assign t[92] = ~(t[165]);
  assign t[93] = ~(t[158] | t[159]);
  assign t[94] = ~(t[166]);
  assign t[95] = ~(t[167]);
  assign t[96] = ~(t[119] | t[120]);
  assign t[97] = ~(t[121] | t[85]);
  assign t[98] = ~(t[122] | t[123]);
  assign t[99] = ~(t[168]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[144];
endmodule

module R1ind134(x, y);
 input [139:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = t[143] ^ x[2];
  assign t[103] = t[144] ^ x[10];
  assign t[104] = t[145] ^ x[13];
  assign t[105] = t[146] ^ x[16];
  assign t[106] = t[147] ^ x[19];
  assign t[107] = t[148] ^ x[22];
  assign t[108] = t[149] ^ x[27];
  assign t[109] = t[150] ^ x[32];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[35];
  assign t[111] = t[152] ^ x[38];
  assign t[112] = t[153] ^ x[41];
  assign t[113] = t[154] ^ x[46];
  assign t[114] = t[155] ^ x[51];
  assign t[115] = t[156] ^ x[54];
  assign t[116] = t[157] ^ x[57];
  assign t[117] = t[158] ^ x[62];
  assign t[118] = t[159] ^ x[67];
  assign t[119] = t[160] ^ x[70];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[73];
  assign t[121] = t[162] ^ x[76];
  assign t[122] = t[163] ^ x[79];
  assign t[123] = t[164] ^ x[82];
  assign t[124] = t[165] ^ x[85];
  assign t[125] = t[166] ^ x[88];
  assign t[126] = t[167] ^ x[91];
  assign t[127] = t[168] ^ x[94];
  assign t[128] = t[169] ^ x[97];
  assign t[129] = t[170] ^ x[100];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[103];
  assign t[131] = t[172] ^ x[106];
  assign t[132] = t[173] ^ x[109];
  assign t[133] = t[174] ^ x[112];
  assign t[134] = t[175] ^ x[115];
  assign t[135] = t[176] ^ x[118];
  assign t[136] = t[177] ^ x[121];
  assign t[137] = t[178] ^ x[124];
  assign t[138] = t[179] ^ x[127];
  assign t[139] = t[180] ^ x[130];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[133];
  assign t[141] = t[182] ^ x[136];
  assign t[142] = t[183] ^ x[139];
  assign t[143] = (x[0] & x[1]);
  assign t[144] = (x[8] & x[9]);
  assign t[145] = (x[11] & x[12]);
  assign t[146] = (x[14] & x[15]);
  assign t[147] = (x[17] & x[18]);
  assign t[148] = (x[20] & x[21]);
  assign t[149] = (x[25] & x[26]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[30] & x[31]);
  assign t[151] = (x[33] & x[34]);
  assign t[152] = (x[36] & x[37]);
  assign t[153] = (x[39] & x[40]);
  assign t[154] = (x[44] & x[45]);
  assign t[155] = (x[49] & x[50]);
  assign t[156] = (x[52] & x[53]);
  assign t[157] = (x[55] & x[56]);
  assign t[158] = (x[60] & x[61]);
  assign t[159] = (x[65] & x[66]);
  assign t[15] = ~(t[103] & t[104]);
  assign t[160] = (x[68] & x[69]);
  assign t[161] = (x[71] & x[72]);
  assign t[162] = (x[74] & x[75]);
  assign t[163] = (x[77] & x[78]);
  assign t[164] = (x[80] & x[81]);
  assign t[165] = (x[83] & x[84]);
  assign t[166] = (x[86] & x[87]);
  assign t[167] = (x[89] & x[90]);
  assign t[168] = (x[92] & x[93]);
  assign t[169] = (x[95] & x[96]);
  assign t[16] = ~(t[105] & t[106]);
  assign t[170] = (x[98] & x[99]);
  assign t[171] = (x[101] & x[102]);
  assign t[172] = (x[104] & x[105]);
  assign t[173] = (x[107] & x[108]);
  assign t[174] = (x[110] & x[111]);
  assign t[175] = (x[113] & x[114]);
  assign t[176] = (x[116] & x[117]);
  assign t[177] = (x[119] & x[120]);
  assign t[178] = (x[122] & x[123]);
  assign t[179] = (x[125] & x[126]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[128] & x[129]);
  assign t[181] = (x[131] & x[132]);
  assign t[182] = (x[134] & x[135]);
  assign t[183] = (x[137] & x[138]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[105]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[107];
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[42];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] | t[108];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[109]);
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[68] & t[69]);
  assign t[49] = t[70] | t[111];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = t[73] | t[112];
  assign t[52] = t[74] ? x[43] : x[42];
  assign t[53] = ~(t[75] & t[76]);
  assign t[54] = t[77] | t[113];
  assign t[55] = t[74] ? x[48] : x[47];
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[78] | t[56]);
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[81] | t[116];
  assign t[61] = t[74] ? x[59] : x[58];
  assign t[62] = ~(t[82] & t[83]);
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = t[86] | t[117];
  assign t[65] = t[17] ? x[64] : x[63];
  assign t[66] = ~(t[87] & t[88]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[121]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[90] | t[71]);
  assign t[74] = ~(t[24]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[91] | t[75]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[92] | t[79]);
  assign t[82] = ~(t[93] & t[94]);
  assign t[83] = t[95] | t[128];
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[137]);
  assign t[95] = ~(t[100] | t[93]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[102];
endmodule

module R1ind135(x, y);
 input [139:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[107] & t[108]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[146] & t[145]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[151]);
  assign t[111] = t[152] ^ x[2];
  assign t[112] = t[153] ^ x[10];
  assign t[113] = t[154] ^ x[13];
  assign t[114] = t[155] ^ x[16];
  assign t[115] = t[156] ^ x[19];
  assign t[116] = t[157] ^ x[22];
  assign t[117] = t[158] ^ x[27];
  assign t[118] = t[159] ^ x[32];
  assign t[119] = t[160] ^ x[35];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[38];
  assign t[121] = t[162] ^ x[41];
  assign t[122] = t[163] ^ x[46];
  assign t[123] = t[164] ^ x[51];
  assign t[124] = t[165] ^ x[54];
  assign t[125] = t[166] ^ x[57];
  assign t[126] = t[167] ^ x[62];
  assign t[127] = t[168] ^ x[67];
  assign t[128] = t[169] ^ x[70];
  assign t[129] = t[170] ^ x[73];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[76];
  assign t[131] = t[172] ^ x[79];
  assign t[132] = t[173] ^ x[82];
  assign t[133] = t[174] ^ x[85];
  assign t[134] = t[175] ^ x[88];
  assign t[135] = t[176] ^ x[91];
  assign t[136] = t[177] ^ x[94];
  assign t[137] = t[178] ^ x[97];
  assign t[138] = t[179] ^ x[100];
  assign t[139] = t[180] ^ x[103];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[106];
  assign t[141] = t[182] ^ x[109];
  assign t[142] = t[183] ^ x[112];
  assign t[143] = t[184] ^ x[115];
  assign t[144] = t[185] ^ x[118];
  assign t[145] = t[186] ^ x[121];
  assign t[146] = t[187] ^ x[124];
  assign t[147] = t[188] ^ x[127];
  assign t[148] = t[189] ^ x[130];
  assign t[149] = t[190] ^ x[133];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[136];
  assign t[151] = t[192] ^ x[139];
  assign t[152] = (x[0] & x[1]);
  assign t[153] = (x[8] & x[9]);
  assign t[154] = (x[11] & x[12]);
  assign t[155] = (x[14] & x[15]);
  assign t[156] = (x[17] & x[18]);
  assign t[157] = (x[20] & x[21]);
  assign t[158] = (x[25] & x[26]);
  assign t[159] = (x[30] & x[31]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[33] & x[34]);
  assign t[161] = (x[36] & x[37]);
  assign t[162] = (x[39] & x[40]);
  assign t[163] = (x[44] & x[45]);
  assign t[164] = (x[49] & x[50]);
  assign t[165] = (x[52] & x[53]);
  assign t[166] = (x[55] & x[56]);
  assign t[167] = (x[60] & x[61]);
  assign t[168] = (x[65] & x[66]);
  assign t[169] = (x[68] & x[69]);
  assign t[16] = ~(t[114] & t[115]);
  assign t[170] = (x[71] & x[72]);
  assign t[171] = (x[74] & x[75]);
  assign t[172] = (x[77] & x[78]);
  assign t[173] = (x[80] & x[81]);
  assign t[174] = (x[83] & x[84]);
  assign t[175] = (x[86] & x[87]);
  assign t[176] = (x[89] & x[90]);
  assign t[177] = (x[92] & x[93]);
  assign t[178] = (x[95] & x[96]);
  assign t[179] = (x[98] & x[99]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[101] & x[102]);
  assign t[181] = (x[104] & x[105]);
  assign t[182] = (x[107] & x[108]);
  assign t[183] = (x[110] & x[111]);
  assign t[184] = (x[113] & x[114]);
  assign t[185] = (x[116] & x[117]);
  assign t[186] = (x[119] & x[120]);
  assign t[187] = (x[122] & x[123]);
  assign t[188] = (x[125] & x[126]);
  assign t[189] = (x[128] & x[129]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[131] & x[132]);
  assign t[191] = (x[134] & x[135]);
  assign t[192] = (x[137] & x[138]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[114]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[116]);
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[42];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = ~(t[58] & t[117]);
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[118]);
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[67] & t[68]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = ~(t[71] & t[120]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[74] & t[121]);
  assign t[52] = t[75] ? x[43] : x[42];
  assign t[53] = ~(t[76] & t[77]);
  assign t[54] = ~(t[78] & t[122]);
  assign t[55] = t[75] ? x[48] : x[47];
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[125]);
  assign t[61] = t[75] ? x[59] : x[58];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[126]);
  assign t[65] = t[17] ? x[64] : x[63];
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[91] & t[92]);
  assign t[72] = ~(t[130]);
  assign t[73] = ~(t[131]);
  assign t[74] = ~(t[93] & t[94]);
  assign t[75] = ~(t[24]);
  assign t[76] = ~(t[132]);
  assign t[77] = ~(t[133]);
  assign t[78] = ~(t[95] & t[96]);
  assign t[79] = ~(t[124] & t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[97] & t[98]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[101] & t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[133] & t[132]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[136] & t[135]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[111];
endmodule

module R1ind136(x, y);
 input [112:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[30];
  assign t[101] = t[133] ^ x[33];
  assign t[102] = t[134] ^ x[38];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[44];
  assign t[105] = t[137] ^ x[47];
  assign t[106] = t[138] ^ x[50];
  assign t[107] = t[139] ^ x[55];
  assign t[108] = t[140] ^ x[58];
  assign t[109] = t[141] ^ x[63];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[66];
  assign t[111] = t[143] ^ x[69];
  assign t[112] = t[144] ^ x[74];
  assign t[113] = t[145] ^ x[77];
  assign t[114] = t[146] ^ x[82];
  assign t[115] = t[147] ^ x[85];
  assign t[116] = t[148] ^ x[88];
  assign t[117] = t[149] ^ x[91];
  assign t[118] = t[150] ^ x[94];
  assign t[119] = t[151] ^ x[97];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[152] ^ x[100];
  assign t[121] = t[153] ^ x[103];
  assign t[122] = t[154] ^ x[106];
  assign t[123] = t[155] ^ x[109];
  assign t[124] = t[156] ^ x[112];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[23] & x[24]);
  assign t[132] = (x[28] & x[29]);
  assign t[133] = (x[31] & x[32]);
  assign t[134] = (x[36] & x[37]);
  assign t[135] = (x[39] & x[40]);
  assign t[136] = (x[42] & x[43]);
  assign t[137] = (x[45] & x[46]);
  assign t[138] = (x[48] & x[49]);
  assign t[139] = (x[53] & x[54]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[56] & x[57]);
  assign t[141] = (x[61] & x[62]);
  assign t[142] = (x[64] & x[65]);
  assign t[143] = (x[67] & x[68]);
  assign t[144] = (x[72] & x[73]);
  assign t[145] = (x[75] & x[76]);
  assign t[146] = (x[80] & x[81]);
  assign t[147] = (x[83] & x[84]);
  assign t[148] = (x[86] & x[87]);
  assign t[149] = (x[89] & x[90]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[92] & x[93]);
  assign t[151] = (x[95] & x[96]);
  assign t[152] = (x[98] & x[99]);
  assign t[153] = (x[101] & x[102]);
  assign t[154] = (x[104] & x[105]);
  assign t[155] = (x[107] & x[108]);
  assign t[156] = (x[110] & x[111]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[46] ? x[27] : x[26];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = t[51] ^ t[42];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[33];
  assign t[37] = ~(t[100] & t[55]);
  assign t[38] = ~(t[101] & t[56]);
  assign t[39] = t[17] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = t[59] ^ t[60];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[65]);
  assign t[46] = ~(t[24]);
  assign t[47] = ~(t[103] & t[66]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[106] & t[69]);
  assign t[51] = t[70] ? x[52] : x[51];
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = t[70] ? x[60] : x[59];
  assign t[55] = ~(t[109]);
  assign t[56] = ~(t[109] & t[73]);
  assign t[57] = ~(t[110] & t[74]);
  assign t[58] = ~(t[111] & t[75]);
  assign t[59] = t[70] ? x[71] : x[70];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[76] & t[77]);
  assign t[61] = ~(t[112] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = t[17] ? x[79] : x[78];
  assign t[64] = ~(t[80] & t[81]);
  assign t[65] = ~(t[98]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[115]);
  assign t[69] = ~(t[115] & t[83]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[24]);
  assign t[71] = ~(t[116]);
  assign t[72] = ~(t[116] & t[84]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[117]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[107]);
  assign t[85] = ~(t[110]);
  assign t[86] = ~(t[123]);
  assign t[87] = ~(t[123] & t[91]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[124]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[124] & t[92]);
  assign t[91] = ~(t[118]);
  assign t[92] = ~(t[121]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[25];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind137(x, y);
 input [139:0] x;
 output y;

 wire [278:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[136] ? x[81] : x[80];
  assign t[101] = ~(t[141] & t[105]);
  assign t[102] = ~(t[220]);
  assign t[103] = ~(t[209] | t[210]);
  assign t[104] = ~(t[124] | t[49]);
  assign t[105] = ~(t[142] | t[138]);
  assign t[106] = ~(t[221]);
  assign t[107] = ~(t[222]);
  assign t[108] = ~(t[143] | t[144]);
  assign t[109] = ~(t[145] | t[146]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[223] | t[147]);
  assign t[111] = t[29] ? x[95] : x[94];
  assign t[112] = ~(t[148] & t[149]);
  assign t[113] = ~(t[224]);
  assign t[114] = ~(t[225]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[152] | t[153]);
  assign t[117] = ~(t[226] | t[154]);
  assign t[118] = t[136] ? x[106] : x[105];
  assign t[119] = ~(t[155] & t[156]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[158]);
  assign t[122] = ~(x[4] & t[160]);
  assign t[123] = ~(t[161] & t[158]);
  assign t[124] = ~(t[78] | t[162]);
  assign t[125] = ~(t[163] | t[164]);
  assign t[126] = ~(t[122] & t[165]);
  assign t[127] = t[201] & t[166];
  assign t[128] = t[157] | t[159];
  assign t[129] = t[198] ? t[122] : t[123];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[227]);
  assign t[131] = ~(t[214] | t[215]);
  assign t[132] = ~(t[167] & t[168]);
  assign t[133] = t[138] | t[169];
  assign t[134] = ~(t[228]);
  assign t[135] = ~(t[216] | t[217]);
  assign t[136] = ~(t[47]);
  assign t[137] = ~(t[30] & t[168]);
  assign t[138] = ~(t[163] | t[170]);
  assign t[139] = ~(t[229]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[218] | t[219]);
  assign t[141] = ~(t[171]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[230]);
  assign t[144] = ~(t[221] | t[222]);
  assign t[145] = ~(t[231]);
  assign t[146] = ~(t[232]);
  assign t[147] = ~(t[173] | t[174]);
  assign t[148] = ~(t[175] | t[176]);
  assign t[149] = ~(t[127] | t[177]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[233]);
  assign t[151] = ~(t[224] | t[225]);
  assign t[152] = ~(t[234]);
  assign t[153] = ~(t[235]);
  assign t[154] = ~(t[178] | t[179]);
  assign t[155] = ~(t[180] | t[181]);
  assign t[156] = ~(t[182]);
  assign t[157] = ~(x[4] | t[199]);
  assign t[158] = ~(t[201]);
  assign t[159] = x[4] & t[199];
  assign t[15] = ~(t[198] & t[199]);
  assign t[160] = ~(t[199] | t[201]);
  assign t[161] = ~(x[4] | t[183]);
  assign t[162] = t[198] ? t[120] : t[121];
  assign t[163] = ~(t[78]);
  assign t[164] = t[198] ? t[123] : t[184];
  assign t[165] = ~(t[201] & t[161]);
  assign t[166] = ~(t[78] | t[198]);
  assign t[167] = ~(t[166] & t[185]);
  assign t[168] = ~(t[186] & t[187]);
  assign t[169] = ~(t[163] | t[188]);
  assign t[16] = ~(t[200] & t[201]);
  assign t[170] = t[198] ? t[165] : t[122];
  assign t[171] = ~(t[163] | t[189]);
  assign t[172] = ~(t[180] | t[176]);
  assign t[173] = ~(t[236]);
  assign t[174] = ~(t[231] | t[232]);
  assign t[175] = ~(t[163] | t[190]);
  assign t[176] = ~(t[163] | t[191]);
  assign t[177] = ~(t[30]);
  assign t[178] = ~(t[237]);
  assign t[179] = ~(t[234] | t[235]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[163] | t[192]);
  assign t[181] = ~(t[193] & t[30]);
  assign t[182] = ~(t[163] | t[194]);
  assign t[183] = ~(t[199]);
  assign t[184] = ~(x[4] & t[186]);
  assign t[185] = ~(t[165] & t[184]);
  assign t[186] = ~(t[199] | t[158]);
  assign t[187] = t[163] & t[198];
  assign t[188] = t[198] ? t[195] : t[121];
  assign t[189] = t[198] ? t[196] : t[120];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[198] ? t[122] : t[165];
  assign t[191] = t[198] ? t[121] : t[195];
  assign t[192] = t[198] ? t[184] : t[123];
  assign t[193] = ~(t[171] | t[50]);
  assign t[194] = t[198] ? t[120] : t[196];
  assign t[195] = ~(t[157] & t[201]);
  assign t[196] = ~(t[159] & t[201]);
  assign t[197] = t[238] ^ x[2];
  assign t[198] = t[239] ^ x[10];
  assign t[199] = t[240] ^ x[13];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[16];
  assign t[201] = t[242] ^ x[19];
  assign t[202] = t[243] ^ x[22];
  assign t[203] = t[244] ^ x[25];
  assign t[204] = t[245] ^ x[28];
  assign t[205] = t[246] ^ x[31];
  assign t[206] = t[247] ^ x[34];
  assign t[207] = t[248] ^ x[39];
  assign t[208] = t[249] ^ x[42];
  assign t[209] = t[250] ^ x[45];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[48];
  assign t[211] = t[252] ^ x[53];
  assign t[212] = t[253] ^ x[56];
  assign t[213] = t[254] ^ x[59];
  assign t[214] = t[255] ^ x[62];
  assign t[215] = t[256] ^ x[65];
  assign t[216] = t[257] ^ x[68];
  assign t[217] = t[258] ^ x[71];
  assign t[218] = t[259] ^ x[76];
  assign t[219] = t[260] ^ x[79];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[84];
  assign t[221] = t[262] ^ x[87];
  assign t[222] = t[263] ^ x[90];
  assign t[223] = t[264] ^ x[93];
  assign t[224] = t[265] ^ x[98];
  assign t[225] = t[266] ^ x[101];
  assign t[226] = t[267] ^ x[104];
  assign t[227] = t[268] ^ x[109];
  assign t[228] = t[269] ^ x[112];
  assign t[229] = t[270] ^ x[115];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[271] ^ x[118];
  assign t[231] = t[272] ^ x[121];
  assign t[232] = t[273] ^ x[124];
  assign t[233] = t[274] ^ x[127];
  assign t[234] = t[275] ^ x[130];
  assign t[235] = t[276] ^ x[133];
  assign t[236] = t[277] ^ x[136];
  assign t[237] = t[278] ^ x[139];
  assign t[238] = (x[0] & x[1]);
  assign t[239] = (x[8] & x[9]);
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = (x[11] & x[12]);
  assign t[241] = (x[14] & x[15]);
  assign t[242] = (x[17] & x[18]);
  assign t[243] = (x[20] & x[21]);
  assign t[244] = (x[23] & x[24]);
  assign t[245] = (x[26] & x[27]);
  assign t[246] = (x[29] & x[30]);
  assign t[247] = (x[32] & x[33]);
  assign t[248] = (x[37] & x[38]);
  assign t[249] = (x[40] & x[41]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[43] & x[44]);
  assign t[251] = (x[46] & x[47]);
  assign t[252] = (x[51] & x[52]);
  assign t[253] = (x[54] & x[55]);
  assign t[254] = (x[57] & x[58]);
  assign t[255] = (x[60] & x[61]);
  assign t[256] = (x[63] & x[64]);
  assign t[257] = (x[66] & x[67]);
  assign t[258] = (x[69] & x[70]);
  assign t[259] = (x[74] & x[75]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[77] & x[78]);
  assign t[261] = (x[82] & x[83]);
  assign t[262] = (x[85] & x[86]);
  assign t[263] = (x[88] & x[89]);
  assign t[264] = (x[91] & x[92]);
  assign t[265] = (x[96] & x[97]);
  assign t[266] = (x[99] & x[100]);
  assign t[267] = (x[102] & x[103]);
  assign t[268] = (x[107] & x[108]);
  assign t[269] = (x[110] & x[111]);
  assign t[26] = ~(t[25] ^ t[42]);
  assign t[270] = (x[113] & x[114]);
  assign t[271] = (x[116] & x[117]);
  assign t[272] = (x[119] & x[120]);
  assign t[273] = (x[122] & x[123]);
  assign t[274] = (x[125] & x[126]);
  assign t[275] = (x[128] & x[129]);
  assign t[276] = (x[131] & x[132]);
  assign t[277] = (x[134] & x[135]);
  assign t[278] = (x[137] & x[138]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[202] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[38] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[43] ^ t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[203] | t[67]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[200]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[78] | t[80]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81] & t[82]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = ~(t[204]);
  assign t[53] = ~(t[205]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[206] | t[89]);
  assign t[57] = t[90] ? x[36] : x[35];
  assign t[58] = ~(t[91] & t[83]);
  assign t[59] = ~(t[92] | t[93]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[207] | t[94]);
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = ~(t[97] | t[98]);
  assign t[63] = ~(t[208] | t[99]);
  assign t[64] = ~(t[100] ^ t[101]);
  assign t[65] = ~(t[209]);
  assign t[66] = ~(t[210]);
  assign t[67] = ~(t[102] | t[103]);
  assign t[68] = t[29] ? x[50] : x[49];
  assign t[69] = ~(t[104] & t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[211] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[212] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[200]);
  assign t[79] = t[198] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[198] ? t[123] : t[122];
  assign t[81] = ~(t[124] | t[125]);
  assign t[82] = ~(t[78] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = t[78] | t[129];
  assign t[85] = ~(t[213]);
  assign t[86] = ~(t[204] | t[205]);
  assign t[87] = ~(t[214]);
  assign t[88] = ~(t[215]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[47]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[216]);
  assign t[93] = ~(t[217]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = t[136] ? x[73] : x[72];
  assign t[96] = t[137] | t[138];
  assign t[97] = ~(t[218]);
  assign t[98] = ~(t[219]);
  assign t[99] = ~(t[139] | t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[197];
endmodule

module R1ind138(x, y);
 input [139:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = t[142] ^ x[2];
  assign t[102] = t[143] ^ x[10];
  assign t[103] = t[144] ^ x[13];
  assign t[104] = t[145] ^ x[16];
  assign t[105] = t[146] ^ x[19];
  assign t[106] = t[147] ^ x[22];
  assign t[107] = t[148] ^ x[27];
  assign t[108] = t[149] ^ x[32];
  assign t[109] = t[150] ^ x[35];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[38];
  assign t[111] = t[152] ^ x[43];
  assign t[112] = t[153] ^ x[48];
  assign t[113] = t[154] ^ x[51];
  assign t[114] = t[155] ^ x[54];
  assign t[115] = t[156] ^ x[57];
  assign t[116] = t[157] ^ x[62];
  assign t[117] = t[158] ^ x[67];
  assign t[118] = t[159] ^ x[70];
  assign t[119] = t[160] ^ x[73];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[76];
  assign t[121] = t[162] ^ x[79];
  assign t[122] = t[163] ^ x[82];
  assign t[123] = t[164] ^ x[85];
  assign t[124] = t[165] ^ x[88];
  assign t[125] = t[166] ^ x[91];
  assign t[126] = t[167] ^ x[94];
  assign t[127] = t[168] ^ x[97];
  assign t[128] = t[169] ^ x[100];
  assign t[129] = t[170] ^ x[103];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[106];
  assign t[131] = t[172] ^ x[109];
  assign t[132] = t[173] ^ x[112];
  assign t[133] = t[174] ^ x[115];
  assign t[134] = t[175] ^ x[118];
  assign t[135] = t[176] ^ x[121];
  assign t[136] = t[177] ^ x[124];
  assign t[137] = t[178] ^ x[127];
  assign t[138] = t[179] ^ x[130];
  assign t[139] = t[180] ^ x[133];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[136];
  assign t[141] = t[182] ^ x[139];
  assign t[142] = (x[0] & x[1]);
  assign t[143] = (x[8] & x[9]);
  assign t[144] = (x[11] & x[12]);
  assign t[145] = (x[14] & x[15]);
  assign t[146] = (x[17] & x[18]);
  assign t[147] = (x[20] & x[21]);
  assign t[148] = (x[25] & x[26]);
  assign t[149] = (x[30] & x[31]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[33] & x[34]);
  assign t[151] = (x[36] & x[37]);
  assign t[152] = (x[41] & x[42]);
  assign t[153] = (x[46] & x[47]);
  assign t[154] = (x[49] & x[50]);
  assign t[155] = (x[52] & x[53]);
  assign t[156] = (x[55] & x[56]);
  assign t[157] = (x[60] & x[61]);
  assign t[158] = (x[65] & x[66]);
  assign t[159] = (x[68] & x[69]);
  assign t[15] = ~(t[102] & t[103]);
  assign t[160] = (x[71] & x[72]);
  assign t[161] = (x[74] & x[75]);
  assign t[162] = (x[77] & x[78]);
  assign t[163] = (x[80] & x[81]);
  assign t[164] = (x[83] & x[84]);
  assign t[165] = (x[86] & x[87]);
  assign t[166] = (x[89] & x[90]);
  assign t[167] = (x[92] & x[93]);
  assign t[168] = (x[95] & x[96]);
  assign t[169] = (x[98] & x[99]);
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = (x[101] & x[102]);
  assign t[171] = (x[104] & x[105]);
  assign t[172] = (x[107] & x[108]);
  assign t[173] = (x[110] & x[111]);
  assign t[174] = (x[113] & x[114]);
  assign t[175] = (x[116] & x[117]);
  assign t[176] = (x[119] & x[120]);
  assign t[177] = (x[122] & x[123]);
  assign t[178] = (x[125] & x[126]);
  assign t[179] = (x[128] & x[129]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[131] & x[132]);
  assign t[181] = (x[134] & x[135]);
  assign t[182] = (x[137] & x[138]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[104]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[106];
  assign t[31] = t[104] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[107];
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[108]);
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[70] | t[110];
  assign t[49] = t[104] ? x[40] : x[39];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = t[75] | t[111];
  assign t[53] = t[104] ? x[45] : x[44];
  assign t[54] = ~(t[112]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[76] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[77] & t[78]);
  assign t[59] = t[79] | t[114];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[80] & t[81]);
  assign t[61] = t[82] | t[115];
  assign t[62] = t[17] ? x[59] : x[58];
  assign t[63] = ~(t[83] & t[84]);
  assign t[64] = t[85] | t[116];
  assign t[65] = t[17] ? x[64] : x[63];
  assign t[66] = ~(t[86] & t[87]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[88] | t[68]);
  assign t[71] = ~(t[89] & t[90]);
  assign t[72] = t[91] | t[120];
  assign t[73] = ~(t[121]);
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[92] | t[73]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[93] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[94] | t[80]);
  assign t[83] = ~(t[128]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[95] | t[83]);
  assign t[86] = ~(t[96] & t[97]);
  assign t[87] = t[98] | t[130];
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[99] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[100] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[101];
endmodule

module R1ind139(x, y);
 input [139:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[108] & t[109]);
  assign t[106] = ~(t[142] & t[141]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[32];
  assign t[118] = t[159] ^ x[35];
  assign t[119] = t[160] ^ x[38];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[43];
  assign t[121] = t[162] ^ x[48];
  assign t[122] = t[163] ^ x[51];
  assign t[123] = t[164] ^ x[54];
  assign t[124] = t[165] ^ x[57];
  assign t[125] = t[166] ^ x[62];
  assign t[126] = t[167] ^ x[67];
  assign t[127] = t[168] ^ x[70];
  assign t[128] = t[169] ^ x[73];
  assign t[129] = t[170] ^ x[76];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[79];
  assign t[131] = t[172] ^ x[82];
  assign t[132] = t[173] ^ x[85];
  assign t[133] = t[174] ^ x[88];
  assign t[134] = t[175] ^ x[91];
  assign t[135] = t[176] ^ x[94];
  assign t[136] = t[177] ^ x[97];
  assign t[137] = t[178] ^ x[100];
  assign t[138] = t[179] ^ x[103];
  assign t[139] = t[180] ^ x[106];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[109];
  assign t[141] = t[182] ^ x[112];
  assign t[142] = t[183] ^ x[115];
  assign t[143] = t[184] ^ x[118];
  assign t[144] = t[185] ^ x[121];
  assign t[145] = t[186] ^ x[124];
  assign t[146] = t[187] ^ x[127];
  assign t[147] = t[188] ^ x[130];
  assign t[148] = t[189] ^ x[133];
  assign t[149] = t[190] ^ x[136];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[139];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[30] & x[31]);
  assign t[159] = (x[33] & x[34]);
  assign t[15] = ~(t[111] & t[112]);
  assign t[160] = (x[36] & x[37]);
  assign t[161] = (x[41] & x[42]);
  assign t[162] = (x[46] & x[47]);
  assign t[163] = (x[49] & x[50]);
  assign t[164] = (x[52] & x[53]);
  assign t[165] = (x[55] & x[56]);
  assign t[166] = (x[60] & x[61]);
  assign t[167] = (x[65] & x[66]);
  assign t[168] = (x[68] & x[69]);
  assign t[169] = (x[71] & x[72]);
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = (x[74] & x[75]);
  assign t[171] = (x[77] & x[78]);
  assign t[172] = (x[80] & x[81]);
  assign t[173] = (x[83] & x[84]);
  assign t[174] = (x[86] & x[87]);
  assign t[175] = (x[89] & x[90]);
  assign t[176] = (x[92] & x[93]);
  assign t[177] = (x[95] & x[96]);
  assign t[178] = (x[98] & x[99]);
  assign t[179] = (x[101] & x[102]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[104] & x[105]);
  assign t[181] = (x[107] & x[108]);
  assign t[182] = (x[110] & x[111]);
  assign t[183] = (x[113] & x[114]);
  assign t[184] = (x[116] & x[117]);
  assign t[185] = (x[119] & x[120]);
  assign t[186] = (x[122] & x[123]);
  assign t[187] = (x[125] & x[126]);
  assign t[188] = (x[128] & x[129]);
  assign t[189] = (x[131] & x[132]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[134] & x[135]);
  assign t[191] = (x[137] & x[138]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[113]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[115]);
  assign t[31] = t[113] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = ~(t[56] & t[116]);
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[117]);
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[67] & t[68]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[71] & t[119]);
  assign t[49] = t[113] ? x[40] : x[39];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = ~(t[76] & t[120]);
  assign t[53] = t[113] ? x[45] : x[44];
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[77] & t[78]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[123]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[124]);
  assign t[62] = t[17] ? x[59] : x[58];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[87] & t[125]);
  assign t[65] = t[17] ? x[64] : x[63];
  assign t[66] = ~(t[88] & t[89]);
  assign t[67] = ~(t[118] & t[117]);
  assign t[68] = ~(t[126]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = ~(t[92] & t[93]);
  assign t[73] = ~(t[94] & t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[122] & t[121]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[97] & t[98]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[101] & t[102]);
  assign t[88] = ~(t[103] & t[104]);
  assign t[89] = ~(t[105] & t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[106] & t[107]);
  assign t[95] = ~(t[131] & t[130]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind140(x, y);
 input [112:0] x;
 output y;

 wire [155:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[33];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[41];
  assign t[103] = t[135] ^ x[44];
  assign t[104] = t[136] ^ x[49];
  assign t[105] = t[137] ^ x[52];
  assign t[106] = t[138] ^ x[57];
  assign t[107] = t[139] ^ x[60];
  assign t[108] = t[140] ^ x[63];
  assign t[109] = t[141] ^ x[66];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[69];
  assign t[111] = t[143] ^ x[74];
  assign t[112] = t[144] ^ x[77];
  assign t[113] = t[145] ^ x[82];
  assign t[114] = t[146] ^ x[85];
  assign t[115] = t[147] ^ x[88];
  assign t[116] = t[148] ^ x[91];
  assign t[117] = t[149] ^ x[94];
  assign t[118] = t[150] ^ x[97];
  assign t[119] = t[151] ^ x[100];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[152] ^ x[103];
  assign t[121] = t[153] ^ x[106];
  assign t[122] = t[154] ^ x[109];
  assign t[123] = t[155] ^ x[112];
  assign t[124] = (x[0] & x[1]);
  assign t[125] = (x[8] & x[9]);
  assign t[126] = (x[11] & x[12]);
  assign t[127] = (x[14] & x[15]);
  assign t[128] = (x[17] & x[18]);
  assign t[129] = (x[20] & x[21]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[23] & x[24]);
  assign t[131] = (x[28] & x[29]);
  assign t[132] = (x[31] & x[32]);
  assign t[133] = (x[36] & x[37]);
  assign t[134] = (x[39] & x[40]);
  assign t[135] = (x[42] & x[43]);
  assign t[136] = (x[47] & x[48]);
  assign t[137] = (x[50] & x[51]);
  assign t[138] = (x[55] & x[56]);
  assign t[139] = (x[58] & x[59]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[61] & x[62]);
  assign t[141] = (x[64] & x[65]);
  assign t[142] = (x[67] & x[68]);
  assign t[143] = (x[72] & x[73]);
  assign t[144] = (x[75] & x[76]);
  assign t[145] = (x[80] & x[81]);
  assign t[146] = (x[83] & x[84]);
  assign t[147] = (x[86] & x[87]);
  assign t[148] = (x[89] & x[90]);
  assign t[149] = (x[92] & x[93]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[95] & x[96]);
  assign t[151] = (x[98] & x[99]);
  assign t[152] = (x[101] & x[102]);
  assign t[153] = (x[104] & x[105]);
  assign t[154] = (x[107] & x[108]);
  assign t[155] = (x[110] & x[111]);
  assign t[15] = ~(t[93] & t[94]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[95]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[97] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[98] & t[45]);
  assign t[31] = t[95] ? x[27] : x[26];
  assign t[32] = ~(t[46] & t[47]);
  assign t[33] = t[48] ^ t[32];
  assign t[34] = ~(t[49] & t[50]);
  assign t[35] = t[51] ^ t[52];
  assign t[36] = ~(t[99] & t[53]);
  assign t[37] = ~(t[100] & t[54]);
  assign t[38] = t[55] ? x[35] : x[34];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[61];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[42];
  assign t[44] = ~(t[101]);
  assign t[45] = ~(t[101] & t[65]);
  assign t[46] = ~(t[102] & t[66]);
  assign t[47] = ~(t[103] & t[67]);
  assign t[48] = t[95] ? x[46] : x[45];
  assign t[49] = ~(t[104] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = t[95] ? x[54] : x[53];
  assign t[52] = ~(t[70] & t[71]);
  assign t[53] = ~(t[106]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[24]);
  assign t[56] = ~(t[107] & t[73]);
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[17] ? x[71] : x[70];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[111] & t[79]);
  assign t[63] = ~(t[112] & t[80]);
  assign t[64] = t[17] ? x[79] : x[78];
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[113]);
  assign t[67] = ~(t[113] & t[81]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[99]);
  assign t[73] = ~(t[117]);
  assign t[74] = ~(t[117] & t[85]);
  assign t[75] = ~(t[118]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[102]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[122]);
  assign t[84] = ~(t[122] & t[90]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[123]);
  assign t[88] = ~(t[123] & t[91]);
  assign t[89] = ~(t[111]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[115]);
  assign t[91] = ~(t[119]);
  assign t[92] = t[124] ^ x[2];
  assign t[93] = t[125] ^ x[10];
  assign t[94] = t[126] ^ x[13];
  assign t[95] = t[127] ^ x[16];
  assign t[96] = t[128] ^ x[19];
  assign t[97] = t[129] ^ x[22];
  assign t[98] = t[130] ^ x[25];
  assign t[99] = t[131] ^ x[30];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[92];
endmodule

module R1ind141(x, y);
 input [139:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[211] | t[212]);
  assign t[101] = ~(t[223]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[139] | t[140]);
  assign t[104] = ~(t[47]);
  assign t[105] = ~(t[128] | t[141]);
  assign t[106] = ~(t[126]);
  assign t[107] = ~(t[225]);
  assign t[108] = ~(t[226]);
  assign t[109] = ~(t[142] | t[143]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[29] ? x[95] : x[94];
  assign t[111] = ~(t[144] & t[145]);
  assign t[112] = ~(t[227]);
  assign t[113] = ~(t[228]);
  assign t[114] = ~(t[146] | t[147]);
  assign t[115] = ~(t[148] | t[149]);
  assign t[116] = ~(t[229] | t[150]);
  assign t[117] = t[29] ? x[106] : x[105];
  assign t[118] = ~(t[82] & t[151]);
  assign t[119] = ~(t[203]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[204] & t[152]);
  assign t[121] = ~(x[4] & t[153]);
  assign t[122] = ~(t[154] & t[204]);
  assign t[123] = ~(t[155] & t[156]);
  assign t[124] = ~(t[119] | t[157]);
  assign t[125] = ~(t[119] | t[158]);
  assign t[126] = ~(t[78] | t[159]);
  assign t[127] = ~(t[160] & t[161]);
  assign t[128] = ~(t[78] | t[162]);
  assign t[129] = ~(t[230]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[217] | t[218]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[163] | t[164]);
  assign t[134] = ~(t[137] | t[165]);
  assign t[135] = ~(t[233]);
  assign t[136] = ~(t[220] | t[221]);
  assign t[137] = ~(t[166] & t[167]);
  assign t[138] = ~(t[168] & t[30]);
  assign t[139] = ~(t[234]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[223] | t[224]);
  assign t[141] = ~(t[169] & t[82]);
  assign t[142] = ~(t[235]);
  assign t[143] = ~(t[225] | t[226]);
  assign t[144] = ~(t[170] | t[125]);
  assign t[145] = ~(t[171] | t[172]);
  assign t[146] = ~(t[236]);
  assign t[147] = ~(t[227] | t[228]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[238]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[173] | t[174]);
  assign t[151] = ~(t[175] | t[176]);
  assign t[152] = ~(x[4] | t[177]);
  assign t[153] = ~(t[202] | t[204]);
  assign t[154] = ~(x[4] | t[202]);
  assign t[155] = x[4] & t[202];
  assign t[156] = ~(t[204]);
  assign t[157] = t[201] ? t[123] : t[178];
  assign t[158] = t[201] ? t[179] : t[121];
  assign t[159] = t[201] ? t[178] : t[180];
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = ~(t[181] | t[48]);
  assign t[161] = ~(t[50] & t[182]);
  assign t[162] = t[201] ? t[183] : t[179];
  assign t[163] = ~(t[239]);
  assign t[164] = ~(t[231] | t[232]);
  assign t[165] = ~(t[184] & t[185]);
  assign t[166] = ~(t[81] & t[186]);
  assign t[167] = ~(t[187] & t[188]);
  assign t[168] = ~(t[126] | t[189]);
  assign t[169] = ~(t[181] | t[175]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[119] | t[190]);
  assign t[171] = ~(t[86]);
  assign t[172] = ~(t[78] | t[191]);
  assign t[173] = ~(t[240]);
  assign t[174] = ~(t[237] | t[238]);
  assign t[175] = ~(t[192] & t[193]);
  assign t[176] = ~(t[161] & t[185]);
  assign t[177] = ~(t[202]);
  assign t[178] = ~(t[154] & t[156]);
  assign t[179] = ~(t[152] & t[156]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[155] & t[204]);
  assign t[181] = ~(t[78] | t[194]);
  assign t[182] = t[154] | t[155];
  assign t[183] = ~(x[4] & t[187]);
  assign t[184] = ~(t[125]);
  assign t[185] = t[119] | t[195];
  assign t[186] = ~(t[120] & t[183]);
  assign t[187] = ~(t[202] | t[156]);
  assign t[188] = t[78] & t[201];
  assign t[189] = ~(t[78] | t[196]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[201] ? t[178] : t[123];
  assign t[191] = t[201] ? t[120] : t[121];
  assign t[192] = ~(t[170] | t[197]);
  assign t[193] = ~(t[119] & t[198]);
  assign t[194] = t[201] ? t[180] : t[178];
  assign t[195] = t[201] ? t[121] : t[179];
  assign t[196] = t[201] ? t[122] : t[123];
  assign t[197] = ~(t[78] | t[199]);
  assign t[198] = ~(t[121] & t[120]);
  assign t[199] = t[201] ? t[179] : t[183];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[10];
  assign t[202] = t[243] ^ x[13];
  assign t[203] = t[244] ^ x[16];
  assign t[204] = t[245] ^ x[19];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[28];
  assign t[208] = t[249] ^ x[31];
  assign t[209] = t[250] ^ x[36];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[39];
  assign t[211] = t[252] ^ x[42];
  assign t[212] = t[253] ^ x[45];
  assign t[213] = t[254] ^ x[48];
  assign t[214] = t[255] ^ x[53];
  assign t[215] = t[256] ^ x[56];
  assign t[216] = t[257] ^ x[59];
  assign t[217] = t[258] ^ x[62];
  assign t[218] = t[259] ^ x[65];
  assign t[219] = t[260] ^ x[68];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[73];
  assign t[221] = t[262] ^ x[76];
  assign t[222] = t[263] ^ x[81];
  assign t[223] = t[264] ^ x[84];
  assign t[224] = t[265] ^ x[87];
  assign t[225] = t[266] ^ x[90];
  assign t[226] = t[267] ^ x[93];
  assign t[227] = t[268] ^ x[98];
  assign t[228] = t[269] ^ x[101];
  assign t[229] = t[270] ^ x[104];
  assign t[22] = ~(t[25] ^ t[34]);
  assign t[230] = t[271] ^ x[109];
  assign t[231] = t[272] ^ x[112];
  assign t[232] = t[273] ^ x[115];
  assign t[233] = t[274] ^ x[118];
  assign t[234] = t[275] ^ x[121];
  assign t[235] = t[276] ^ x[124];
  assign t[236] = t[277] ^ x[127];
  assign t[237] = t[278] ^ x[130];
  assign t[238] = t[279] ^ x[133];
  assign t[239] = t[280] ^ x[136];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[281] ^ x[139];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[8] & x[9]);
  assign t[243] = (x[11] & x[12]);
  assign t[244] = (x[14] & x[15]);
  assign t[245] = (x[17] & x[18]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[26] & x[27]);
  assign t[249] = (x[29] & x[30]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[34] & x[35]);
  assign t[251] = (x[37] & x[38]);
  assign t[252] = (x[40] & x[41]);
  assign t[253] = (x[43] & x[44]);
  assign t[254] = (x[46] & x[47]);
  assign t[255] = (x[51] & x[52]);
  assign t[256] = (x[54] & x[55]);
  assign t[257] = (x[57] & x[58]);
  assign t[258] = (x[60] & x[61]);
  assign t[259] = (x[63] & x[64]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[66] & x[67]);
  assign t[261] = (x[71] & x[72]);
  assign t[262] = (x[74] & x[75]);
  assign t[263] = (x[79] & x[80]);
  assign t[264] = (x[82] & x[83]);
  assign t[265] = (x[85] & x[86]);
  assign t[266] = (x[88] & x[89]);
  assign t[267] = (x[91] & x[92]);
  assign t[268] = (x[96] & x[97]);
  assign t[269] = (x[99] & x[100]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[102] & x[103]);
  assign t[271] = (x[107] & x[108]);
  assign t[272] = (x[110] & x[111]);
  assign t[273] = (x[113] & x[114]);
  assign t[274] = (x[116] & x[117]);
  assign t[275] = (x[119] & x[120]);
  assign t[276] = (x[122] & x[123]);
  assign t[277] = (x[125] & x[126]);
  assign t[278] = (x[128] & x[129]);
  assign t[279] = (x[131] & x[132]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[134] & x[135]);
  assign t[281] = (x[137] & x[138]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[205] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[37] = ~(t[61] | t[62]);
  assign t[38] = ~(t[37] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[206] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[43] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[203]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[78] | t[80]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[204] & t[81];
  assign t[51] = ~(t[82]);
  assign t[52] = ~(t[207]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[83] | t[84]);
  assign t[55] = t[203] ? x[33] : x[32];
  assign t[56] = ~(t[85] & t[86]);
  assign t[57] = ~(t[87] | t[88]);
  assign t[58] = ~(t[209] | t[89]);
  assign t[59] = ~(t[90] | t[91]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[92] ^ t[93]);
  assign t[61] = ~(t[94] | t[95]);
  assign t[62] = ~(t[210] | t[96]);
  assign t[63] = ~(t[97] ^ t[98]);
  assign t[64] = ~(t[211]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[99] | t[100]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[213] | t[103]);
  assign t[69] = t[104] ? x[50] : x[49];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[214] | t[109]);
  assign t[73] = ~(t[110] ^ t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[215] | t[114]);
  assign t[76] = ~(t[115] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119]);
  assign t[79] = t[201] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[201] ? t[123] : t[122];
  assign t[81] = ~(t[119] | t[201]);
  assign t[82] = ~(t[124] | t[125]);
  assign t[83] = ~(t[216]);
  assign t[84] = ~(t[207] | t[208]);
  assign t[85] = ~(t[126] | t[127]);
  assign t[86] = ~(t[128] | t[49]);
  assign t[87] = ~(t[217]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[219] | t[133]);
  assign t[92] = t[104] ? x[70] : x[69];
  assign t[93] = ~(t[134] & t[106]);
  assign t[94] = ~(t[220]);
  assign t[95] = ~(t[221]);
  assign t[96] = ~(t[135] | t[136]);
  assign t[97] = t[203] ? x[78] : x[77];
  assign t[98] = t[137] | t[138];
  assign t[99] = ~(t[222]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind142(x, y);
 input [151:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[32];
  assign t[117] = t[162] ^ x[35];
  assign t[118] = t[163] ^ x[38];
  assign t[119] = t[164] ^ x[41];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[46];
  assign t[121] = t[166] ^ x[51];
  assign t[122] = t[167] ^ x[54];
  assign t[123] = t[168] ^ x[57];
  assign t[124] = t[169] ^ x[60];
  assign t[125] = t[170] ^ x[65];
  assign t[126] = t[171] ^ x[70];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[76];
  assign t[129] = t[174] ^ x[79];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[82];
  assign t[131] = t[176] ^ x[85];
  assign t[132] = t[177] ^ x[88];
  assign t[133] = t[178] ^ x[91];
  assign t[134] = t[179] ^ x[94];
  assign t[135] = t[180] ^ x[97];
  assign t[136] = t[181] ^ x[100];
  assign t[137] = t[182] ^ x[103];
  assign t[138] = t[183] ^ x[106];
  assign t[139] = t[184] ^ x[109];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[112];
  assign t[141] = t[186] ^ x[115];
  assign t[142] = t[187] ^ x[118];
  assign t[143] = t[188] ^ x[121];
  assign t[144] = t[189] ^ x[124];
  assign t[145] = t[190] ^ x[127];
  assign t[146] = t[191] ^ x[130];
  assign t[147] = t[192] ^ x[133];
  assign t[148] = t[193] ^ x[136];
  assign t[149] = t[194] ^ x[139];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[142];
  assign t[151] = t[196] ^ x[145];
  assign t[152] = t[197] ^ x[148];
  assign t[153] = t[198] ^ x[151];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[30] & x[31]);
  assign t[162] = (x[33] & x[34]);
  assign t[163] = (x[36] & x[37]);
  assign t[164] = (x[39] & x[40]);
  assign t[165] = (x[44] & x[45]);
  assign t[166] = (x[49] & x[50]);
  assign t[167] = (x[52] & x[53]);
  assign t[168] = (x[55] & x[56]);
  assign t[169] = (x[58] & x[59]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[63] & x[64]);
  assign t[171] = (x[68] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[74] & x[75]);
  assign t[174] = (x[77] & x[78]);
  assign t[175] = (x[80] & x[81]);
  assign t[176] = (x[83] & x[84]);
  assign t[177] = (x[86] & x[87]);
  assign t[178] = (x[89] & x[90]);
  assign t[179] = (x[92] & x[93]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[95] & x[96]);
  assign t[181] = (x[98] & x[99]);
  assign t[182] = (x[101] & x[102]);
  assign t[183] = (x[104] & x[105]);
  assign t[184] = (x[107] & x[108]);
  assign t[185] = (x[110] & x[111]);
  assign t[186] = (x[113] & x[114]);
  assign t[187] = (x[116] & x[117]);
  assign t[188] = (x[119] & x[120]);
  assign t[189] = (x[122] & x[123]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[125] & x[126]);
  assign t[191] = (x[128] & x[129]);
  assign t[192] = (x[131] & x[132]);
  assign t[193] = (x[134] & x[135]);
  assign t[194] = (x[137] & x[138]);
  assign t[195] = (x[140] & x[141]);
  assign t[196] = (x[143] & x[144]);
  assign t[197] = (x[146] & x[147]);
  assign t[198] = (x[149] & x[150]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[43];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = t[60] | t[115];
  assign t[39] = t[61] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] & t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[71] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[74] | t[118];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[119];
  assign t[53] = t[48] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = t[82] | t[120];
  assign t[57] = t[61] ? x[48] : x[47];
  assign t[58] = ~(t[121]);
  assign t[59] = ~(t[122]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] | t[58]);
  assign t[61] = ~(t[24]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[123];
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = t[89] | t[124];
  assign t[66] = t[61] ? x[62] : x[61];
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = t[92] | t[125];
  assign t[69] = t[61] ? x[67] : x[66];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[93] & t[94]);
  assign t[71] = ~(t[126]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[95] | t[72]);
  assign t[75] = ~(t[129]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[96] | t[75]);
  assign t[78] = ~(t[97] & t[98]);
  assign t[79] = t[99] | t[131];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[132]);
  assign t[81] = ~(t[133]);
  assign t[82] = ~(t[100] | t[80]);
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[101] | t[84]);
  assign t[87] = ~(t[137]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[102] | t[87]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[107] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind143(x, y);
 input [151:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[115] & t[116]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[156]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[155] & t[154]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = t[164] ^ x[2];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[10];
  assign t[121] = t[166] ^ x[13];
  assign t[122] = t[167] ^ x[16];
  assign t[123] = t[168] ^ x[19];
  assign t[124] = t[169] ^ x[22];
  assign t[125] = t[170] ^ x[27];
  assign t[126] = t[171] ^ x[32];
  assign t[127] = t[172] ^ x[35];
  assign t[128] = t[173] ^ x[38];
  assign t[129] = t[174] ^ x[41];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[46];
  assign t[131] = t[176] ^ x[51];
  assign t[132] = t[177] ^ x[54];
  assign t[133] = t[178] ^ x[57];
  assign t[134] = t[179] ^ x[60];
  assign t[135] = t[180] ^ x[65];
  assign t[136] = t[181] ^ x[70];
  assign t[137] = t[182] ^ x[73];
  assign t[138] = t[183] ^ x[76];
  assign t[139] = t[184] ^ x[79];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[82];
  assign t[141] = t[186] ^ x[85];
  assign t[142] = t[187] ^ x[88];
  assign t[143] = t[188] ^ x[91];
  assign t[144] = t[189] ^ x[94];
  assign t[145] = t[190] ^ x[97];
  assign t[146] = t[191] ^ x[100];
  assign t[147] = t[192] ^ x[103];
  assign t[148] = t[193] ^ x[106];
  assign t[149] = t[194] ^ x[109];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[112];
  assign t[151] = t[196] ^ x[115];
  assign t[152] = t[197] ^ x[118];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = t[199] ^ x[124];
  assign t[155] = t[200] ^ x[127];
  assign t[156] = t[201] ^ x[130];
  assign t[157] = t[202] ^ x[133];
  assign t[158] = t[203] ^ x[136];
  assign t[159] = t[204] ^ x[139];
  assign t[15] = ~(t[120] & t[121]);
  assign t[160] = t[205] ^ x[142];
  assign t[161] = t[206] ^ x[145];
  assign t[162] = t[207] ^ x[148];
  assign t[163] = t[208] ^ x[151];
  assign t[164] = (x[0] & x[1]);
  assign t[165] = (x[8] & x[9]);
  assign t[166] = (x[11] & x[12]);
  assign t[167] = (x[14] & x[15]);
  assign t[168] = (x[17] & x[18]);
  assign t[169] = (x[20] & x[21]);
  assign t[16] = ~(t[122] & t[123]);
  assign t[170] = (x[25] & x[26]);
  assign t[171] = (x[30] & x[31]);
  assign t[172] = (x[33] & x[34]);
  assign t[173] = (x[36] & x[37]);
  assign t[174] = (x[39] & x[40]);
  assign t[175] = (x[44] & x[45]);
  assign t[176] = (x[49] & x[50]);
  assign t[177] = (x[52] & x[53]);
  assign t[178] = (x[55] & x[56]);
  assign t[179] = (x[58] & x[59]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[63] & x[64]);
  assign t[181] = (x[68] & x[69]);
  assign t[182] = (x[71] & x[72]);
  assign t[183] = (x[74] & x[75]);
  assign t[184] = (x[77] & x[78]);
  assign t[185] = (x[80] & x[81]);
  assign t[186] = (x[83] & x[84]);
  assign t[187] = (x[86] & x[87]);
  assign t[188] = (x[89] & x[90]);
  assign t[189] = (x[92] & x[93]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[95] & x[96]);
  assign t[191] = (x[98] & x[99]);
  assign t[192] = (x[101] & x[102]);
  assign t[193] = (x[104] & x[105]);
  assign t[194] = (x[107] & x[108]);
  assign t[195] = (x[110] & x[111]);
  assign t[196] = (x[113] & x[114]);
  assign t[197] = (x[116] & x[117]);
  assign t[198] = (x[119] & x[120]);
  assign t[199] = (x[122] & x[123]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[125] & x[126]);
  assign t[201] = (x[128] & x[129]);
  assign t[202] = (x[131] & x[132]);
  assign t[203] = (x[134] & x[135]);
  assign t[204] = (x[137] & x[138]);
  assign t[205] = (x[140] & x[141]);
  assign t[206] = (x[143] & x[144]);
  assign t[207] = (x[146] & x[147]);
  assign t[208] = (x[149] & x[150]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[122]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[124]);
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[43];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = ~(t[60] & t[125]);
  assign t[39] = t[61] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] & t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[126]);
  assign t[46] = ~(t[127]);
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[129]);
  assign t[53] = t[48] ? x[43] : x[42];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = ~(t[81] & t[82]);
  assign t[56] = ~(t[83] & t[130]);
  assign t[57] = t[17] ? x[48] : x[47];
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[132]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[24]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[61] ? x[62] : x[61];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[135]);
  assign t[69] = t[61] ? x[67] : x[66];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[95] & t[96]);
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[101] & t[102]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[103] & t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[104] & t[105]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[110] & t[111]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[119];
endmodule

module R1ind144(x, y);
 input [121:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[25];
  assign t[106] = t[141] ^ x[30];
  assign t[107] = t[142] ^ x[33];
  assign t[108] = t[143] ^ x[38];
  assign t[109] = t[144] ^ x[41];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[44];
  assign t[111] = t[146] ^ x[47];
  assign t[112] = t[147] ^ x[50];
  assign t[113] = t[148] ^ x[55];
  assign t[114] = t[149] ^ x[58];
  assign t[115] = t[150] ^ x[63];
  assign t[116] = t[151] ^ x[66];
  assign t[117] = t[152] ^ x[69];
  assign t[118] = t[153] ^ x[72];
  assign t[119] = t[154] ^ x[75];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[155] ^ x[80];
  assign t[121] = t[156] ^ x[83];
  assign t[122] = t[157] ^ x[88];
  assign t[123] = t[158] ^ x[91];
  assign t[124] = t[159] ^ x[94];
  assign t[125] = t[160] ^ x[97];
  assign t[126] = t[161] ^ x[100];
  assign t[127] = t[162] ^ x[103];
  assign t[128] = t[163] ^ x[106];
  assign t[129] = t[164] ^ x[109];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[112];
  assign t[131] = t[166] ^ x[115];
  assign t[132] = t[167] ^ x[118];
  assign t[133] = t[168] ^ x[121];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[23] & x[24]);
  assign t[141] = (x[28] & x[29]);
  assign t[142] = (x[31] & x[32]);
  assign t[143] = (x[36] & x[37]);
  assign t[144] = (x[39] & x[40]);
  assign t[145] = (x[42] & x[43]);
  assign t[146] = (x[45] & x[46]);
  assign t[147] = (x[48] & x[49]);
  assign t[148] = (x[53] & x[54]);
  assign t[149] = (x[56] & x[57]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[61] & x[62]);
  assign t[151] = (x[64] & x[65]);
  assign t[152] = (x[67] & x[68]);
  assign t[153] = (x[70] & x[71]);
  assign t[154] = (x[73] & x[74]);
  assign t[155] = (x[78] & x[79]);
  assign t[156] = (x[81] & x[82]);
  assign t[157] = (x[86] & x[87]);
  assign t[158] = (x[89] & x[90]);
  assign t[159] = (x[92] & x[93]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[95] & x[96]);
  assign t[161] = (x[98] & x[99]);
  assign t[162] = (x[101] & x[102]);
  assign t[163] = (x[104] & x[105]);
  assign t[164] = (x[107] & x[108]);
  assign t[165] = (x[110] & x[111]);
  assign t[166] = (x[113] & x[114]);
  assign t[167] = (x[116] & x[117]);
  assign t[168] = (x[119] & x[120]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[27] : x[26];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[41];
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = t[59] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[43];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[70]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = t[59] ? x[52] : x[51];
  assign t[53] = ~(t[74] & t[75]);
  assign t[54] = ~(t[113] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = t[47] ? x[60] : x[59];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[24]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[116] & t[79]);
  assign t[61] = ~(t[117] & t[80]);
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = t[59] ? x[77] : x[76];
  assign t[65] = ~(t[83] & t[84]);
  assign t[66] = ~(t[120] & t[85]);
  assign t[67] = ~(t[121] & t[86]);
  assign t[68] = t[59] ? x[85] : x[84];
  assign t[69] = ~(t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[132] & t[97]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[133]);
  assign t[95] = ~(t[133] & t[98]);
  assign t[96] = ~(t[120]);
  assign t[97] = ~(t[124]);
  assign t[98] = ~(t[129]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind145(x, y);
 input [151:0] x;
 output y;

 wire [299:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[143] | t[144]);
  assign t[101] = ~(t[145] | t[146]);
  assign t[102] = ~(t[234] | t[147]);
  assign t[103] = t[90] ? x[87] : x[86];
  assign t[104] = ~(t[148] & t[149]);
  assign t[105] = ~(t[235]);
  assign t[106] = ~(t[222] | t[223]);
  assign t[107] = ~(t[236]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[150] | t[151]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[48]);
  assign t[111] = ~(t[136] | t[152]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[238]);
  assign t[114] = ~(t[239]);
  assign t[115] = ~(t[155] | t[156]);
  assign t[116] = t[110] ? x[104] : x[103];
  assign t[117] = ~(t[157] & t[158]);
  assign t[118] = ~(t[240]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[159] | t[160]);
  assign t[121] = ~(t[161] | t[162]);
  assign t[122] = ~(t[242] | t[163]);
  assign t[123] = t[110] ? x[115] : x[114];
  assign t[124] = ~(t[83] & t[148]);
  assign t[125] = ~(t[213]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(x[4] & t[166]);
  assign t[128] = ~(t[80] | t[167]);
  assign t[129] = ~(t[141] & t[168]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[125] | t[169]);
  assign t[131] = ~(t[125] | t[170]);
  assign t[132] = ~(t[171] & t[214]);
  assign t[133] = ~(t[172] & t[165]);
  assign t[134] = ~(t[243]);
  assign t[135] = ~(t[228] | t[229]);
  assign t[136] = ~(t[80] | t[173]);
  assign t[137] = t[174] | t[175];
  assign t[138] = ~(t[176] & t[177]);
  assign t[139] = ~(t[244]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[230] | t[231]);
  assign t[141] = ~(t[178] | t[179]);
  assign t[142] = ~(t[180] | t[181]);
  assign t[143] = ~(t[245]);
  assign t[144] = ~(t[232] | t[233]);
  assign t[145] = ~(t[246]);
  assign t[146] = ~(t[247]);
  assign t[147] = ~(t[182] | t[183]);
  assign t[148] = ~(t[129] | t[184]);
  assign t[149] = ~(t[128] | t[152]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[248]);
  assign t[151] = ~(t[236] | t[237]);
  assign t[152] = ~(t[80] | t[185]);
  assign t[153] = t[214] & t[186];
  assign t[154] = ~(t[83]);
  assign t[155] = ~(t[249]);
  assign t[156] = ~(t[238] | t[239]);
  assign t[157] = ~(t[178] | t[131]);
  assign t[158] = ~(t[187] | t[175]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[211] & t[212]);
  assign t[160] = ~(t[240] | t[241]);
  assign t[161] = ~(t[251]);
  assign t[162] = ~(t[252]);
  assign t[163] = ~(t[188] | t[189]);
  assign t[164] = ~(x[4] | t[190]);
  assign t[165] = ~(t[214]);
  assign t[166] = ~(t[212] | t[165]);
  assign t[167] = t[211] ? t[132] : t[133];
  assign t[168] = ~(t[125] & t[191]);
  assign t[169] = t[211] ? t[192] : t[133];
  assign t[16] = ~(t[213] & t[214]);
  assign t[170] = t[211] ? t[126] : t[193];
  assign t[171] = x[4] & t[212];
  assign t[172] = ~(x[4] | t[212]);
  assign t[173] = t[211] ? t[193] : t[194];
  assign t[174] = ~(t[83] & t[195]);
  assign t[175] = ~(t[80] | t[196]);
  assign t[176] = ~(t[197] | t[49]);
  assign t[177] = t[125] | t[198];
  assign t[178] = ~(t[125] | t[199]);
  assign t[179] = ~(t[80] | t[200]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[80] | t[201]);
  assign t[181] = ~(t[149] & t[177]);
  assign t[182] = ~(t[253]);
  assign t[183] = ~(t[246] | t[247]);
  assign t[184] = ~(t[202] & t[177]);
  assign t[185] = t[211] ? t[192] : t[203];
  assign t[186] = ~(t[125] | t[211]);
  assign t[187] = ~(t[204]);
  assign t[188] = ~(t[254]);
  assign t[189] = ~(t[251] | t[252]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[212]);
  assign t[191] = ~(t[193] & t[194]);
  assign t[192] = ~(t[171] & t[165]);
  assign t[193] = ~(x[4] & t[205]);
  assign t[194] = ~(t[214] & t[164]);
  assign t[195] = ~(t[166] & t[206]);
  assign t[196] = t[211] ? t[194] : t[193];
  assign t[197] = ~(t[207]);
  assign t[198] = t[211] ? t[193] : t[126];
  assign t[199] = t[211] ? t[133] : t[192];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[211] ? t[126] : t[127];
  assign t[201] = t[211] ? t[203] : t[192];
  assign t[202] = ~(t[153] & t[208]);
  assign t[203] = ~(t[172] & t[214]);
  assign t[204] = ~(t[49] | t[152]);
  assign t[205] = ~(t[212] | t[214]);
  assign t[206] = t[80] & t[211];
  assign t[207] = ~(t[186] & t[209]);
  assign t[208] = t[172] | t[171];
  assign t[209] = ~(t[194] & t[127]);
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[2];
  assign t[211] = t[256] ^ x[10];
  assign t[212] = t[257] ^ x[13];
  assign t[213] = t[258] ^ x[16];
  assign t[214] = t[259] ^ x[19];
  assign t[215] = t[260] ^ x[22];
  assign t[216] = t[261] ^ x[25];
  assign t[217] = t[262] ^ x[28];
  assign t[218] = t[263] ^ x[31];
  assign t[219] = t[264] ^ x[34];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[39];
  assign t[221] = t[266] ^ x[42];
  assign t[222] = t[267] ^ x[45];
  assign t[223] = t[268] ^ x[48];
  assign t[224] = t[269] ^ x[51];
  assign t[225] = t[270] ^ x[56];
  assign t[226] = t[271] ^ x[59];
  assign t[227] = t[272] ^ x[62];
  assign t[228] = t[273] ^ x[65];
  assign t[229] = t[274] ^ x[68];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[71];
  assign t[231] = t[276] ^ x[74];
  assign t[232] = t[277] ^ x[79];
  assign t[233] = t[278] ^ x[82];
  assign t[234] = t[279] ^ x[85];
  assign t[235] = t[280] ^ x[90];
  assign t[236] = t[281] ^ x[93];
  assign t[237] = t[282] ^ x[96];
  assign t[238] = t[283] ^ x[99];
  assign t[239] = t[284] ^ x[102];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[107];
  assign t[241] = t[286] ^ x[110];
  assign t[242] = t[287] ^ x[113];
  assign t[243] = t[288] ^ x[118];
  assign t[244] = t[289] ^ x[121];
  assign t[245] = t[290] ^ x[124];
  assign t[246] = t[291] ^ x[127];
  assign t[247] = t[292] ^ x[130];
  assign t[248] = t[293] ^ x[133];
  assign t[249] = t[294] ^ x[136];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = t[295] ^ x[139];
  assign t[251] = t[296] ^ x[142];
  assign t[252] = t[297] ^ x[145];
  assign t[253] = t[298] ^ x[148];
  assign t[254] = t[299] ^ x[151];
  assign t[255] = (x[0] & x[1]);
  assign t[256] = (x[8] & x[9]);
  assign t[257] = (x[11] & x[12]);
  assign t[258] = (x[14] & x[15]);
  assign t[259] = (x[17] & x[18]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[20] & x[21]);
  assign t[261] = (x[23] & x[24]);
  assign t[262] = (x[26] & x[27]);
  assign t[263] = (x[29] & x[30]);
  assign t[264] = (x[32] & x[33]);
  assign t[265] = (x[37] & x[38]);
  assign t[266] = (x[40] & x[41]);
  assign t[267] = (x[43] & x[44]);
  assign t[268] = (x[46] & x[47]);
  assign t[269] = (x[49] & x[50]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[54] & x[55]);
  assign t[271] = (x[57] & x[58]);
  assign t[272] = (x[60] & x[61]);
  assign t[273] = (x[63] & x[64]);
  assign t[274] = (x[66] & x[67]);
  assign t[275] = (x[69] & x[70]);
  assign t[276] = (x[72] & x[73]);
  assign t[277] = (x[77] & x[78]);
  assign t[278] = (x[80] & x[81]);
  assign t[279] = (x[83] & x[84]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[88] & x[89]);
  assign t[281] = (x[91] & x[92]);
  assign t[282] = (x[94] & x[95]);
  assign t[283] = (x[97] & x[98]);
  assign t[284] = (x[100] & x[101]);
  assign t[285] = (x[105] & x[106]);
  assign t[286] = (x[108] & x[109]);
  assign t[287] = (x[111] & x[112]);
  assign t[288] = (x[116] & x[117]);
  assign t[289] = (x[119] & x[120]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[122] & x[123]);
  assign t[291] = (x[125] & x[126]);
  assign t[292] = (x[128] & x[129]);
  assign t[293] = (x[131] & x[132]);
  assign t[294] = (x[134] & x[135]);
  assign t[295] = (x[137] & x[138]);
  assign t[296] = (x[140] & x[141]);
  assign t[297] = (x[143] & x[144]);
  assign t[298] = (x[146] & x[147]);
  assign t[299] = (x[149] & x[150]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[215] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[46] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[64] ^ t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[66] | t[67]);
  assign t[41] = ~(t[216] | t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[44] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] ^ t[79]);
  assign t[48] = ~(t[213]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = ~(t[80] | t[84]);
  assign t[52] = ~(t[217]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[219] | t[89]);
  assign t[57] = t[90] ? x[36] : x[35];
  assign t[58] = ~(t[91] & t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[220] | t[95]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[221] | t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[103] ^ t[104]);
  assign t[66] = ~(t[222]);
  assign t[67] = ~(t[223]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[224] | t[109]);
  assign t[71] = t[110] ? x[53] : x[52];
  assign t[72] = ~(t[111] & t[112]);
  assign t[73] = ~(t[113] | t[114]);
  assign t[74] = ~(t[225] | t[115]);
  assign t[75] = ~(t[116] ^ t[117]);
  assign t[76] = ~(t[118] | t[119]);
  assign t[77] = ~(t[226] | t[120]);
  assign t[78] = ~(t[121] | t[122]);
  assign t[79] = ~(t[123] ^ t[124]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[125]);
  assign t[81] = t[211] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] | t[131]);
  assign t[84] = t[211] ? t[133] : t[132];
  assign t[85] = ~(t[227]);
  assign t[86] = ~(t[217] | t[218]);
  assign t[87] = ~(t[228]);
  assign t[88] = ~(t[229]);
  assign t[89] = ~(t[134] | t[135]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[48]);
  assign t[91] = ~(t[128] | t[136]);
  assign t[92] = ~(t[137] | t[138]);
  assign t[93] = ~(t[230]);
  assign t[94] = ~(t[231]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = t[90] ? x[76] : x[75];
  assign t[97] = ~(t[141] & t[142]);
  assign t[98] = ~(t[232]);
  assign t[99] = ~(t[233]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[210];
endmodule

module R1ind146(x, y);
 input [106:0] x;
 output y;

 wire [142:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[76];
  assign t[101] = t[133] ^ x[79];
  assign t[102] = t[134] ^ x[82];
  assign t[103] = t[135] ^ x[85];
  assign t[104] = t[136] ^ x[88];
  assign t[105] = t[137] ^ x[91];
  assign t[106] = t[138] ^ x[94];
  assign t[107] = t[139] ^ x[97];
  assign t[108] = t[140] ^ x[100];
  assign t[109] = t[141] ^ x[103];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[106];
  assign t[111] = (x[0] & x[1]);
  assign t[112] = (x[8] & x[9]);
  assign t[113] = (x[11] & x[12]);
  assign t[114] = (x[14] & x[15]);
  assign t[115] = (x[17] & x[18]);
  assign t[116] = (x[20] & x[21]);
  assign t[117] = (x[23] & x[24]);
  assign t[118] = (x[28] & x[29]);
  assign t[119] = (x[31] & x[32]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[34] & x[35]);
  assign t[121] = (x[39] & x[40]);
  assign t[122] = (x[44] & x[45]);
  assign t[123] = (x[47] & x[48]);
  assign t[124] = (x[50] & x[51]);
  assign t[125] = (x[53] & x[54]);
  assign t[126] = (x[56] & x[57]);
  assign t[127] = (x[59] & x[60]);
  assign t[128] = (x[62] & x[63]);
  assign t[129] = (x[65] & x[66]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[68] & x[69]);
  assign t[131] = (x[71] & x[72]);
  assign t[132] = (x[74] & x[75]);
  assign t[133] = (x[77] & x[78]);
  assign t[134] = (x[80] & x[81]);
  assign t[135] = (x[83] & x[84]);
  assign t[136] = (x[86] & x[87]);
  assign t[137] = (x[89] & x[90]);
  assign t[138] = (x[92] & x[93]);
  assign t[139] = (x[95] & x[96]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[98] & x[99]);
  assign t[141] = (x[101] & x[102]);
  assign t[142] = (x[104] & x[105]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[80] & t[81]);
  assign t[16] = ~(t[82] & t[83]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[82]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = t[38] | t[84];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] | t[85];
  assign t[34] = t[17] ? x[27] : x[26];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[86]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[52] | t[36]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[88];
  assign t[41] = t[56] ? x[38] : x[37];
  assign t[42] = ~(t[57] & t[58]);
  assign t[43] = ~(t[59] & t[60]);
  assign t[44] = t[61] | t[89];
  assign t[45] = t[56] ? x[43] : x[42];
  assign t[46] = ~(t[62] & t[63]);
  assign t[47] = ~(t[79]);
  assign t[48] = ~(t[90]);
  assign t[49] = ~(t[64] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[65] & t[66]);
  assign t[51] = t[67] | t[91];
  assign t[52] = ~(t[92]);
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[68] | t[53]);
  assign t[56] = ~(t[23]);
  assign t[57] = ~(t[69] & t[70]);
  assign t[58] = t[71] | t[95];
  assign t[59] = ~(t[96]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[97]);
  assign t[61] = ~(t[72] | t[59]);
  assign t[62] = ~(t[73] & t[74]);
  assign t[63] = t[75] | t[98];
  assign t[64] = ~(t[99]);
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[76] | t[65]);
  assign t[68] = ~(t[102]);
  assign t[69] = ~(t[103]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[77] | t[69]);
  assign t[72] = ~(t[105]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[78] | t[73]);
  assign t[76] = ~(t[108]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = t[111] ^ x[2];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[112] ^ x[10];
  assign t[81] = t[113] ^ x[13];
  assign t[82] = t[114] ^ x[16];
  assign t[83] = t[115] ^ x[19];
  assign t[84] = t[116] ^ x[22];
  assign t[85] = t[117] ^ x[25];
  assign t[86] = t[118] ^ x[30];
  assign t[87] = t[119] ^ x[33];
  assign t[88] = t[120] ^ x[36];
  assign t[89] = t[121] ^ x[41];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[46];
  assign t[91] = t[123] ^ x[49];
  assign t[92] = t[124] ^ x[52];
  assign t[93] = t[125] ^ x[55];
  assign t[94] = t[126] ^ x[58];
  assign t[95] = t[127] ^ x[61];
  assign t[96] = t[128] ^ x[64];
  assign t[97] = t[129] ^ x[67];
  assign t[98] = t[130] ^ x[70];
  assign t[99] = t[131] ^ x[73];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[79];
endmodule

module R1ind147(x, y);
 input [106:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[55];
  assign t[101] = t[133] ^ x[58];
  assign t[102] = t[134] ^ x[61];
  assign t[103] = t[135] ^ x[64];
  assign t[104] = t[136] ^ x[67];
  assign t[105] = t[137] ^ x[70];
  assign t[106] = t[138] ^ x[73];
  assign t[107] = t[139] ^ x[76];
  assign t[108] = t[140] ^ x[79];
  assign t[109] = t[141] ^ x[82];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[85];
  assign t[111] = t[143] ^ x[88];
  assign t[112] = t[144] ^ x[91];
  assign t[113] = t[145] ^ x[94];
  assign t[114] = t[146] ^ x[97];
  assign t[115] = t[147] ^ x[100];
  assign t[116] = t[148] ^ x[103];
  assign t[117] = t[149] ^ x[106];
  assign t[118] = (x[0] & x[1]);
  assign t[119] = (x[8] & x[9]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[11] & x[12]);
  assign t[121] = (x[14] & x[15]);
  assign t[122] = (x[17] & x[18]);
  assign t[123] = (x[20] & x[21]);
  assign t[124] = (x[23] & x[24]);
  assign t[125] = (x[28] & x[29]);
  assign t[126] = (x[31] & x[32]);
  assign t[127] = (x[34] & x[35]);
  assign t[128] = (x[39] & x[40]);
  assign t[129] = (x[44] & x[45]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[47] & x[48]);
  assign t[131] = (x[50] & x[51]);
  assign t[132] = (x[53] & x[54]);
  assign t[133] = (x[56] & x[57]);
  assign t[134] = (x[59] & x[60]);
  assign t[135] = (x[62] & x[63]);
  assign t[136] = (x[65] & x[66]);
  assign t[137] = (x[68] & x[69]);
  assign t[138] = (x[71] & x[72]);
  assign t[139] = (x[74] & x[75]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[77] & x[78]);
  assign t[141] = (x[80] & x[81]);
  assign t[142] = (x[83] & x[84]);
  assign t[143] = (x[86] & x[87]);
  assign t[144] = (x[89] & x[90]);
  assign t[145] = (x[92] & x[93]);
  assign t[146] = (x[95] & x[96]);
  assign t[147] = (x[98] & x[99]);
  assign t[148] = (x[101] & x[102]);
  assign t[149] = (x[104] & x[105]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[87] & t[88]);
  assign t[16] = ~(t[89] & t[90]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[89]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = ~(t[38] & t[91]);
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[92]);
  assign t[34] = t[17] ? x[27] : x[26];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[93]);
  assign t[37] = ~(t[94]);
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[95]);
  assign t[41] = t[57] ? x[38] : x[37];
  assign t[42] = ~(t[58] & t[59]);
  assign t[43] = ~(t[60] & t[61]);
  assign t[44] = ~(t[62] & t[96]);
  assign t[45] = t[57] ? x[43] : x[42];
  assign t[46] = ~(t[63] & t[64]);
  assign t[47] = ~(t[97]);
  assign t[48] = ~(t[98]);
  assign t[49] = ~(t[65] & t[66]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[67] & t[68]);
  assign t[51] = ~(t[69] & t[99]);
  assign t[52] = ~(t[94] & t[93]);
  assign t[53] = ~(t[100]);
  assign t[54] = ~(t[101]);
  assign t[55] = ~(t[102]);
  assign t[56] = ~(t[70] & t[71]);
  assign t[57] = ~(t[23]);
  assign t[58] = ~(t[72] & t[73]);
  assign t[59] = ~(t[74] & t[103]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[104]);
  assign t[61] = ~(t[105]);
  assign t[62] = ~(t[75] & t[76]);
  assign t[63] = ~(t[77] & t[78]);
  assign t[64] = ~(t[79] & t[106]);
  assign t[65] = ~(t[98] & t[97]);
  assign t[66] = ~(t[86]);
  assign t[67] = ~(t[107]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[80] & t[81]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[102] & t[101]);
  assign t[71] = ~(t[109]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[82] & t[83]);
  assign t[75] = ~(t[105] & t[104]);
  assign t[76] = ~(t[112]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[84] & t[85]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[108] & t[107]);
  assign t[81] = ~(t[115]);
  assign t[82] = ~(t[111] & t[110]);
  assign t[83] = ~(t[116]);
  assign t[84] = ~(t[114] & t[113]);
  assign t[85] = ~(t[117]);
  assign t[86] = t[118] ^ x[2];
  assign t[87] = t[119] ^ x[10];
  assign t[88] = t[120] ^ x[13];
  assign t[89] = t[121] ^ x[16];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[19];
  assign t[91] = t[123] ^ x[22];
  assign t[92] = t[124] ^ x[25];
  assign t[93] = t[125] ^ x[30];
  assign t[94] = t[126] ^ x[33];
  assign t[95] = t[127] ^ x[36];
  assign t[96] = t[128] ^ x[41];
  assign t[97] = t[129] ^ x[46];
  assign t[98] = t[130] ^ x[49];
  assign t[99] = t[131] ^ x[52];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[86];
endmodule

module R1ind148(x, y);
 input [88:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[11] & x[12]);
  assign t[101] = (x[14] & x[15]);
  assign t[102] = (x[17] & x[18]);
  assign t[103] = (x[20] & x[21]);
  assign t[104] = (x[23] & x[24]);
  assign t[105] = (x[26] & x[27]);
  assign t[106] = (x[29] & x[30]);
  assign t[107] = (x[34] & x[35]);
  assign t[108] = (x[37] & x[38]);
  assign t[109] = (x[40] & x[41]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[45] & x[46]);
  assign t[111] = (x[48] & x[49]);
  assign t[112] = (x[53] & x[54]);
  assign t[113] = (x[56] & x[57]);
  assign t[114] = (x[59] & x[60]);
  assign t[115] = (x[62] & x[63]);
  assign t[116] = (x[65] & x[66]);
  assign t[117] = (x[68] & x[69]);
  assign t[118] = (x[71] & x[72]);
  assign t[119] = (x[74] & x[75]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[77] & x[78]);
  assign t[121] = (x[80] & x[81]);
  assign t[122] = (x[83] & x[84]);
  assign t[123] = (x[86] & x[87]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[73] & t[74]);
  assign t[16] = ~(t[75] & t[76]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[75]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[77] & t[36]);
  assign t[27] = ~(t[78] & t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[79] & t[46]);
  assign t[33] = ~(t[80] & t[47]);
  assign t[34] = t[17] ? x[33] : x[32];
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[81]);
  assign t[37] = ~(t[81] & t[50]);
  assign t[38] = ~(t[82] & t[51]);
  assign t[39] = ~(t[83] & t[52]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[53] ? x[44] : x[43];
  assign t[41] = ~(t[54] & t[55]);
  assign t[42] = ~(t[84] & t[56]);
  assign t[43] = ~(t[85] & t[57]);
  assign t[44] = t[53] ? x[52] : x[51];
  assign t[45] = ~(t[58] & t[59]);
  assign t[46] = ~(t[86]);
  assign t[47] = ~(t[86] & t[60]);
  assign t[48] = ~(t[87] & t[61]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[77]);
  assign t[51] = ~(t[89]);
  assign t[52] = ~(t[89] & t[63]);
  assign t[53] = ~(t[23]);
  assign t[54] = ~(t[90] & t[64]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92]);
  assign t[57] = ~(t[92] & t[66]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[79]);
  assign t[61] = ~(t[95]);
  assign t[62] = ~(t[95] & t[69]);
  assign t[63] = ~(t[82]);
  assign t[64] = ~(t[96]);
  assign t[65] = ~(t[96] & t[70]);
  assign t[66] = ~(t[84]);
  assign t[67] = ~(t[97]);
  assign t[68] = ~(t[97] & t[71]);
  assign t[69] = ~(t[87]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[90]);
  assign t[71] = ~(t[93]);
  assign t[72] = t[98] ^ x[2];
  assign t[73] = t[99] ^ x[10];
  assign t[74] = t[100] ^ x[13];
  assign t[75] = t[101] ^ x[16];
  assign t[76] = t[102] ^ x[19];
  assign t[77] = t[103] ^ x[22];
  assign t[78] = t[104] ^ x[25];
  assign t[79] = t[105] ^ x[28];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] ^ x[31];
  assign t[81] = t[107] ^ x[36];
  assign t[82] = t[108] ^ x[39];
  assign t[83] = t[109] ^ x[42];
  assign t[84] = t[110] ^ x[47];
  assign t[85] = t[111] ^ x[50];
  assign t[86] = t[112] ^ x[55];
  assign t[87] = t[113] ^ x[58];
  assign t[88] = t[114] ^ x[61];
  assign t[89] = t[115] ^ x[64];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[116] ^ x[67];
  assign t[91] = t[117] ^ x[70];
  assign t[92] = t[118] ^ x[73];
  assign t[93] = t[119] ^ x[76];
  assign t[94] = t[120] ^ x[79];
  assign t[95] = t[121] ^ x[82];
  assign t[96] = t[122] ^ x[85];
  assign t[97] = t[123] ^ x[88];
  assign t[98] = (x[0] & x[1]);
  assign t[99] = (x[8] & x[9]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[72];
endmodule

module R1ind149(x, y);
 input [106:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[176]);
  assign t[101] = ~(t[119] | t[120]);
  assign t[102] = ~(t[39]);
  assign t[103] = ~(t[121] | t[122]);
  assign t[104] = ~(t[123] & t[124]);
  assign t[105] = ~(t[177]);
  assign t[106] = ~(t[169] | t[170]);
  assign t[107] = ~(t[178]);
  assign t[108] = ~(t[179]);
  assign t[109] = ~(t[125] | t[126]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[113] | t[127]);
  assign t[111] = ~(t[180]);
  assign t[112] = ~(t[172] | t[173]);
  assign t[113] = ~(t[42] | t[128]);
  assign t[114] = ~(t[129]);
  assign t[115] = ~(t[130] & t[94]);
  assign t[116] = ~(t[131] & t[94]);
  assign t[117] = ~(t[96] & t[94]);
  assign t[118] = ~(t[153]);
  assign t[119] = ~(t[181]);
  assign t[11] = ~(t[17] ^ t[14]);
  assign t[120] = ~(t[175] | t[176]);
  assign t[121] = ~(t[132] & t[41]);
  assign t[122] = t[28] | t[133];
  assign t[123] = t[155] & t[134];
  assign t[124] = t[130] | t[131];
  assign t[125] = ~(t[182]);
  assign t[126] = ~(t[178] | t[179]);
  assign t[127] = ~(t[135] & t[136]);
  assign t[128] = t[152] ? t[137] : t[115];
  assign t[129] = ~(t[138] | t[139]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(x[4] | t[153]);
  assign t[131] = x[4] & t[153];
  assign t[132] = ~(t[134] & t[140]);
  assign t[133] = ~(t[42] | t[141]);
  assign t[134] = ~(t[66] | t[152]);
  assign t[135] = ~(t[142] | t[143]);
  assign t[136] = ~(t[66] & t[144]);
  assign t[137] = ~(t[131] & t[155]);
  assign t[138] = ~(t[42] | t[145]);
  assign t[139] = ~(t[42] | t[146]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = ~(t[68] & t[147]);
  assign t[141] = t[152] ? t[148] : t[116];
  assign t[142] = ~(t[66] | t[149]);
  assign t[143] = ~(t[42] | t[150]);
  assign t[144] = ~(t[67] & t[68]);
  assign t[145] = t[152] ? t[147] : t[117];
  assign t[146] = t[152] ? t[116] : t[148];
  assign t[147] = ~(x[4] & t[64]);
  assign t[148] = ~(t[130] & t[155]);
  assign t[149] = t[152] ? t[115] : t[116];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[152] ? t[117] : t[147];
  assign t[151] = t[183] ^ x[2];
  assign t[152] = t[184] ^ x[10];
  assign t[153] = t[185] ^ x[13];
  assign t[154] = t[186] ^ x[16];
  assign t[155] = t[187] ^ x[19];
  assign t[156] = t[188] ^ x[22];
  assign t[157] = t[189] ^ x[25];
  assign t[158] = t[190] ^ x[28];
  assign t[159] = t[191] ^ x[31];
  assign t[15] = ~(t[152] & t[153]);
  assign t[160] = t[192] ^ x[34];
  assign t[161] = t[193] ^ x[37];
  assign t[162] = t[194] ^ x[40];
  assign t[163] = t[195] ^ x[43];
  assign t[164] = t[196] ^ x[46];
  assign t[165] = t[197] ^ x[51];
  assign t[166] = t[198] ^ x[54];
  assign t[167] = t[199] ^ x[57];
  assign t[168] = t[200] ^ x[60];
  assign t[169] = t[201] ^ x[65];
  assign t[16] = ~(t[154] & t[155]);
  assign t[170] = t[202] ^ x[68];
  assign t[171] = t[203] ^ x[71];
  assign t[172] = t[204] ^ x[76];
  assign t[173] = t[205] ^ x[79];
  assign t[174] = t[206] ^ x[82];
  assign t[175] = t[207] ^ x[85];
  assign t[176] = t[208] ^ x[88];
  assign t[177] = t[209] ^ x[91];
  assign t[178] = t[210] ^ x[94];
  assign t[179] = t[211] ^ x[97];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[212] ^ x[100];
  assign t[181] = t[213] ^ x[103];
  assign t[182] = t[214] ^ x[106];
  assign t[183] = (x[0] & x[1]);
  assign t[184] = (x[8] & x[9]);
  assign t[185] = (x[11] & x[12]);
  assign t[186] = (x[14] & x[15]);
  assign t[187] = (x[17] & x[18]);
  assign t[188] = (x[20] & x[21]);
  assign t[189] = (x[23] & x[24]);
  assign t[18] = t[26] ? x[7] : x[6];
  assign t[190] = (x[26] & x[27]);
  assign t[191] = (x[29] & x[30]);
  assign t[192] = (x[32] & x[33]);
  assign t[193] = (x[35] & x[36]);
  assign t[194] = (x[38] & x[39]);
  assign t[195] = (x[41] & x[42]);
  assign t[196] = (x[44] & x[45]);
  assign t[197] = (x[49] & x[50]);
  assign t[198] = (x[52] & x[53]);
  assign t[199] = (x[55] & x[56]);
  assign t[19] = t[27] | t[28];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[58] & x[59]);
  assign t[201] = (x[63] & x[64]);
  assign t[202] = (x[66] & x[67]);
  assign t[203] = (x[69] & x[70]);
  assign t[204] = (x[74] & x[75]);
  assign t[205] = (x[77] & x[78]);
  assign t[206] = (x[80] & x[81]);
  assign t[207] = (x[83] & x[84]);
  assign t[208] = (x[86] & x[87]);
  assign t[209] = (x[89] & x[90]);
  assign t[20] = ~(t[29] | t[30]);
  assign t[210] = (x[92] & x[93]);
  assign t[211] = (x[95] & x[96]);
  assign t[212] = (x[98] & x[99]);
  assign t[213] = (x[101] & x[102]);
  assign t[214] = (x[104] & x[105]);
  assign t[21] = ~(t[24] ^ t[12]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[40] & t[41]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[29] = ~(t[44] | t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[156] | t[46]);
  assign t[31] = ~(t[47] | t[48]);
  assign t[32] = ~(t[49] ^ t[50]);
  assign t[33] = ~(t[51] | t[52]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[157] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] ^ t[61]);
  assign t[39] = ~(t[154]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] | t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = ~(t[66]);
  assign t[43] = t[152] ? t[68] : t[67];
  assign t[44] = ~(t[158]);
  assign t[45] = ~(t[159]);
  assign t[46] = ~(t[69] | t[70]);
  assign t[47] = ~(t[71] | t[72]);
  assign t[48] = ~(t[160] | t[73]);
  assign t[49] = ~(t[74] | t[75]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[76] ^ t[77]);
  assign t[51] = ~(t[78] | t[79]);
  assign t[52] = ~(t[161] | t[80]);
  assign t[53] = ~(t[81] | t[82]);
  assign t[54] = ~(t[83] ^ t[84]);
  assign t[55] = ~(t[162]);
  assign t[56] = ~(t[163]);
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[87] | t[88]);
  assign t[59] = ~(t[164] | t[89]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[26] ? x[48] : x[47];
  assign t[61] = ~(t[90] & t[91]);
  assign t[62] = ~(t[66] | t[92]);
  assign t[63] = ~(t[66] | t[93]);
  assign t[64] = ~(t[153] | t[94]);
  assign t[65] = t[42] & t[152];
  assign t[66] = ~(t[154]);
  assign t[67] = ~(x[4] & t[95]);
  assign t[68] = ~(t[155] & t[96]);
  assign t[69] = ~(t[165]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[158] | t[159]);
  assign t[71] = ~(t[166]);
  assign t[72] = ~(t[167]);
  assign t[73] = ~(t[97] | t[98]);
  assign t[74] = ~(t[99] | t[100]);
  assign t[75] = ~(t[168] | t[101]);
  assign t[76] = t[102] ? x[62] : x[61];
  assign t[77] = ~(t[103] & t[104]);
  assign t[78] = ~(t[169]);
  assign t[79] = ~(t[170]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[105] | t[106]);
  assign t[81] = ~(t[107] | t[108]);
  assign t[82] = ~(t[171] | t[109]);
  assign t[83] = t[102] ? x[73] : x[72];
  assign t[84] = ~(t[110] & t[41]);
  assign t[85] = ~(t[151]);
  assign t[86] = ~(t[162] | t[163]);
  assign t[87] = ~(t[172]);
  assign t[88] = ~(t[173]);
  assign t[89] = ~(t[111] | t[112]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[113]);
  assign t[91] = ~(t[114] | t[28]);
  assign t[92] = t[152] ? t[116] : t[115];
  assign t[93] = t[152] ? t[117] : t[67];
  assign t[94] = ~(t[155]);
  assign t[95] = ~(t[153] | t[155]);
  assign t[96] = ~(x[4] | t[118]);
  assign t[97] = ~(t[174]);
  assign t[98] = ~(t[166] | t[167]);
  assign t[99] = ~(t[175]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[151];
endmodule

module R1ind150(x, y);
 input [151:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[107] | t[100]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[32];
  assign t[117] = t[162] ^ x[35];
  assign t[118] = t[163] ^ x[38];
  assign t[119] = t[164] ^ x[41];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[46];
  assign t[121] = t[166] ^ x[51];
  assign t[122] = t[167] ^ x[54];
  assign t[123] = t[168] ^ x[57];
  assign t[124] = t[169] ^ x[60];
  assign t[125] = t[170] ^ x[65];
  assign t[126] = t[171] ^ x[70];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[76];
  assign t[129] = t[174] ^ x[79];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[82];
  assign t[131] = t[176] ^ x[85];
  assign t[132] = t[177] ^ x[88];
  assign t[133] = t[178] ^ x[91];
  assign t[134] = t[179] ^ x[94];
  assign t[135] = t[180] ^ x[97];
  assign t[136] = t[181] ^ x[100];
  assign t[137] = t[182] ^ x[103];
  assign t[138] = t[183] ^ x[106];
  assign t[139] = t[184] ^ x[109];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[112];
  assign t[141] = t[186] ^ x[115];
  assign t[142] = t[187] ^ x[118];
  assign t[143] = t[188] ^ x[121];
  assign t[144] = t[189] ^ x[124];
  assign t[145] = t[190] ^ x[127];
  assign t[146] = t[191] ^ x[130];
  assign t[147] = t[192] ^ x[133];
  assign t[148] = t[193] ^ x[136];
  assign t[149] = t[194] ^ x[139];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[142];
  assign t[151] = t[196] ^ x[145];
  assign t[152] = t[197] ^ x[148];
  assign t[153] = t[198] ^ x[151];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[30] & x[31]);
  assign t[162] = (x[33] & x[34]);
  assign t[163] = (x[36] & x[37]);
  assign t[164] = (x[39] & x[40]);
  assign t[165] = (x[44] & x[45]);
  assign t[166] = (x[49] & x[50]);
  assign t[167] = (x[52] & x[53]);
  assign t[168] = (x[55] & x[56]);
  assign t[169] = (x[58] & x[59]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[63] & x[64]);
  assign t[171] = (x[68] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[74] & x[75]);
  assign t[174] = (x[77] & x[78]);
  assign t[175] = (x[80] & x[81]);
  assign t[176] = (x[83] & x[84]);
  assign t[177] = (x[86] & x[87]);
  assign t[178] = (x[89] & x[90]);
  assign t[179] = (x[92] & x[93]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[95] & x[96]);
  assign t[181] = (x[98] & x[99]);
  assign t[182] = (x[101] & x[102]);
  assign t[183] = (x[104] & x[105]);
  assign t[184] = (x[107] & x[108]);
  assign t[185] = (x[110] & x[111]);
  assign t[186] = (x[113] & x[114]);
  assign t[187] = (x[116] & x[117]);
  assign t[188] = (x[119] & x[120]);
  assign t[189] = (x[122] & x[123]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[125] & x[126]);
  assign t[191] = (x[128] & x[129]);
  assign t[192] = (x[131] & x[132]);
  assign t[193] = (x[134] & x[135]);
  assign t[194] = (x[137] & x[138]);
  assign t[195] = (x[140] & x[141]);
  assign t[196] = (x[143] & x[144]);
  assign t[197] = (x[146] & x[147]);
  assign t[198] = (x[149] & x[150]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[41];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[69] | t[45]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = t[72] | t[118];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = t[75] | t[119];
  assign t[52] = t[76] ? x[43] : x[42];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = t[79] | t[120];
  assign t[55] = t[76] ? x[48] : x[47];
  assign t[56] = ~(t[121]);
  assign t[57] = ~(t[122]);
  assign t[58] = ~(t[80] | t[56]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[83] | t[123];
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = t[86] | t[124];
  assign t[63] = t[87] ? x[62] : x[61];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = t[92] | t[125];
  assign t[67] = t[87] ? x[67] : x[66];
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = ~(t[126]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[95] | t[70]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[96] | t[73]);
  assign t[76] = ~(t[24]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[97] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[24]);
  assign t[88] = ~(t[100] & t[101]);
  assign t[89] = t[102] | t[138];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind151(x, y);
 input [151:0] x;
 output y;

 wire [206:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[143] & t[142]);
  assign t[102] = ~(t[153]);
  assign t[103] = ~(t[145] & t[144]);
  assign t[104] = ~(t[154]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[113] & t[114]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[157]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[115] & t[116]);
  assign t[113] = ~(t[156] & t[155]);
  assign t[114] = ~(t[160]);
  assign t[115] = ~(t[159] & t[158]);
  assign t[116] = ~(t[161]);
  assign t[117] = t[162] ^ x[2];
  assign t[118] = t[163] ^ x[8];
  assign t[119] = t[164] ^ x[11];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[165] ^ x[14];
  assign t[121] = t[166] ^ x[17];
  assign t[122] = t[167] ^ x[22];
  assign t[123] = t[168] ^ x[27];
  assign t[124] = t[169] ^ x[32];
  assign t[125] = t[170] ^ x[35];
  assign t[126] = t[171] ^ x[38];
  assign t[127] = t[172] ^ x[41];
  assign t[128] = t[173] ^ x[46];
  assign t[129] = t[174] ^ x[51];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[54];
  assign t[131] = t[176] ^ x[57];
  assign t[132] = t[177] ^ x[60];
  assign t[133] = t[178] ^ x[65];
  assign t[134] = t[179] ^ x[70];
  assign t[135] = t[180] ^ x[73];
  assign t[136] = t[181] ^ x[76];
  assign t[137] = t[182] ^ x[79];
  assign t[138] = t[183] ^ x[82];
  assign t[139] = t[184] ^ x[85];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[88];
  assign t[141] = t[186] ^ x[91];
  assign t[142] = t[187] ^ x[94];
  assign t[143] = t[188] ^ x[97];
  assign t[144] = t[189] ^ x[100];
  assign t[145] = t[190] ^ x[103];
  assign t[146] = t[191] ^ x[106];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[112];
  assign t[149] = t[194] ^ x[115];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[118];
  assign t[151] = t[196] ^ x[121];
  assign t[152] = t[197] ^ x[124];
  assign t[153] = t[198] ^ x[127];
  assign t[154] = t[199] ^ x[130];
  assign t[155] = t[200] ^ x[133];
  assign t[156] = t[201] ^ x[136];
  assign t[157] = t[202] ^ x[139];
  assign t[158] = t[203] ^ x[142];
  assign t[159] = t[204] ^ x[145];
  assign t[15] = ~(t[22]);
  assign t[160] = t[205] ^ x[148];
  assign t[161] = t[206] ^ x[151];
  assign t[162] = (x[0] & x[1]);
  assign t[163] = (x[6] & x[7]);
  assign t[164] = (x[9] & x[10]);
  assign t[165] = (x[12] & x[13]);
  assign t[166] = (x[15] & x[16]);
  assign t[167] = (x[20] & x[21]);
  assign t[168] = (x[25] & x[26]);
  assign t[169] = (x[30] & x[31]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[33] & x[34]);
  assign t[171] = (x[36] & x[37]);
  assign t[172] = (x[39] & x[40]);
  assign t[173] = (x[44] & x[45]);
  assign t[174] = (x[49] & x[50]);
  assign t[175] = (x[52] & x[53]);
  assign t[176] = (x[55] & x[56]);
  assign t[177] = (x[58] & x[59]);
  assign t[178] = (x[63] & x[64]);
  assign t[179] = (x[68] & x[69]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[71] & x[72]);
  assign t[181] = (x[74] & x[75]);
  assign t[182] = (x[77] & x[78]);
  assign t[183] = (x[80] & x[81]);
  assign t[184] = (x[83] & x[84]);
  assign t[185] = (x[86] & x[87]);
  assign t[186] = (x[89] & x[90]);
  assign t[187] = (x[92] & x[93]);
  assign t[188] = (x[95] & x[96]);
  assign t[189] = (x[98] & x[99]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[101] & x[102]);
  assign t[191] = (x[104] & x[105]);
  assign t[192] = (x[107] & x[108]);
  assign t[193] = (x[110] & x[111]);
  assign t[194] = (x[113] & x[114]);
  assign t[195] = (x[116] & x[117]);
  assign t[196] = (x[119] & x[120]);
  assign t[197] = (x[122] & x[123]);
  assign t[198] = (x[125] & x[126]);
  assign t[199] = (x[128] & x[129]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = (x[131] & x[132]);
  assign t[201] = (x[134] & x[135]);
  assign t[202] = (x[137] & x[138]);
  assign t[203] = (x[140] & x[141]);
  assign t[204] = (x[143] & x[144]);
  assign t[205] = (x[146] & x[147]);
  assign t[206] = (x[149] & x[150]);
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[120]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = ~(t[45] & t[122]);
  assign t[29] = t[15] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[31];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[39];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = ~(t[56] & t[123]);
  assign t[37] = t[15] ? x[29] : x[28];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[124]);
  assign t[44] = ~(t[125]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[126]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[74] & t[127]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[75] ? x[43] : x[42];
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[128]);
  assign t[53] = t[75] ? x[48] : x[47];
  assign t[54] = ~(t[129]);
  assign t[55] = ~(t[130]);
  assign t[56] = ~(t[79] & t[80]);
  assign t[57] = ~(t[81] & t[82]);
  assign t[58] = ~(t[83] & t[131]);
  assign t[59] = ~(t[84] & t[85]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[86] & t[132]);
  assign t[61] = t[87] ? x[62] : x[61];
  assign t[62] = ~(t[88] & t[89]);
  assign t[63] = ~(t[90] & t[91]);
  assign t[64] = ~(t[92] & t[133]);
  assign t[65] = t[87] ? x[67] : x[66];
  assign t[66] = ~(t[93] & t[94]);
  assign t[67] = ~(t[125] & t[124]);
  assign t[68] = ~(t[134]);
  assign t[69] = ~(t[135]);
  assign t[6] = ~(t[118] & t[119]);
  assign t[70] = ~(t[136]);
  assign t[71] = ~(t[95] & t[96]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[97] & t[98]);
  assign t[75] = ~(t[22]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[130] & t[129]);
  assign t[7] = ~(t[120] & t[121]);
  assign t[80] = ~(t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[101] & t[102]);
  assign t[84] = ~(t[144]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[103] & t[104]);
  assign t[87] = ~(t[22]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[146]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[147]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[108] & t[109]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[112] & t[149]);
  assign t[95] = ~(t[136] & t[135]);
  assign t[96] = ~(t[150]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[151]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[117];
endmodule

module R1ind152(x, y);
 input [121:0] x;
 output y;

 wire [166:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[135] ^ x[14];
  assign t[101] = t[136] ^ x[17];
  assign t[102] = t[137] ^ x[22];
  assign t[103] = t[138] ^ x[25];
  assign t[104] = t[139] ^ x[30];
  assign t[105] = t[140] ^ x[33];
  assign t[106] = t[141] ^ x[38];
  assign t[107] = t[142] ^ x[41];
  assign t[108] = t[143] ^ x[44];
  assign t[109] = t[144] ^ x[47];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[145] ^ x[50];
  assign t[111] = t[146] ^ x[55];
  assign t[112] = t[147] ^ x[58];
  assign t[113] = t[148] ^ x[63];
  assign t[114] = t[149] ^ x[66];
  assign t[115] = t[150] ^ x[69];
  assign t[116] = t[151] ^ x[72];
  assign t[117] = t[152] ^ x[75];
  assign t[118] = t[153] ^ x[80];
  assign t[119] = t[154] ^ x[83];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[155] ^ x[88];
  assign t[121] = t[156] ^ x[91];
  assign t[122] = t[157] ^ x[94];
  assign t[123] = t[158] ^ x[97];
  assign t[124] = t[159] ^ x[100];
  assign t[125] = t[160] ^ x[103];
  assign t[126] = t[161] ^ x[106];
  assign t[127] = t[162] ^ x[109];
  assign t[128] = t[163] ^ x[112];
  assign t[129] = t[164] ^ x[115];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[165] ^ x[118];
  assign t[131] = t[166] ^ x[121];
  assign t[132] = (x[0] & x[1]);
  assign t[133] = (x[6] & x[7]);
  assign t[134] = (x[9] & x[10]);
  assign t[135] = (x[12] & x[13]);
  assign t[136] = (x[15] & x[16]);
  assign t[137] = (x[20] & x[21]);
  assign t[138] = (x[23] & x[24]);
  assign t[139] = (x[28] & x[29]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[31] & x[32]);
  assign t[141] = (x[36] & x[37]);
  assign t[142] = (x[39] & x[40]);
  assign t[143] = (x[42] & x[43]);
  assign t[144] = (x[45] & x[46]);
  assign t[145] = (x[48] & x[49]);
  assign t[146] = (x[53] & x[54]);
  assign t[147] = (x[56] & x[57]);
  assign t[148] = (x[61] & x[62]);
  assign t[149] = (x[64] & x[65]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (x[67] & x[68]);
  assign t[151] = (x[70] & x[71]);
  assign t[152] = (x[73] & x[74]);
  assign t[153] = (x[78] & x[79]);
  assign t[154] = (x[81] & x[82]);
  assign t[155] = (x[86] & x[87]);
  assign t[156] = (x[89] & x[90]);
  assign t[157] = (x[92] & x[93]);
  assign t[158] = (x[95] & x[96]);
  assign t[159] = (x[98] & x[99]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[101] & x[102]);
  assign t[161] = (x[104] & x[105]);
  assign t[162] = (x[107] & x[108]);
  assign t[163] = (x[110] & x[111]);
  assign t[164] = (x[113] & x[114]);
  assign t[165] = (x[116] & x[117]);
  assign t[166] = (x[119] & x[120]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[100]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[102] & t[43]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[29] = t[15] ? x[27] : x[26];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[32] = t[49] ^ t[39];
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[104] & t[53]);
  assign t[36] = ~(t[105] & t[54]);
  assign t[37] = t[15] ? x[35] : x[34];
  assign t[38] = ~(t[55] & t[56]);
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[59] ^ t[60];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[106]);
  assign t[44] = ~(t[106] & t[65]);
  assign t[45] = ~(t[107] & t[66]);
  assign t[46] = ~(t[108] & t[67]);
  assign t[47] = ~(t[109] & t[68]);
  assign t[48] = ~(t[110] & t[69]);
  assign t[49] = t[70] ? x[52] : x[51];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[70] ? x[60] : x[59];
  assign t[53] = ~(t[113]);
  assign t[54] = ~(t[113] & t[73]);
  assign t[55] = ~(t[114] & t[74]);
  assign t[56] = ~(t[115] & t[75]);
  assign t[57] = ~(t[116] & t[76]);
  assign t[58] = ~(t[117] & t[77]);
  assign t[59] = t[78] ? x[77] : x[76];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[79] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[78] ? x[85] : x[84];
  assign t[64] = ~(t[83] & t[84]);
  assign t[65] = ~(t[102]);
  assign t[66] = ~(t[120]);
  assign t[67] = ~(t[120] & t[85]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = ~(t[98] & t[99]);
  assign t[70] = ~(t[22]);
  assign t[71] = ~(t[122]);
  assign t[72] = ~(t[122] & t[87]);
  assign t[73] = ~(t[104]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[123] & t[88]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[124] & t[89]);
  assign t[78] = ~(t[22]);
  assign t[79] = ~(t[125] & t[90]);
  assign t[7] = ~(t[100] & t[101]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[127] & t[92]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[114]);
  assign t[89] = ~(t[116]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[130]);
  assign t[91] = ~(t[130] & t[95]);
  assign t[92] = ~(t[118]);
  assign t[93] = ~(t[131]);
  assign t[94] = ~(t[131] & t[96]);
  assign t[95] = ~(t[125]);
  assign t[96] = ~(t[128]);
  assign t[97] = t[132] ^ x[2];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[11];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[97];
endmodule

module R1ind153(x, y);
 input [151:0] x;
 output y;

 wire [289:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[138] & t[139]);
  assign t[101] = ~(t[224]);
  assign t[102] = ~(t[212] | t[213]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[140] | t[141]);
  assign t[106] = ~(t[138] & t[142]);
  assign t[107] = ~(t[227]);
  assign t[108] = ~(t[228]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[145] | t[146]);
  assign t[111] = ~(t[229] | t[147]);
  assign t[112] = t[148] ? x[104] : x[103];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[230]);
  assign t[115] = ~(t[231]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[232] | t[155]);
  assign t[119] = t[148] ? x[115] : x[114];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[156] & t[142]);
  assign t[121] = ~(t[203]);
  assign t[122] = ~(t[157] & t[158]);
  assign t[123] = ~(t[159] & t[204]);
  assign t[124] = ~(t[80] | t[160]);
  assign t[125] = ~(t[80] | t[161]);
  assign t[126] = ~(x[4] & t[162]);
  assign t[127] = ~(t[204] & t[163]);
  assign t[128] = ~(t[233]);
  assign t[129] = ~(t[218] | t[219]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[156] & t[138]);
  assign t[131] = ~(t[80] | t[164]);
  assign t[132] = ~(t[234]);
  assign t[133] = ~(t[220] | t[221]);
  assign t[134] = ~(t[48]);
  assign t[135] = ~(t[165] | t[166]);
  assign t[136] = ~(t[235]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[167] | t[166]);
  assign t[139] = ~(t[168] | t[169]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[236]);
  assign t[141] = ~(t[225] | t[226]);
  assign t[142] = ~(t[170] & t[171]);
  assign t[143] = ~(t[237]);
  assign t[144] = ~(t[227] | t[228]);
  assign t[145] = ~(t[238]);
  assign t[146] = ~(t[239]);
  assign t[147] = ~(t[172] | t[173]);
  assign t[148] = ~(t[48]);
  assign t[149] = ~(t[174] | t[175]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[176] & t[177]);
  assign t[151] = ~(t[240]);
  assign t[152] = ~(t[230] | t[231]);
  assign t[153] = ~(t[241]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[178] | t[179]);
  assign t[156] = ~(t[49] | t[168]);
  assign t[157] = ~(x[4] | t[202]);
  assign t[158] = ~(t[204]);
  assign t[159] = x[4] & t[202];
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = t[201] ? t[181] : t[180];
  assign t[161] = t[201] ? t[183] : t[182];
  assign t[162] = ~(t[202] | t[204]);
  assign t[163] = ~(x[4] | t[184]);
  assign t[164] = t[201] ? t[122] : t[123];
  assign t[165] = ~(t[121] | t[185]);
  assign t[166] = ~(t[121] | t[186]);
  assign t[167] = ~(t[121] | t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[150] & t[190]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[202] | t[158]);
  assign t[171] = t[80] & t[201];
  assign t[172] = ~(t[243]);
  assign t[173] = ~(t[238] | t[239]);
  assign t[174] = ~(t[191] & t[142]);
  assign t[175] = t[51] | t[192];
  assign t[176] = t[204] & t[193];
  assign t[177] = t[157] | t[159];
  assign t[178] = ~(t[244]);
  assign t[179] = ~(t[241] | t[242]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[163] & t[158]);
  assign t[181] = ~(x[4] & t[170]);
  assign t[182] = ~(t[157] & t[204]);
  assign t[183] = ~(t[159] & t[158]);
  assign t[184] = ~(t[202]);
  assign t[185] = t[201] ? t[122] : t[183];
  assign t[186] = t[201] ? t[180] : t[126];
  assign t[187] = t[201] ? t[183] : t[122];
  assign t[188] = ~(t[165] | t[194]);
  assign t[189] = ~(t[121] & t[195]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[121] | t[196];
  assign t[191] = ~(t[193] & t[197]);
  assign t[192] = ~(t[80] | t[198]);
  assign t[193] = ~(t[121] | t[201]);
  assign t[194] = ~(t[80] | t[199]);
  assign t[195] = ~(t[126] & t[127]);
  assign t[196] = t[201] ? t[126] : t[180];
  assign t[197] = ~(t[127] & t[181]);
  assign t[198] = t[201] ? t[182] : t[183];
  assign t[199] = t[201] ? t[180] : t[181];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[245] ^ x[2];
  assign t[201] = t[246] ^ x[10];
  assign t[202] = t[247] ^ x[13];
  assign t[203] = t[248] ^ x[16];
  assign t[204] = t[249] ^ x[19];
  assign t[205] = t[250] ^ x[22];
  assign t[206] = t[251] ^ x[25];
  assign t[207] = t[252] ^ x[28];
  assign t[208] = t[253] ^ x[31];
  assign t[209] = t[254] ^ x[34];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[39];
  assign t[211] = t[256] ^ x[42];
  assign t[212] = t[257] ^ x[45];
  assign t[213] = t[258] ^ x[48];
  assign t[214] = t[259] ^ x[51];
  assign t[215] = t[260] ^ x[56];
  assign t[216] = t[261] ^ x[59];
  assign t[217] = t[262] ^ x[62];
  assign t[218] = t[263] ^ x[65];
  assign t[219] = t[264] ^ x[68];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[71];
  assign t[221] = t[266] ^ x[74];
  assign t[222] = t[267] ^ x[79];
  assign t[223] = t[268] ^ x[82];
  assign t[224] = t[269] ^ x[87];
  assign t[225] = t[270] ^ x[90];
  assign t[226] = t[271] ^ x[93];
  assign t[227] = t[272] ^ x[96];
  assign t[228] = t[273] ^ x[99];
  assign t[229] = t[274] ^ x[102];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[107];
  assign t[231] = t[276] ^ x[110];
  assign t[232] = t[277] ^ x[113];
  assign t[233] = t[278] ^ x[118];
  assign t[234] = t[279] ^ x[121];
  assign t[235] = t[280] ^ x[124];
  assign t[236] = t[281] ^ x[127];
  assign t[237] = t[282] ^ x[130];
  assign t[238] = t[283] ^ x[133];
  assign t[239] = t[284] ^ x[136];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[139];
  assign t[241] = t[286] ^ x[142];
  assign t[242] = t[287] ^ x[145];
  assign t[243] = t[288] ^ x[148];
  assign t[244] = t[289] ^ x[151];
  assign t[245] = (x[0] & x[1]);
  assign t[246] = (x[8] & x[9]);
  assign t[247] = (x[11] & x[12]);
  assign t[248] = (x[14] & x[15]);
  assign t[249] = (x[17] & x[18]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[20] & x[21]);
  assign t[251] = (x[23] & x[24]);
  assign t[252] = (x[26] & x[27]);
  assign t[253] = (x[29] & x[30]);
  assign t[254] = (x[32] & x[33]);
  assign t[255] = (x[37] & x[38]);
  assign t[256] = (x[40] & x[41]);
  assign t[257] = (x[43] & x[44]);
  assign t[258] = (x[46] & x[47]);
  assign t[259] = (x[49] & x[50]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[54] & x[55]);
  assign t[261] = (x[57] & x[58]);
  assign t[262] = (x[60] & x[61]);
  assign t[263] = (x[63] & x[64]);
  assign t[264] = (x[66] & x[67]);
  assign t[265] = (x[69] & x[70]);
  assign t[266] = (x[72] & x[73]);
  assign t[267] = (x[77] & x[78]);
  assign t[268] = (x[80] & x[81]);
  assign t[269] = (x[85] & x[86]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[88] & x[89]);
  assign t[271] = (x[91] & x[92]);
  assign t[272] = (x[94] & x[95]);
  assign t[273] = (x[97] & x[98]);
  assign t[274] = (x[100] & x[101]);
  assign t[275] = (x[105] & x[106]);
  assign t[276] = (x[108] & x[109]);
  assign t[277] = (x[111] & x[112]);
  assign t[278] = (x[116] & x[117]);
  assign t[279] = (x[119] & x[120]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[122] & x[123]);
  assign t[281] = (x[125] & x[126]);
  assign t[282] = (x[128] & x[129]);
  assign t[283] = (x[131] & x[132]);
  assign t[284] = (x[134] & x[135]);
  assign t[285] = (x[137] & x[138]);
  assign t[286] = (x[140] & x[141]);
  assign t[287] = (x[143] & x[144]);
  assign t[288] = (x[146] & x[147]);
  assign t[289] = (x[149] & x[150]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[205] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[36] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[206] | t[67]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] ^ t[79]);
  assign t[48] = ~(t[203]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[82]);
  assign t[51] = ~(t[80] | t[83]);
  assign t[52] = ~(t[207]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[209] | t[88]);
  assign t[57] = t[29] ? x[36] : x[35];
  assign t[58] = ~(t[89] & t[90]);
  assign t[59] = ~(t[91] | t[92]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[210] | t[93]);
  assign t[61] = ~(t[94] ^ t[95]);
  assign t[62] = ~(t[96] | t[97]);
  assign t[63] = ~(t[211] | t[98]);
  assign t[64] = ~(t[99] ^ t[100]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[214] | t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[29] ? x[53] : x[52];
  assign t[71] = t[106] | t[51];
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[215] | t[109]);
  assign t[74] = ~(t[110] | t[111]);
  assign t[75] = ~(t[112] ^ t[113]);
  assign t[76] = ~(t[114] | t[115]);
  assign t[77] = ~(t[216] | t[116]);
  assign t[78] = ~(t[117] | t[118]);
  assign t[79] = ~(t[119] ^ t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121]);
  assign t[81] = t[201] ? t[123] : t[122];
  assign t[82] = ~(t[124] | t[125]);
  assign t[83] = t[201] ? t[127] : t[126];
  assign t[84] = ~(t[217]);
  assign t[85] = ~(t[207] | t[208]);
  assign t[86] = ~(t[218]);
  assign t[87] = ~(t[219]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[124] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131]);
  assign t[91] = ~(t[220]);
  assign t[92] = ~(t[221]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = t[134] ? x[76] : x[75];
  assign t[95] = ~(t[135] & t[31]);
  assign t[96] = ~(t[222]);
  assign t[97] = ~(t[223]);
  assign t[98] = ~(t[136] | t[137]);
  assign t[99] = t[134] ? x[84] : x[83];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind154(x, y);
 input [151:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[32];
  assign t[117] = t[162] ^ x[35];
  assign t[118] = t[163] ^ x[38];
  assign t[119] = t[164] ^ x[41];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[46];
  assign t[121] = t[166] ^ x[51];
  assign t[122] = t[167] ^ x[54];
  assign t[123] = t[168] ^ x[57];
  assign t[124] = t[169] ^ x[60];
  assign t[125] = t[170] ^ x[65];
  assign t[126] = t[171] ^ x[70];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[76];
  assign t[129] = t[174] ^ x[79];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[82];
  assign t[131] = t[176] ^ x[85];
  assign t[132] = t[177] ^ x[88];
  assign t[133] = t[178] ^ x[91];
  assign t[134] = t[179] ^ x[94];
  assign t[135] = t[180] ^ x[97];
  assign t[136] = t[181] ^ x[100];
  assign t[137] = t[182] ^ x[103];
  assign t[138] = t[183] ^ x[106];
  assign t[139] = t[184] ^ x[109];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[112];
  assign t[141] = t[186] ^ x[115];
  assign t[142] = t[187] ^ x[118];
  assign t[143] = t[188] ^ x[121];
  assign t[144] = t[189] ^ x[124];
  assign t[145] = t[190] ^ x[127];
  assign t[146] = t[191] ^ x[130];
  assign t[147] = t[192] ^ x[133];
  assign t[148] = t[193] ^ x[136];
  assign t[149] = t[194] ^ x[139];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[142];
  assign t[151] = t[196] ^ x[145];
  assign t[152] = t[197] ^ x[148];
  assign t[153] = t[198] ^ x[151];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[30] & x[31]);
  assign t[162] = (x[33] & x[34]);
  assign t[163] = (x[36] & x[37]);
  assign t[164] = (x[39] & x[40]);
  assign t[165] = (x[44] & x[45]);
  assign t[166] = (x[49] & x[50]);
  assign t[167] = (x[52] & x[53]);
  assign t[168] = (x[55] & x[56]);
  assign t[169] = (x[58] & x[59]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[63] & x[64]);
  assign t[171] = (x[68] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[74] & x[75]);
  assign t[174] = (x[77] & x[78]);
  assign t[175] = (x[80] & x[81]);
  assign t[176] = (x[83] & x[84]);
  assign t[177] = (x[86] & x[87]);
  assign t[178] = (x[89] & x[90]);
  assign t[179] = (x[92] & x[93]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[95] & x[96]);
  assign t[181] = (x[98] & x[99]);
  assign t[182] = (x[101] & x[102]);
  assign t[183] = (x[104] & x[105]);
  assign t[184] = (x[107] & x[108]);
  assign t[185] = (x[110] & x[111]);
  assign t[186] = (x[113] & x[114]);
  assign t[187] = (x[116] & x[117]);
  assign t[188] = (x[119] & x[120]);
  assign t[189] = (x[122] & x[123]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[125] & x[126]);
  assign t[191] = (x[128] & x[129]);
  assign t[192] = (x[131] & x[132]);
  assign t[193] = (x[134] & x[135]);
  assign t[194] = (x[137] & x[138]);
  assign t[195] = (x[140] & x[141]);
  assign t[196] = (x[143] & x[144]);
  assign t[197] = (x[146] & x[147]);
  assign t[198] = (x[149] & x[150]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[33];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = t[60] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[43];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[73] | t[118];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[119];
  assign t[53] = t[17] ? x[43] : x[42];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = t[81] | t[120];
  assign t[57] = t[17] ? x[48] : x[47];
  assign t[58] = ~(t[121]);
  assign t[59] = ~(t[122]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] | t[58]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = t[85] | t[123];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = t[88] | t[124];
  assign t[65] = t[89] ? x[62] : x[61];
  assign t[66] = ~(t[90] & t[91]);
  assign t[67] = t[92] | t[125];
  assign t[68] = t[89] ? x[67] : x[66];
  assign t[69] = ~(t[93] & t[94]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[97] & t[98]);
  assign t[78] = t[99] | t[131];
  assign t[79] = ~(t[132]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[100] | t[79]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[101] | t[83]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[102] | t[86]);
  assign t[89] = ~(t[24]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[107] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind155(x, y);
 input [151:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[114] & t[115]);
  assign t[103] = ~(t[142] & t[141]);
  assign t[104] = ~(t[155]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[154] & t[153]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[32];
  assign t[126] = t[171] ^ x[35];
  assign t[127] = t[172] ^ x[38];
  assign t[128] = t[173] ^ x[41];
  assign t[129] = t[174] ^ x[46];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[51];
  assign t[131] = t[176] ^ x[54];
  assign t[132] = t[177] ^ x[57];
  assign t[133] = t[178] ^ x[60];
  assign t[134] = t[179] ^ x[65];
  assign t[135] = t[180] ^ x[70];
  assign t[136] = t[181] ^ x[73];
  assign t[137] = t[182] ^ x[76];
  assign t[138] = t[183] ^ x[79];
  assign t[139] = t[184] ^ x[82];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[85];
  assign t[141] = t[186] ^ x[88];
  assign t[142] = t[187] ^ x[91];
  assign t[143] = t[188] ^ x[94];
  assign t[144] = t[189] ^ x[97];
  assign t[145] = t[190] ^ x[100];
  assign t[146] = t[191] ^ x[103];
  assign t[147] = t[192] ^ x[106];
  assign t[148] = t[193] ^ x[109];
  assign t[149] = t[194] ^ x[112];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[118];
  assign t[152] = t[197] ^ x[121];
  assign t[153] = t[198] ^ x[124];
  assign t[154] = t[199] ^ x[127];
  assign t[155] = t[200] ^ x[130];
  assign t[156] = t[201] ^ x[133];
  assign t[157] = t[202] ^ x[136];
  assign t[158] = t[203] ^ x[139];
  assign t[159] = t[204] ^ x[142];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[145];
  assign t[161] = t[206] ^ x[148];
  assign t[162] = t[207] ^ x[151];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[30] & x[31]);
  assign t[171] = (x[33] & x[34]);
  assign t[172] = (x[36] & x[37]);
  assign t[173] = (x[39] & x[40]);
  assign t[174] = (x[44] & x[45]);
  assign t[175] = (x[49] & x[50]);
  assign t[176] = (x[52] & x[53]);
  assign t[177] = (x[55] & x[56]);
  assign t[178] = (x[58] & x[59]);
  assign t[179] = (x[63] & x[64]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[68] & x[69]);
  assign t[181] = (x[71] & x[72]);
  assign t[182] = (x[74] & x[75]);
  assign t[183] = (x[77] & x[78]);
  assign t[184] = (x[80] & x[81]);
  assign t[185] = (x[83] & x[84]);
  assign t[186] = (x[86] & x[87]);
  assign t[187] = (x[89] & x[90]);
  assign t[188] = (x[92] & x[93]);
  assign t[189] = (x[95] & x[96]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[98] & x[99]);
  assign t[191] = (x[101] & x[102]);
  assign t[192] = (x[104] & x[105]);
  assign t[193] = (x[107] & x[108]);
  assign t[194] = (x[110] & x[111]);
  assign t[195] = (x[113] & x[114]);
  assign t[196] = (x[116] & x[117]);
  assign t[197] = (x[119] & x[120]);
  assign t[198] = (x[122] & x[123]);
  assign t[199] = (x[125] & x[126]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[128] & x[129]);
  assign t[201] = (x[131] & x[132]);
  assign t[202] = (x[134] & x[135]);
  assign t[203] = (x[137] & x[138]);
  assign t[204] = (x[140] & x[141]);
  assign t[205] = (x[143] & x[144]);
  assign t[206] = (x[146] & x[147]);
  assign t[207] = (x[149] & x[150]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[33];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = ~(t[60] & t[124]);
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[43];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[127]);
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = ~(t[77] & t[128]);
  assign t[53] = t[17] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = ~(t[82] & t[129]);
  assign t[57] = t[121] ? x[48] : x[47];
  assign t[58] = ~(t[130]);
  assign t[59] = ~(t[131]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[132]);
  assign t[63] = ~(t[88] & t[89]);
  assign t[64] = ~(t[90] & t[133]);
  assign t[65] = t[48] ? x[62] : x[61];
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[134]);
  assign t[68] = t[48] ? x[67] : x[66];
  assign t[69] = ~(t[94] & t[95]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126] & t[125]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[96] & t[97]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[98] & t[99]);
  assign t[78] = ~(t[100] & t[101]);
  assign t[79] = ~(t[102] & t[140]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[103] & t[104]);
  assign t[83] = ~(t[131] & t[130]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[105] & t[106]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[107] & t[108]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[109] & t[110]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind156(x, y);
 input [121:0] x;
 output y;

 wire [167:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[13];
  assign t[101] = t[136] ^ x[16];
  assign t[102] = t[137] ^ x[19];
  assign t[103] = t[138] ^ x[22];
  assign t[104] = t[139] ^ x[25];
  assign t[105] = t[140] ^ x[30];
  assign t[106] = t[141] ^ x[33];
  assign t[107] = t[142] ^ x[38];
  assign t[108] = t[143] ^ x[41];
  assign t[109] = t[144] ^ x[44];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[47];
  assign t[111] = t[146] ^ x[50];
  assign t[112] = t[147] ^ x[55];
  assign t[113] = t[148] ^ x[58];
  assign t[114] = t[149] ^ x[63];
  assign t[115] = t[150] ^ x[66];
  assign t[116] = t[151] ^ x[69];
  assign t[117] = t[152] ^ x[72];
  assign t[118] = t[153] ^ x[75];
  assign t[119] = t[154] ^ x[80];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[155] ^ x[83];
  assign t[121] = t[156] ^ x[88];
  assign t[122] = t[157] ^ x[91];
  assign t[123] = t[158] ^ x[94];
  assign t[124] = t[159] ^ x[97];
  assign t[125] = t[160] ^ x[100];
  assign t[126] = t[161] ^ x[103];
  assign t[127] = t[162] ^ x[106];
  assign t[128] = t[163] ^ x[109];
  assign t[129] = t[164] ^ x[112];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[115];
  assign t[131] = t[166] ^ x[118];
  assign t[132] = t[167] ^ x[121];
  assign t[133] = (x[0] & x[1]);
  assign t[134] = (x[8] & x[9]);
  assign t[135] = (x[11] & x[12]);
  assign t[136] = (x[14] & x[15]);
  assign t[137] = (x[17] & x[18]);
  assign t[138] = (x[20] & x[21]);
  assign t[139] = (x[23] & x[24]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[28] & x[29]);
  assign t[141] = (x[31] & x[32]);
  assign t[142] = (x[36] & x[37]);
  assign t[143] = (x[39] & x[40]);
  assign t[144] = (x[42] & x[43]);
  assign t[145] = (x[45] & x[46]);
  assign t[146] = (x[48] & x[49]);
  assign t[147] = (x[53] & x[54]);
  assign t[148] = (x[56] & x[57]);
  assign t[149] = (x[61] & x[62]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[64] & x[65]);
  assign t[151] = (x[67] & x[68]);
  assign t[152] = (x[70] & x[71]);
  assign t[153] = (x[73] & x[74]);
  assign t[154] = (x[78] & x[79]);
  assign t[155] = (x[81] & x[82]);
  assign t[156] = (x[86] & x[87]);
  assign t[157] = (x[89] & x[90]);
  assign t[158] = (x[92] & x[93]);
  assign t[159] = (x[95] & x[96]);
  assign t[15] = ~(t[99] & t[100]);
  assign t[160] = (x[98] & x[99]);
  assign t[161] = (x[101] & x[102]);
  assign t[162] = (x[104] & x[105]);
  assign t[163] = (x[107] & x[108]);
  assign t[164] = (x[110] & x[111]);
  assign t[165] = (x[113] & x[114]);
  assign t[166] = (x[116] & x[117]);
  assign t[167] = (x[119] & x[120]);
  assign t[16] = ~(t[101] & t[102]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[101]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[103] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[104] & t[46]);
  assign t[31] = t[17] ? x[27] : x[26];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = t[51] ^ t[35];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[55];
  assign t[37] = ~(t[105] & t[56]);
  assign t[38] = ~(t[106] & t[57]);
  assign t[39] = t[17] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[41];
  assign t[45] = ~(t[107]);
  assign t[46] = ~(t[107] & t[67]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = t[72] ? x[52] : x[51];
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = t[17] ? x[60] : x[59];
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = t[72] ? x[77] : x[76];
  assign t[63] = ~(t[82] & t[83]);
  assign t[64] = ~(t[119] & t[84]);
  assign t[65] = ~(t[120] & t[85]);
  assign t[66] = t[72] ? x[85] : x[84];
  assign t[67] = ~(t[103]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[24]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131] & t[96]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[132]);
  assign t[94] = ~(t[132] & t[97]);
  assign t[95] = ~(t[119]);
  assign t[96] = ~(t[124]);
  assign t[97] = ~(t[128]);
  assign t[98] = t[133] ^ x[2];
  assign t[99] = t[134] ^ x[10];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[98];
endmodule

module R1ind157(x, y);
 input [151:0] x;
 output y;

 wire [294:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[29] ? x[79] : x[78];
  assign t[101] = ~(t[142] & t[143]);
  assign t[102] = ~(t[228]);
  assign t[103] = ~(t[229]);
  assign t[104] = ~(t[144] | t[145]);
  assign t[105] = t[29] ? x[87] : x[86];
  assign t[106] = ~(t[146] & t[147]);
  assign t[107] = ~(t[230]);
  assign t[108] = ~(t[217] | t[218]);
  assign t[109] = ~(t[231]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[232]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[233]);
  assign t[114] = ~(t[234]);
  assign t[115] = ~(t[152] | t[153]);
  assign t[116] = t[154] ? x[104] : x[103];
  assign t[117] = t[155] | t[83];
  assign t[118] = ~(t[235]);
  assign t[119] = ~(t[236]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[156] | t[157]);
  assign t[121] = ~(t[158] | t[159]);
  assign t[122] = ~(t[237] | t[160]);
  assign t[123] = t[154] ? x[115] : x[114];
  assign t[124] = ~(t[161] & t[162]);
  assign t[125] = ~(t[163] & t[164]);
  assign t[126] = ~(t[207] | t[165]);
  assign t[127] = t[128] & t[206];
  assign t[128] = ~(t[131]);
  assign t[129] = t[206] ? t[163] : t[166];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[206] ? t[168] : t[167];
  assign t[131] = ~(t[208]);
  assign t[132] = ~(t[238]);
  assign t[133] = ~(t[223] | t[224]);
  assign t[134] = ~(t[131] | t[169]);
  assign t[135] = ~(t[128] | t[170]);
  assign t[136] = ~(t[171] & t[172]);
  assign t[137] = ~(t[239]);
  assign t[138] = ~(t[225] | t[226]);
  assign t[139] = ~(t[240]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[241]);
  assign t[141] = ~(t[173] | t[174]);
  assign t[142] = ~(t[150] | t[175]);
  assign t[143] = ~(t[117] | t[176]);
  assign t[144] = ~(t[242]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[177] | t[84]);
  assign t[147] = ~(t[134] | t[155]);
  assign t[148] = ~(t[243]);
  assign t[149] = ~(t[231] | t[232]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[93] & t[179]);
  assign t[152] = ~(t[244]);
  assign t[153] = ~(t[233] | t[234]);
  assign t[154] = ~(t[48]);
  assign t[155] = ~(t[180] & t[82]);
  assign t[156] = ~(t[245]);
  assign t[157] = ~(t[235] | t[236]);
  assign t[158] = ~(t[246]);
  assign t[159] = ~(t[247]);
  assign t[15] = ~(t[206] & t[207]);
  assign t[160] = ~(t[181] | t[182]);
  assign t[161] = ~(t[150]);
  assign t[162] = ~(t[183] | t[83]);
  assign t[163] = ~(t[209] & t[184]);
  assign t[164] = ~(x[4] & t[126]);
  assign t[165] = ~(t[209]);
  assign t[166] = ~(x[4] & t[185]);
  assign t[167] = ~(t[87] & t[165]);
  assign t[168] = ~(t[86] & t[209]);
  assign t[169] = t[206] ? t[186] : t[167];
  assign t[16] = ~(t[208] & t[209]);
  assign t[170] = t[206] ? t[187] : t[164];
  assign t[171] = ~(t[150] | t[188]);
  assign t[172] = t[131] | t[189];
  assign t[173] = ~(t[248]);
  assign t[174] = ~(t[240] | t[241]);
  assign t[175] = ~(t[128] | t[190]);
  assign t[176] = ~(t[191] & t[172]);
  assign t[177] = ~(t[128] | t[192]);
  assign t[178] = t[206] ? t[193] : t[186];
  assign t[179] = ~(t[131] & t[194]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[195] | t[196]);
  assign t[181] = ~(t[249]);
  assign t[182] = ~(t[246] | t[247]);
  assign t[183] = ~(t[197]);
  assign t[184] = ~(x[4] | t[198]);
  assign t[185] = ~(t[207] | t[209]);
  assign t[186] = ~(t[86] & t[165]);
  assign t[187] = ~(t[184] & t[165]);
  assign t[188] = ~(t[128] | t[199]);
  assign t[189] = t[206] ? t[166] : t[187];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[206] ? t[166] : t[163];
  assign t[191] = ~(t[200] | t[201]);
  assign t[192] = t[206] ? t[186] : t[193];
  assign t[193] = ~(t[87] & t[209]);
  assign t[194] = ~(t[166] & t[163]);
  assign t[195] = ~(t[131] | t[202]);
  assign t[196] = ~(t[131] | t[203]);
  assign t[197] = ~(t[201] | t[188]);
  assign t[198] = ~(t[207]);
  assign t[199] = t[206] ? t[167] : t[168];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[81]);
  assign t[201] = ~(t[128] | t[204]);
  assign t[202] = t[206] ? t[167] : t[186];
  assign t[203] = t[206] ? t[187] : t[166];
  assign t[204] = t[206] ? t[164] : t[187];
  assign t[205] = t[250] ^ x[2];
  assign t[206] = t[251] ^ x[10];
  assign t[207] = t[252] ^ x[13];
  assign t[208] = t[253] ^ x[16];
  assign t[209] = t[254] ^ x[19];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[22];
  assign t[211] = t[256] ^ x[25];
  assign t[212] = t[257] ^ x[28];
  assign t[213] = t[258] ^ x[31];
  assign t[214] = t[259] ^ x[34];
  assign t[215] = t[260] ^ x[39];
  assign t[216] = t[261] ^ x[42];
  assign t[217] = t[262] ^ x[45];
  assign t[218] = t[263] ^ x[48];
  assign t[219] = t[264] ^ x[51];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[56];
  assign t[221] = t[266] ^ x[59];
  assign t[222] = t[267] ^ x[62];
  assign t[223] = t[268] ^ x[65];
  assign t[224] = t[269] ^ x[68];
  assign t[225] = t[270] ^ x[71];
  assign t[226] = t[271] ^ x[74];
  assign t[227] = t[272] ^ x[77];
  assign t[228] = t[273] ^ x[82];
  assign t[229] = t[274] ^ x[85];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[90];
  assign t[231] = t[276] ^ x[93];
  assign t[232] = t[277] ^ x[96];
  assign t[233] = t[278] ^ x[99];
  assign t[234] = t[279] ^ x[102];
  assign t[235] = t[280] ^ x[107];
  assign t[236] = t[281] ^ x[110];
  assign t[237] = t[282] ^ x[113];
  assign t[238] = t[283] ^ x[118];
  assign t[239] = t[284] ^ x[121];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[124];
  assign t[241] = t[286] ^ x[127];
  assign t[242] = t[287] ^ x[130];
  assign t[243] = t[288] ^ x[133];
  assign t[244] = t[289] ^ x[136];
  assign t[245] = t[290] ^ x[139];
  assign t[246] = t[291] ^ x[142];
  assign t[247] = t[292] ^ x[145];
  assign t[248] = t[293] ^ x[148];
  assign t[249] = t[294] ^ x[151];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[0] & x[1]);
  assign t[251] = (x[8] & x[9]);
  assign t[252] = (x[11] & x[12]);
  assign t[253] = (x[14] & x[15]);
  assign t[254] = (x[17] & x[18]);
  assign t[255] = (x[20] & x[21]);
  assign t[256] = (x[23] & x[24]);
  assign t[257] = (x[26] & x[27]);
  assign t[258] = (x[29] & x[30]);
  assign t[259] = (x[32] & x[33]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[37] & x[38]);
  assign t[261] = (x[40] & x[41]);
  assign t[262] = (x[43] & x[44]);
  assign t[263] = (x[46] & x[47]);
  assign t[264] = (x[49] & x[50]);
  assign t[265] = (x[54] & x[55]);
  assign t[266] = (x[57] & x[58]);
  assign t[267] = (x[60] & x[61]);
  assign t[268] = (x[63] & x[64]);
  assign t[269] = (x[66] & x[67]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[69] & x[70]);
  assign t[271] = (x[72] & x[73]);
  assign t[272] = (x[75] & x[76]);
  assign t[273] = (x[80] & x[81]);
  assign t[274] = (x[83] & x[84]);
  assign t[275] = (x[88] & x[89]);
  assign t[276] = (x[91] & x[92]);
  assign t[277] = (x[94] & x[95]);
  assign t[278] = (x[97] & x[98]);
  assign t[279] = (x[100] & x[101]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[105] & x[106]);
  assign t[281] = (x[108] & x[109]);
  assign t[282] = (x[111] & x[112]);
  assign t[283] = (x[116] & x[117]);
  assign t[284] = (x[119] & x[120]);
  assign t[285] = (x[122] & x[123]);
  assign t[286] = (x[125] & x[126]);
  assign t[287] = (x[128] & x[129]);
  assign t[288] = (x[131] & x[132]);
  assign t[289] = (x[134] & x[135]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[137] & x[138]);
  assign t[291] = (x[140] & x[141]);
  assign t[292] = (x[143] & x[144]);
  assign t[293] = (x[146] & x[147]);
  assign t[294] = (x[149] & x[150]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] & t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[210] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[62] ^ t[63]);
  assign t[38] = ~(t[64] | t[65]);
  assign t[39] = ~(t[36] ^ t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[67] | t[68]);
  assign t[41] = ~(t[211] | t[69]);
  assign t[42] = ~(t[70] | t[71]);
  assign t[43] = ~(t[72] ^ t[73]);
  assign t[44] = ~(t[74] | t[75]);
  assign t[45] = ~(t[46] ^ t[76]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[47] = ~(t[79] ^ t[80]);
  assign t[48] = ~(t[208]);
  assign t[49] = ~(t[81] & t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[83] | t[84];
  assign t[51] = t[209] & t[85];
  assign t[52] = t[86] | t[87];
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[214] | t[92]);
  assign t[58] = t[29] ? x[36] : x[35];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[215] | t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[100] ^ t[101]);
  assign t[64] = ~(t[102] | t[103]);
  assign t[65] = ~(t[216] | t[104]);
  assign t[66] = ~(t[105] ^ t[106]);
  assign t[67] = ~(t[217]);
  assign t[68] = ~(t[218]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[109] | t[110]);
  assign t[71] = ~(t[219] | t[111]);
  assign t[72] = t[29] ? x[53] : x[52];
  assign t[73] = ~(t[112] & t[82]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[220] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118] | t[119]);
  assign t[78] = ~(t[221] | t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[123] ^ t[124]);
  assign t[81] = ~(t[85] & t[125]);
  assign t[82] = ~(t[126] & t[127]);
  assign t[83] = ~(t[128] | t[129]);
  assign t[84] = ~(t[128] | t[130]);
  assign t[85] = ~(t[131] | t[206]);
  assign t[86] = ~(x[4] | t[207]);
  assign t[87] = x[4] & t[207];
  assign t[88] = ~(t[222]);
  assign t[89] = ~(t[212] | t[213]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = ~(t[134] | t[135]);
  assign t[94] = ~(t[84] | t[136]);
  assign t[95] = ~(t[225]);
  assign t[96] = ~(t[226]);
  assign t[97] = ~(t[137] | t[138]);
  assign t[98] = ~(t[139] | t[140]);
  assign t[99] = ~(t[227] | t[141]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[205];
endmodule

module R1ind158(x, y);
 input [139:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = t[142] ^ x[2];
  assign t[102] = t[143] ^ x[10];
  assign t[103] = t[144] ^ x[13];
  assign t[104] = t[145] ^ x[16];
  assign t[105] = t[146] ^ x[19];
  assign t[106] = t[147] ^ x[22];
  assign t[107] = t[148] ^ x[27];
  assign t[108] = t[149] ^ x[32];
  assign t[109] = t[150] ^ x[35];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[38];
  assign t[111] = t[152] ^ x[43];
  assign t[112] = t[153] ^ x[48];
  assign t[113] = t[154] ^ x[51];
  assign t[114] = t[155] ^ x[54];
  assign t[115] = t[156] ^ x[57];
  assign t[116] = t[157] ^ x[62];
  assign t[117] = t[158] ^ x[67];
  assign t[118] = t[159] ^ x[70];
  assign t[119] = t[160] ^ x[73];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[76];
  assign t[121] = t[162] ^ x[79];
  assign t[122] = t[163] ^ x[82];
  assign t[123] = t[164] ^ x[85];
  assign t[124] = t[165] ^ x[88];
  assign t[125] = t[166] ^ x[91];
  assign t[126] = t[167] ^ x[94];
  assign t[127] = t[168] ^ x[97];
  assign t[128] = t[169] ^ x[100];
  assign t[129] = t[170] ^ x[103];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[106];
  assign t[131] = t[172] ^ x[109];
  assign t[132] = t[173] ^ x[112];
  assign t[133] = t[174] ^ x[115];
  assign t[134] = t[175] ^ x[118];
  assign t[135] = t[176] ^ x[121];
  assign t[136] = t[177] ^ x[124];
  assign t[137] = t[178] ^ x[127];
  assign t[138] = t[179] ^ x[130];
  assign t[139] = t[180] ^ x[133];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[136];
  assign t[141] = t[182] ^ x[139];
  assign t[142] = (x[0] & x[1]);
  assign t[143] = (x[8] & x[9]);
  assign t[144] = (x[11] & x[12]);
  assign t[145] = (x[14] & x[15]);
  assign t[146] = (x[17] & x[18]);
  assign t[147] = (x[20] & x[21]);
  assign t[148] = (x[25] & x[26]);
  assign t[149] = (x[30] & x[31]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[33] & x[34]);
  assign t[151] = (x[36] & x[37]);
  assign t[152] = (x[41] & x[42]);
  assign t[153] = (x[46] & x[47]);
  assign t[154] = (x[49] & x[50]);
  assign t[155] = (x[52] & x[53]);
  assign t[156] = (x[55] & x[56]);
  assign t[157] = (x[60] & x[61]);
  assign t[158] = (x[65] & x[66]);
  assign t[159] = (x[68] & x[69]);
  assign t[15] = ~(t[102] & t[103]);
  assign t[160] = (x[71] & x[72]);
  assign t[161] = (x[74] & x[75]);
  assign t[162] = (x[77] & x[78]);
  assign t[163] = (x[80] & x[81]);
  assign t[164] = (x[83] & x[84]);
  assign t[165] = (x[86] & x[87]);
  assign t[166] = (x[89] & x[90]);
  assign t[167] = (x[92] & x[93]);
  assign t[168] = (x[95] & x[96]);
  assign t[169] = (x[98] & x[99]);
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = (x[101] & x[102]);
  assign t[171] = (x[104] & x[105]);
  assign t[172] = (x[107] & x[108]);
  assign t[173] = (x[110] & x[111]);
  assign t[174] = (x[113] & x[114]);
  assign t[175] = (x[116] & x[117]);
  assign t[176] = (x[119] & x[120]);
  assign t[177] = (x[122] & x[123]);
  assign t[178] = (x[125] & x[126]);
  assign t[179] = (x[128] & x[129]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[131] & x[132]);
  assign t[181] = (x[134] & x[135]);
  assign t[182] = (x[137] & x[138]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[104]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[106];
  assign t[31] = t[104] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[40];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[107];
  assign t[38] = t[17] ? x[29] : x[28];
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[42];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[108]);
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[66] | t[44]);
  assign t[47] = ~(t[67] & t[68]);
  assign t[48] = t[69] | t[110];
  assign t[49] = t[104] ? x[40] : x[39];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[70] & t[71]);
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = t[74] | t[111];
  assign t[53] = t[75] ? x[45] : x[44];
  assign t[54] = ~(t[112]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[76] | t[54]);
  assign t[57] = ~(t[77] & t[78]);
  assign t[58] = t[79] | t[114];
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[82] | t[115];
  assign t[61] = t[75] ? x[59] : x[58];
  assign t[62] = ~(t[83] & t[84]);
  assign t[63] = t[85] | t[116];
  assign t[64] = t[75] ? x[64] : x[63];
  assign t[65] = ~(t[86] & t[87]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[88] | t[67]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] & t[90]);
  assign t[71] = t[91] | t[120];
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[92] | t[72]);
  assign t[75] = ~(t[24]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[93] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[94] | t[80]);
  assign t[83] = ~(t[128]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[95] | t[83]);
  assign t[86] = ~(t[96] & t[97]);
  assign t[87] = t[98] | t[130];
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[99] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[100] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[101];
endmodule

module R1ind159(x, y);
 input [139:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[108] & t[109]);
  assign t[106] = ~(t[142] & t[141]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[32];
  assign t[118] = t[159] ^ x[35];
  assign t[119] = t[160] ^ x[38];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[43];
  assign t[121] = t[162] ^ x[48];
  assign t[122] = t[163] ^ x[51];
  assign t[123] = t[164] ^ x[54];
  assign t[124] = t[165] ^ x[57];
  assign t[125] = t[166] ^ x[62];
  assign t[126] = t[167] ^ x[67];
  assign t[127] = t[168] ^ x[70];
  assign t[128] = t[169] ^ x[73];
  assign t[129] = t[170] ^ x[76];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[79];
  assign t[131] = t[172] ^ x[82];
  assign t[132] = t[173] ^ x[85];
  assign t[133] = t[174] ^ x[88];
  assign t[134] = t[175] ^ x[91];
  assign t[135] = t[176] ^ x[94];
  assign t[136] = t[177] ^ x[97];
  assign t[137] = t[178] ^ x[100];
  assign t[138] = t[179] ^ x[103];
  assign t[139] = t[180] ^ x[106];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[109];
  assign t[141] = t[182] ^ x[112];
  assign t[142] = t[183] ^ x[115];
  assign t[143] = t[184] ^ x[118];
  assign t[144] = t[185] ^ x[121];
  assign t[145] = t[186] ^ x[124];
  assign t[146] = t[187] ^ x[127];
  assign t[147] = t[188] ^ x[130];
  assign t[148] = t[189] ^ x[133];
  assign t[149] = t[190] ^ x[136];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[139];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[30] & x[31]);
  assign t[159] = (x[33] & x[34]);
  assign t[15] = ~(t[111] & t[112]);
  assign t[160] = (x[36] & x[37]);
  assign t[161] = (x[41] & x[42]);
  assign t[162] = (x[46] & x[47]);
  assign t[163] = (x[49] & x[50]);
  assign t[164] = (x[52] & x[53]);
  assign t[165] = (x[55] & x[56]);
  assign t[166] = (x[60] & x[61]);
  assign t[167] = (x[65] & x[66]);
  assign t[168] = (x[68] & x[69]);
  assign t[169] = (x[71] & x[72]);
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = (x[74] & x[75]);
  assign t[171] = (x[77] & x[78]);
  assign t[172] = (x[80] & x[81]);
  assign t[173] = (x[83] & x[84]);
  assign t[174] = (x[86] & x[87]);
  assign t[175] = (x[89] & x[90]);
  assign t[176] = (x[92] & x[93]);
  assign t[177] = (x[95] & x[96]);
  assign t[178] = (x[98] & x[99]);
  assign t[179] = (x[101] & x[102]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[104] & x[105]);
  assign t[181] = (x[107] & x[108]);
  assign t[182] = (x[110] & x[111]);
  assign t[183] = (x[113] & x[114]);
  assign t[184] = (x[116] & x[117]);
  assign t[185] = (x[119] & x[120]);
  assign t[186] = (x[122] & x[123]);
  assign t[187] = (x[125] & x[126]);
  assign t[188] = (x[128] & x[129]);
  assign t[189] = (x[131] & x[132]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[134] & x[135]);
  assign t[191] = (x[137] & x[138]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[113]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[115]);
  assign t[31] = t[113] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[40];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = ~(t[56] & t[116]);
  assign t[38] = t[17] ? x[29] : x[28];
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[42];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[117]);
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[66] & t[67]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[70] & t[119]);
  assign t[49] = t[113] ? x[40] : x[39];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[120]);
  assign t[53] = t[17] ? x[45] : x[44];
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[80] & t[123]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[124]);
  assign t[61] = t[84] ? x[59] : x[58];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[87] & t[125]);
  assign t[64] = t[84] ? x[64] : x[63];
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = ~(t[118] & t[117]);
  assign t[67] = ~(t[126]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[90] & t[91]);
  assign t[71] = ~(t[92] & t[93]);
  assign t[72] = ~(t[94] & t[129]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[95] & t[96]);
  assign t[76] = ~(t[122] & t[121]);
  assign t[77] = ~(t[132]);
  assign t[78] = ~(t[133]);
  assign t[79] = ~(t[134]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[97] & t[98]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[99] & t[100]);
  assign t[84] = ~(t[24]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[101] & t[102]);
  assign t[88] = ~(t[103] & t[104]);
  assign t[89] = ~(t[105] & t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[106] & t[107]);
  assign t[95] = ~(t[131] & t[130]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind160(x, y);
 input [112:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[30];
  assign t[101] = t[133] ^ x[33];
  assign t[102] = t[134] ^ x[38];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[44];
  assign t[105] = t[137] ^ x[49];
  assign t[106] = t[138] ^ x[52];
  assign t[107] = t[139] ^ x[57];
  assign t[108] = t[140] ^ x[60];
  assign t[109] = t[141] ^ x[63];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[66];
  assign t[111] = t[143] ^ x[69];
  assign t[112] = t[144] ^ x[74];
  assign t[113] = t[145] ^ x[77];
  assign t[114] = t[146] ^ x[82];
  assign t[115] = t[147] ^ x[85];
  assign t[116] = t[148] ^ x[88];
  assign t[117] = t[149] ^ x[91];
  assign t[118] = t[150] ^ x[94];
  assign t[119] = t[151] ^ x[97];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[152] ^ x[100];
  assign t[121] = t[153] ^ x[103];
  assign t[122] = t[154] ^ x[106];
  assign t[123] = t[155] ^ x[109];
  assign t[124] = t[156] ^ x[112];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[23] & x[24]);
  assign t[132] = (x[28] & x[29]);
  assign t[133] = (x[31] & x[32]);
  assign t[134] = (x[36] & x[37]);
  assign t[135] = (x[39] & x[40]);
  assign t[136] = (x[42] & x[43]);
  assign t[137] = (x[47] & x[48]);
  assign t[138] = (x[50] & x[51]);
  assign t[139] = (x[55] & x[56]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[58] & x[59]);
  assign t[141] = (x[61] & x[62]);
  assign t[142] = (x[64] & x[65]);
  assign t[143] = (x[67] & x[68]);
  assign t[144] = (x[72] & x[73]);
  assign t[145] = (x[75] & x[76]);
  assign t[146] = (x[80] & x[81]);
  assign t[147] = (x[83] & x[84]);
  assign t[148] = (x[86] & x[87]);
  assign t[149] = (x[89] & x[90]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[92] & x[93]);
  assign t[151] = (x[95] & x[96]);
  assign t[152] = (x[98] & x[99]);
  assign t[153] = (x[101] & x[102]);
  assign t[154] = (x[104] & x[105]);
  assign t[155] = (x[107] & x[108]);
  assign t[156] = (x[110] & x[111]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[96] ? x[27] : x[26];
  assign t[32] = ~(t[46] & t[47]);
  assign t[33] = t[48] ^ t[49];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[42];
  assign t[36] = ~(t[100] & t[53]);
  assign t[37] = ~(t[101] & t[54]);
  assign t[38] = t[17] ? x[35] : x[34];
  assign t[39] = ~(t[55] & t[56]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = t[59] ^ t[60];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[40];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[64]);
  assign t[46] = ~(t[103] & t[65]);
  assign t[47] = ~(t[104] & t[66]);
  assign t[48] = t[96] ? x[46] : x[45];
  assign t[49] = ~(t[67] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[71] ? x[54] : x[53];
  assign t[53] = ~(t[107]);
  assign t[54] = ~(t[107] & t[72]);
  assign t[55] = ~(t[108] & t[73]);
  assign t[56] = ~(t[109] & t[74]);
  assign t[57] = ~(t[110] & t[75]);
  assign t[58] = ~(t[111] & t[76]);
  assign t[59] = t[77] ? x[71] : x[70];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[78] & t[79]);
  assign t[61] = ~(t[112] & t[80]);
  assign t[62] = ~(t[113] & t[81]);
  assign t[63] = t[77] ? x[79] : x[78];
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[114]);
  assign t[66] = ~(t[114] & t[82]);
  assign t[67] = ~(t[115] & t[83]);
  assign t[68] = ~(t[116] & t[84]);
  assign t[69] = ~(t[117]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[117] & t[85]);
  assign t[71] = ~(t[24]);
  assign t[72] = ~(t[100]);
  assign t[73] = ~(t[118]);
  assign t[74] = ~(t[118] & t[86]);
  assign t[75] = ~(t[119]);
  assign t[76] = ~(t[119] & t[87]);
  assign t[77] = ~(t[24]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[122]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[123]);
  assign t[84] = ~(t[123] & t[91]);
  assign t[85] = ~(t[105]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[124]);
  assign t[89] = ~(t[124] & t[92]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[120]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[25];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind161(x, y);
 input [139:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[205] | t[206]);
  assign t[101] = ~(t[217]);
  assign t[102] = ~(t[218]);
  assign t[103] = ~(t[137] | t[138]);
  assign t[104] = ~(t[85] | t[139]);
  assign t[105] = ~(t[140] & t[141]);
  assign t[106] = ~(t[219]);
  assign t[107] = ~(t[220]);
  assign t[108] = ~(t[142] | t[143]);
  assign t[109] = t[144] ? x[95] : x[94];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] | t[146];
  assign t[111] = ~(t[221]);
  assign t[112] = ~(t[222]);
  assign t[113] = ~(t[147] | t[148]);
  assign t[114] = ~(t[149] | t[150]);
  assign t[115] = ~(t[223] | t[151]);
  assign t[116] = t[144] ? x[106] : x[105];
  assign t[117] = ~(t[152] & t[153]);
  assign t[118] = ~(t[197]);
  assign t[119] = ~(t[154] & t[82]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[155] & t[198]);
  assign t[121] = ~(t[118] | t[156]);
  assign t[122] = ~(t[78] | t[157]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[161]);
  assign t[125] = ~(t[162] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[224]);
  assign t[128] = ~(t[211] | t[212]);
  assign t[129] = ~(t[162] | t[166]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[167] | t[168]);
  assign t[131] = ~(t[225]);
  assign t[132] = ~(t[213] | t[214]);
  assign t[133] = ~(t[226]);
  assign t[134] = ~(t[227]);
  assign t[135] = ~(t[169] | t[170]);
  assign t[136] = ~(t[171] | t[165]);
  assign t[137] = ~(t[228]);
  assign t[138] = ~(t[217] | t[218]);
  assign t[139] = t[146] | t[163];
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = t[198] & t[160];
  assign t[141] = t[154] | t[155];
  assign t[142] = ~(t[229]);
  assign t[143] = ~(t[219] | t[220]);
  assign t[144] = ~(t[47]);
  assign t[145] = ~(t[172] & t[31]);
  assign t[146] = ~(t[78] | t[173]);
  assign t[147] = ~(t[230]);
  assign t[148] = ~(t[221] | t[222]);
  assign t[149] = ~(t[231]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[232]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[48]);
  assign t[153] = ~(t[176] | t[146]);
  assign t[154] = ~(x[4] | t[196]);
  assign t[155] = x[4] & t[196];
  assign t[156] = t[195] ? t[119] : t[177];
  assign t[157] = t[195] ? t[179] : t[178];
  assign t[158] = ~(x[4] & t[180]);
  assign t[159] = ~(t[198] & t[181]);
  assign t[15] = ~(t[195] & t[196]);
  assign t[160] = ~(t[118] | t[195]);
  assign t[161] = ~(t[159] & t[178]);
  assign t[162] = ~(t[78] | t[182]);
  assign t[163] = ~(t[78] | t[183]);
  assign t[164] = ~(t[78] | t[184]);
  assign t[165] = ~(t[78] | t[185]);
  assign t[166] = ~(t[186] & t[105]);
  assign t[167] = ~(t[118] | t[187]);
  assign t[168] = t[163] | t[188];
  assign t[169] = ~(t[233]);
  assign t[16] = ~(t[197] & t[198]);
  assign t[170] = ~(t[226] | t[227]);
  assign t[171] = ~(t[78] | t[189]);
  assign t[172] = ~(t[190] | t[167]);
  assign t[173] = t[195] ? t[159] : t[158];
  assign t[174] = ~(t[234]);
  assign t[175] = ~(t[231] | t[232]);
  assign t[176] = ~(t[136]);
  assign t[177] = ~(t[155] & t[82]);
  assign t[178] = ~(x[4] & t[50]);
  assign t[179] = ~(t[181] & t[82]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[196] | t[198]);
  assign t[181] = ~(x[4] | t[191]);
  assign t[182] = t[195] ? t[119] : t[120];
  assign t[183] = t[195] ? t[192] : t[177];
  assign t[184] = t[195] ? t[158] : t[159];
  assign t[185] = t[195] ? t[177] : t[192];
  assign t[186] = ~(t[48] | t[164]);
  assign t[187] = t[195] ? t[179] : t[158];
  assign t[188] = ~(t[124]);
  assign t[189] = t[195] ? t[178] : t[179];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[118] | t[193]);
  assign t[191] = ~(t[196]);
  assign t[192] = ~(t[154] & t[198]);
  assign t[193] = t[195] ? t[177] : t[119];
  assign t[194] = t[235] ^ x[2];
  assign t[195] = t[236] ^ x[10];
  assign t[196] = t[237] ^ x[13];
  assign t[197] = t[238] ^ x[16];
  assign t[198] = t[239] ^ x[19];
  assign t[199] = t[240] ^ x[22];
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[25];
  assign t[201] = t[242] ^ x[28];
  assign t[202] = t[243] ^ x[31];
  assign t[203] = t[244] ^ x[36];
  assign t[204] = t[245] ^ x[39];
  assign t[205] = t[246] ^ x[42];
  assign t[206] = t[247] ^ x[45];
  assign t[207] = t[248] ^ x[48];
  assign t[208] = t[249] ^ x[53];
  assign t[209] = t[250] ^ x[56];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[59];
  assign t[211] = t[252] ^ x[62];
  assign t[212] = t[253] ^ x[65];
  assign t[213] = t[254] ^ x[70];
  assign t[214] = t[255] ^ x[73];
  assign t[215] = t[256] ^ x[76];
  assign t[216] = t[257] ^ x[81];
  assign t[217] = t[258] ^ x[84];
  assign t[218] = t[259] ^ x[87];
  assign t[219] = t[260] ^ x[90];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[93];
  assign t[221] = t[262] ^ x[98];
  assign t[222] = t[263] ^ x[101];
  assign t[223] = t[264] ^ x[104];
  assign t[224] = t[265] ^ x[109];
  assign t[225] = t[266] ^ x[112];
  assign t[226] = t[267] ^ x[115];
  assign t[227] = t[268] ^ x[118];
  assign t[228] = t[269] ^ x[121];
  assign t[229] = t[270] ^ x[124];
  assign t[22] = ~(t[21] ^ t[34]);
  assign t[230] = t[271] ^ x[127];
  assign t[231] = t[272] ^ x[130];
  assign t[232] = t[273] ^ x[133];
  assign t[233] = t[274] ^ x[136];
  assign t[234] = t[275] ^ x[139];
  assign t[235] = (x[0] & x[1]);
  assign t[236] = (x[8] & x[9]);
  assign t[237] = (x[11] & x[12]);
  assign t[238] = (x[14] & x[15]);
  assign t[239] = (x[17] & x[18]);
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = (x[20] & x[21]);
  assign t[241] = (x[23] & x[24]);
  assign t[242] = (x[26] & x[27]);
  assign t[243] = (x[29] & x[30]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[46] & x[47]);
  assign t[249] = (x[51] & x[52]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[54] & x[55]);
  assign t[251] = (x[57] & x[58]);
  assign t[252] = (x[60] & x[61]);
  assign t[253] = (x[63] & x[64]);
  assign t[254] = (x[68] & x[69]);
  assign t[255] = (x[71] & x[72]);
  assign t[256] = (x[74] & x[75]);
  assign t[257] = (x[79] & x[80]);
  assign t[258] = (x[82] & x[83]);
  assign t[259] = (x[85] & x[86]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[88] & x[89]);
  assign t[261] = (x[91] & x[92]);
  assign t[262] = (x[96] & x[97]);
  assign t[263] = (x[99] & x[100]);
  assign t[264] = (x[102] & x[103]);
  assign t[265] = (x[107] & x[108]);
  assign t[266] = (x[110] & x[111]);
  assign t[267] = (x[113] & x[114]);
  assign t[268] = (x[116] & x[117]);
  assign t[269] = (x[119] & x[120]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[122] & x[123]);
  assign t[271] = (x[125] & x[126]);
  assign t[272] = (x[128] & x[129]);
  assign t[273] = (x[131] & x[132]);
  assign t[274] = (x[134] & x[135]);
  assign t[275] = (x[137] & x[138]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] & t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[199] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[43] ^ t[59]);
  assign t[37] = ~(t[60] | t[61]);
  assign t[38] = ~(t[62] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[200] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[45] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[197]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[80] & t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[196] | t[82]);
  assign t[51] = t[78] & t[195];
  assign t[52] = ~(t[201]);
  assign t[53] = ~(t[202]);
  assign t[54] = ~(t[83] | t[84]);
  assign t[55] = t[197] ? x[33] : x[32];
  assign t[56] = t[85] | t[86];
  assign t[57] = ~(t[87] | t[88]);
  assign t[58] = ~(t[203] | t[89]);
  assign t[59] = ~(t[90] ^ t[91]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[92] | t[93]);
  assign t[61] = ~(t[204] | t[94]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[63] = ~(t[97] ^ t[98]);
  assign t[64] = ~(t[205]);
  assign t[65] = ~(t[206]);
  assign t[66] = ~(t[99] | t[100]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[207] | t[103]);
  assign t[69] = t[29] ? x[50] : x[49];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[104] & t[105]);
  assign t[71] = ~(t[106] | t[107]);
  assign t[72] = ~(t[208] | t[108]);
  assign t[73] = ~(t[109] ^ t[110]);
  assign t[74] = ~(t[111] | t[112]);
  assign t[75] = ~(t[209] | t[113]);
  assign t[76] = ~(t[114] | t[115]);
  assign t[77] = ~(t[116] ^ t[117]);
  assign t[78] = ~(t[118]);
  assign t[79] = t[195] ? t[120] : t[119];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] | t[122]);
  assign t[81] = ~(t[118] & t[123]);
  assign t[82] = ~(t[198]);
  assign t[83] = ~(t[210]);
  assign t[84] = ~(t[201] | t[202]);
  assign t[85] = ~(t[124] & t[31]);
  assign t[86] = ~(t[125] & t[126]);
  assign t[87] = ~(t[211]);
  assign t[88] = ~(t[212]);
  assign t[89] = ~(t[127] | t[128]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[197] ? x[67] : x[66];
  assign t[91] = ~(t[129] & t[130]);
  assign t[92] = ~(t[213]);
  assign t[93] = ~(t[214]);
  assign t[94] = ~(t[131] | t[132]);
  assign t[95] = ~(t[133] | t[134]);
  assign t[96] = ~(t[215] | t[135]);
  assign t[97] = t[197] ? x[78] : x[77];
  assign t[98] = ~(t[129] & t[136]);
  assign t[99] = ~(t[216]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[194];
endmodule

module R1ind162(x, y);
 input [151:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[107] | t[100]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[32];
  assign t[117] = t[162] ^ x[35];
  assign t[118] = t[163] ^ x[38];
  assign t[119] = t[164] ^ x[41];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[46];
  assign t[121] = t[166] ^ x[51];
  assign t[122] = t[167] ^ x[54];
  assign t[123] = t[168] ^ x[57];
  assign t[124] = t[169] ^ x[60];
  assign t[125] = t[170] ^ x[65];
  assign t[126] = t[171] ^ x[70];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[76];
  assign t[129] = t[174] ^ x[79];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[82];
  assign t[131] = t[176] ^ x[85];
  assign t[132] = t[177] ^ x[88];
  assign t[133] = t[178] ^ x[91];
  assign t[134] = t[179] ^ x[94];
  assign t[135] = t[180] ^ x[97];
  assign t[136] = t[181] ^ x[100];
  assign t[137] = t[182] ^ x[103];
  assign t[138] = t[183] ^ x[106];
  assign t[139] = t[184] ^ x[109];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[112];
  assign t[141] = t[186] ^ x[115];
  assign t[142] = t[187] ^ x[118];
  assign t[143] = t[188] ^ x[121];
  assign t[144] = t[189] ^ x[124];
  assign t[145] = t[190] ^ x[127];
  assign t[146] = t[191] ^ x[130];
  assign t[147] = t[192] ^ x[133];
  assign t[148] = t[193] ^ x[136];
  assign t[149] = t[194] ^ x[139];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[142];
  assign t[151] = t[196] ^ x[145];
  assign t[152] = t[197] ^ x[148];
  assign t[153] = t[198] ^ x[151];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[30] & x[31]);
  assign t[162] = (x[33] & x[34]);
  assign t[163] = (x[36] & x[37]);
  assign t[164] = (x[39] & x[40]);
  assign t[165] = (x[44] & x[45]);
  assign t[166] = (x[49] & x[50]);
  assign t[167] = (x[52] & x[53]);
  assign t[168] = (x[55] & x[56]);
  assign t[169] = (x[58] & x[59]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[63] & x[64]);
  assign t[171] = (x[68] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[74] & x[75]);
  assign t[174] = (x[77] & x[78]);
  assign t[175] = (x[80] & x[81]);
  assign t[176] = (x[83] & x[84]);
  assign t[177] = (x[86] & x[87]);
  assign t[178] = (x[89] & x[90]);
  assign t[179] = (x[92] & x[93]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[95] & x[96]);
  assign t[181] = (x[98] & x[99]);
  assign t[182] = (x[101] & x[102]);
  assign t[183] = (x[104] & x[105]);
  assign t[184] = (x[107] & x[108]);
  assign t[185] = (x[110] & x[111]);
  assign t[186] = (x[113] & x[114]);
  assign t[187] = (x[116] & x[117]);
  assign t[188] = (x[119] & x[120]);
  assign t[189] = (x[122] & x[123]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[125] & x[126]);
  assign t[191] = (x[128] & x[129]);
  assign t[192] = (x[131] & x[132]);
  assign t[193] = (x[134] & x[135]);
  assign t[194] = (x[137] & x[138]);
  assign t[195] = (x[140] & x[141]);
  assign t[196] = (x[143] & x[144]);
  assign t[197] = (x[146] & x[147]);
  assign t[198] = (x[149] & x[150]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[43];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[35];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = t[59] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[73] | t[118];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[119];
  assign t[53] = t[112] ? x[43] : x[42];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = t[79] | t[120];
  assign t[56] = t[112] ? x[48] : x[47];
  assign t[57] = ~(t[121]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[80] | t[57]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[123];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[124];
  assign t[64] = t[17] ? x[62] : x[61];
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = t[91] | t[125];
  assign t[68] = t[92] ? x[67] : x[66];
  assign t[69] = ~(t[93] & t[94]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[97] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[100] & t[101]);
  assign t[88] = t[102] | t[138];
  assign t[89] = ~(t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[140]);
  assign t[91] = ~(t[103] | t[89]);
  assign t[92] = ~(t[24]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind163(x, y);
 input [151:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[144] & t[143]);
  assign t[103] = ~(t[154]);
  assign t[104] = ~(t[146] & t[145]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[114] & t[115]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[32];
  assign t[126] = t[171] ^ x[35];
  assign t[127] = t[172] ^ x[38];
  assign t[128] = t[173] ^ x[41];
  assign t[129] = t[174] ^ x[46];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[51];
  assign t[131] = t[176] ^ x[54];
  assign t[132] = t[177] ^ x[57];
  assign t[133] = t[178] ^ x[60];
  assign t[134] = t[179] ^ x[65];
  assign t[135] = t[180] ^ x[70];
  assign t[136] = t[181] ^ x[73];
  assign t[137] = t[182] ^ x[76];
  assign t[138] = t[183] ^ x[79];
  assign t[139] = t[184] ^ x[82];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[85];
  assign t[141] = t[186] ^ x[88];
  assign t[142] = t[187] ^ x[91];
  assign t[143] = t[188] ^ x[94];
  assign t[144] = t[189] ^ x[97];
  assign t[145] = t[190] ^ x[100];
  assign t[146] = t[191] ^ x[103];
  assign t[147] = t[192] ^ x[106];
  assign t[148] = t[193] ^ x[109];
  assign t[149] = t[194] ^ x[112];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[118];
  assign t[152] = t[197] ^ x[121];
  assign t[153] = t[198] ^ x[124];
  assign t[154] = t[199] ^ x[127];
  assign t[155] = t[200] ^ x[130];
  assign t[156] = t[201] ^ x[133];
  assign t[157] = t[202] ^ x[136];
  assign t[158] = t[203] ^ x[139];
  assign t[159] = t[204] ^ x[142];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[145];
  assign t[161] = t[206] ^ x[148];
  assign t[162] = t[207] ^ x[151];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[30] & x[31]);
  assign t[171] = (x[33] & x[34]);
  assign t[172] = (x[36] & x[37]);
  assign t[173] = (x[39] & x[40]);
  assign t[174] = (x[44] & x[45]);
  assign t[175] = (x[49] & x[50]);
  assign t[176] = (x[52] & x[53]);
  assign t[177] = (x[55] & x[56]);
  assign t[178] = (x[58] & x[59]);
  assign t[179] = (x[63] & x[64]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[68] & x[69]);
  assign t[181] = (x[71] & x[72]);
  assign t[182] = (x[74] & x[75]);
  assign t[183] = (x[77] & x[78]);
  assign t[184] = (x[80] & x[81]);
  assign t[185] = (x[83] & x[84]);
  assign t[186] = (x[86] & x[87]);
  assign t[187] = (x[89] & x[90]);
  assign t[188] = (x[92] & x[93]);
  assign t[189] = (x[95] & x[96]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[98] & x[99]);
  assign t[191] = (x[101] & x[102]);
  assign t[192] = (x[104] & x[105]);
  assign t[193] = (x[107] & x[108]);
  assign t[194] = (x[110] & x[111]);
  assign t[195] = (x[113] & x[114]);
  assign t[196] = (x[116] & x[117]);
  assign t[197] = (x[119] & x[120]);
  assign t[198] = (x[122] & x[123]);
  assign t[199] = (x[125] & x[126]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[128] & x[129]);
  assign t[201] = (x[131] & x[132]);
  assign t[202] = (x[134] & x[135]);
  assign t[203] = (x[137] & x[138]);
  assign t[204] = (x[140] & x[141]);
  assign t[205] = (x[143] & x[144]);
  assign t[206] = (x[146] & x[147]);
  assign t[207] = (x[149] & x[150]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[43];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[35];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = ~(t[58] & t[124]);
  assign t[39] = t[121] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[127]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[128]);
  assign t[52] = t[121] ? x[43] : x[42];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = ~(t[79] & t[129]);
  assign t[55] = t[121] ? x[48] : x[47];
  assign t[56] = ~(t[130]);
  assign t[57] = ~(t[131]);
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[132]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[133]);
  assign t[63] = t[17] ? x[62] : x[61];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[134]);
  assign t[67] = t[93] ? x[67] : x[66];
  assign t[68] = ~(t[94] & t[95]);
  assign t[69] = ~(t[126] & t[125]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[135]);
  assign t[71] = ~(t[136]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[96] & t[97]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[98] & t[99]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[131] & t[130]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[102] & t[103]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[104] & t[105]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[108] & t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[109] & t[110]);
  assign t[93] = ~(t[24]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind164(x, y);
 input [121:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[25];
  assign t[106] = t[141] ^ x[30];
  assign t[107] = t[142] ^ x[33];
  assign t[108] = t[143] ^ x[38];
  assign t[109] = t[144] ^ x[41];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[44];
  assign t[111] = t[146] ^ x[47];
  assign t[112] = t[147] ^ x[50];
  assign t[113] = t[148] ^ x[55];
  assign t[114] = t[149] ^ x[58];
  assign t[115] = t[150] ^ x[63];
  assign t[116] = t[151] ^ x[66];
  assign t[117] = t[152] ^ x[69];
  assign t[118] = t[153] ^ x[72];
  assign t[119] = t[154] ^ x[75];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[155] ^ x[80];
  assign t[121] = t[156] ^ x[83];
  assign t[122] = t[157] ^ x[88];
  assign t[123] = t[158] ^ x[91];
  assign t[124] = t[159] ^ x[94];
  assign t[125] = t[160] ^ x[97];
  assign t[126] = t[161] ^ x[100];
  assign t[127] = t[162] ^ x[103];
  assign t[128] = t[163] ^ x[106];
  assign t[129] = t[164] ^ x[109];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[112];
  assign t[131] = t[166] ^ x[115];
  assign t[132] = t[167] ^ x[118];
  assign t[133] = t[168] ^ x[121];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[23] & x[24]);
  assign t[141] = (x[28] & x[29]);
  assign t[142] = (x[31] & x[32]);
  assign t[143] = (x[36] & x[37]);
  assign t[144] = (x[39] & x[40]);
  assign t[145] = (x[42] & x[43]);
  assign t[146] = (x[45] & x[46]);
  assign t[147] = (x[48] & x[49]);
  assign t[148] = (x[53] & x[54]);
  assign t[149] = (x[56] & x[57]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[61] & x[62]);
  assign t[151] = (x[64] & x[65]);
  assign t[152] = (x[67] & x[68]);
  assign t[153] = (x[70] & x[71]);
  assign t[154] = (x[73] & x[74]);
  assign t[155] = (x[78] & x[79]);
  assign t[156] = (x[81] & x[82]);
  assign t[157] = (x[86] & x[87]);
  assign t[158] = (x[89] & x[90]);
  assign t[159] = (x[92] & x[93]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[95] & x[96]);
  assign t[161] = (x[98] & x[99]);
  assign t[162] = (x[101] & x[102]);
  assign t[163] = (x[104] & x[105]);
  assign t[164] = (x[107] & x[108]);
  assign t[165] = (x[110] & x[111]);
  assign t[166] = (x[113] & x[114]);
  assign t[167] = (x[116] & x[117]);
  assign t[168] = (x[119] & x[120]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[27] : x[26];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[43];
  assign t[37] = ~(t[106] & t[56]);
  assign t[38] = ~(t[107] & t[57]);
  assign t[39] = t[58] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[70]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = t[102] ? x[52] : x[51];
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = t[102] ? x[60] : x[59];
  assign t[56] = ~(t[115]);
  assign t[57] = ~(t[115] & t[76]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[116] & t[77]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[78]);
  assign t[61] = ~(t[118] & t[79]);
  assign t[62] = ~(t[119] & t[80]);
  assign t[63] = t[47] ? x[77] : x[76];
  assign t[64] = ~(t[81] & t[82]);
  assign t[65] = ~(t[120] & t[83]);
  assign t[66] = ~(t[121] & t[84]);
  assign t[67] = t[17] ? x[85] : x[84];
  assign t[68] = ~(t[85] & t[86]);
  assign t[69] = ~(t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[124]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[106]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[116]);
  assign t[91] = ~(t[118]);
  assign t[92] = ~(t[132]);
  assign t[93] = ~(t[132] & t[97]);
  assign t[94] = ~(t[120]);
  assign t[95] = ~(t[133]);
  assign t[96] = ~(t[133] & t[98]);
  assign t[97] = ~(t[127]);
  assign t[98] = ~(t[130]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind165(x, y);
 input [151:0] x;
 output y;

 wire [300:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[233]);
  assign t[101] = ~(t[234]);
  assign t[102] = ~(t[148] | t[149]);
  assign t[103] = t[214] ? x[84] : x[83];
  assign t[104] = t[150] | t[151];
  assign t[105] = ~(t[235]);
  assign t[106] = ~(t[223] | t[224]);
  assign t[107] = ~(t[236]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[152] | t[153]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[139] | t[154]);
  assign t[111] = ~(t[155] | t[84]);
  assign t[112] = ~(t[238]);
  assign t[113] = ~(t[239]);
  assign t[114] = ~(t[156] | t[157]);
  assign t[115] = ~(t[158] | t[159]);
  assign t[116] = ~(t[240] | t[160]);
  assign t[117] = t[29] ? x[104] : x[103];
  assign t[118] = ~(t[161] & t[162]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[163] | t[164]);
  assign t[122] = ~(t[165] | t[166]);
  assign t[123] = ~(t[243] | t[167]);
  assign t[124] = t[29] ? x[115] : x[114];
  assign t[125] = ~(t[168] & t[169]);
  assign t[126] = ~(t[214]);
  assign t[127] = ~(t[170] & t[171]);
  assign t[128] = ~(t[172] & t[215]);
  assign t[129] = ~(t[215] & t[173]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(x[4] & t[174]);
  assign t[131] = ~(t[175] | t[141]);
  assign t[132] = ~(t[176] & t[177]);
  assign t[133] = t[212] ? t[129] : t[130];
  assign t[134] = ~(t[178]);
  assign t[135] = ~(t[81] | t[179]);
  assign t[136] = t[212] ? t[130] : t[180];
  assign t[137] = ~(t[244]);
  assign t[138] = ~(t[229] | t[230]);
  assign t[139] = ~(t[81] | t[181]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[30] & t[182]);
  assign t[141] = ~(t[126] | t[183]);
  assign t[142] = t[154] | t[134];
  assign t[143] = ~(t[245]);
  assign t[144] = ~(t[231] | t[232]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[150] | t[184]);
  assign t[147] = ~(t[139]);
  assign t[148] = ~(t[246]);
  assign t[149] = ~(t[233] | t[234]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[178] & t[132]);
  assign t[151] = ~(t[110] & t[185]);
  assign t[152] = ~(t[247]);
  assign t[153] = ~(t[236] | t[237]);
  assign t[154] = ~(t[81] | t[186]);
  assign t[155] = ~(t[126] | t[187]);
  assign t[156] = ~(t[248]);
  assign t[157] = ~(t[238] | t[239]);
  assign t[158] = ~(t[249]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[212] & t[213]);
  assign t[160] = ~(t[188] | t[189]);
  assign t[161] = ~(t[155] | t[190]);
  assign t[162] = ~(t[154] | t[191]);
  assign t[163] = ~(t[251]);
  assign t[164] = ~(t[241] | t[242]);
  assign t[165] = ~(t[252]);
  assign t[166] = ~(t[253]);
  assign t[167] = ~(t[192] | t[193]);
  assign t[168] = ~(t[194] | t[195]);
  assign t[169] = ~(t[49] | t[196]);
  assign t[16] = ~(t[214] & t[215]);
  assign t[170] = ~(x[4] | t[213]);
  assign t[171] = ~(t[215]);
  assign t[172] = x[4] & t[213];
  assign t[173] = ~(x[4] | t[197]);
  assign t[174] = ~(t[213] | t[215]);
  assign t[175] = ~(t[126] | t[198]);
  assign t[176] = ~(t[213] | t[171]);
  assign t[177] = t[81] & t[212];
  assign t[178] = ~(t[199] & t[200]);
  assign t[179] = t[212] ? t[201] : t[180];
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[173] & t[171]);
  assign t[181] = t[212] ? t[127] : t[128];
  assign t[182] = ~(t[202] & t[203]);
  assign t[183] = t[212] ? t[180] : t[130];
  assign t[184] = ~(t[204] & t[87]);
  assign t[185] = ~(t[50] | t[196]);
  assign t[186] = t[212] ? t[206] : t[205];
  assign t[187] = t[212] ? t[127] : t[205];
  assign t[188] = ~(t[254]);
  assign t[189] = ~(t[249] | t[250]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[81] | t[207]);
  assign t[191] = ~(t[169] & t[87]);
  assign t[192] = ~(t[255]);
  assign t[193] = ~(t[252] | t[253]);
  assign t[194] = ~(t[161] & t[208]);
  assign t[195] = ~(t[182] & t[87]);
  assign t[196] = ~(t[81] | t[209]);
  assign t[197] = ~(t[213]);
  assign t[198] = t[212] ? t[205] : t[127];
  assign t[199] = ~(t[126] | t[212]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[129] & t[201]);
  assign t[201] = ~(x[4] & t[176]);
  assign t[202] = t[215] & t[199];
  assign t[203] = t[170] | t[172];
  assign t[204] = ~(t[141]);
  assign t[205] = ~(t[172] & t[171]);
  assign t[206] = ~(t[170] & t[215]);
  assign t[207] = t[212] ? t[180] : t[201];
  assign t[208] = ~(t[126] & t[210]);
  assign t[209] = t[212] ? t[205] : t[206];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = ~(t[130] & t[129]);
  assign t[211] = t[256] ^ x[2];
  assign t[212] = t[257] ^ x[10];
  assign t[213] = t[258] ^ x[13];
  assign t[214] = t[259] ^ x[16];
  assign t[215] = t[260] ^ x[19];
  assign t[216] = t[261] ^ x[22];
  assign t[217] = t[262] ^ x[25];
  assign t[218] = t[263] ^ x[28];
  assign t[219] = t[264] ^ x[31];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[34];
  assign t[221] = t[266] ^ x[39];
  assign t[222] = t[267] ^ x[42];
  assign t[223] = t[268] ^ x[45];
  assign t[224] = t[269] ^ x[48];
  assign t[225] = t[270] ^ x[51];
  assign t[226] = t[271] ^ x[56];
  assign t[227] = t[272] ^ x[59];
  assign t[228] = t[273] ^ x[62];
  assign t[229] = t[274] ^ x[65];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[68];
  assign t[231] = t[276] ^ x[71];
  assign t[232] = t[277] ^ x[74];
  assign t[233] = t[278] ^ x[79];
  assign t[234] = t[279] ^ x[82];
  assign t[235] = t[280] ^ x[87];
  assign t[236] = t[281] ^ x[90];
  assign t[237] = t[282] ^ x[93];
  assign t[238] = t[283] ^ x[96];
  assign t[239] = t[284] ^ x[99];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[102];
  assign t[241] = t[286] ^ x[107];
  assign t[242] = t[287] ^ x[110];
  assign t[243] = t[288] ^ x[113];
  assign t[244] = t[289] ^ x[118];
  assign t[245] = t[290] ^ x[121];
  assign t[246] = t[291] ^ x[124];
  assign t[247] = t[292] ^ x[127];
  assign t[248] = t[293] ^ x[130];
  assign t[249] = t[294] ^ x[133];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = t[295] ^ x[136];
  assign t[251] = t[296] ^ x[139];
  assign t[252] = t[297] ^ x[142];
  assign t[253] = t[298] ^ x[145];
  assign t[254] = t[299] ^ x[148];
  assign t[255] = t[300] ^ x[151];
  assign t[256] = (x[0] & x[1]);
  assign t[257] = (x[8] & x[9]);
  assign t[258] = (x[11] & x[12]);
  assign t[259] = (x[14] & x[15]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[17] & x[18]);
  assign t[261] = (x[20] & x[21]);
  assign t[262] = (x[23] & x[24]);
  assign t[263] = (x[26] & x[27]);
  assign t[264] = (x[29] & x[30]);
  assign t[265] = (x[32] & x[33]);
  assign t[266] = (x[37] & x[38]);
  assign t[267] = (x[40] & x[41]);
  assign t[268] = (x[43] & x[44]);
  assign t[269] = (x[46] & x[47]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[49] & x[50]);
  assign t[271] = (x[54] & x[55]);
  assign t[272] = (x[57] & x[58]);
  assign t[273] = (x[60] & x[61]);
  assign t[274] = (x[63] & x[64]);
  assign t[275] = (x[66] & x[67]);
  assign t[276] = (x[69] & x[70]);
  assign t[277] = (x[72] & x[73]);
  assign t[278] = (x[77] & x[78]);
  assign t[279] = (x[80] & x[81]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[85] & x[86]);
  assign t[281] = (x[88] & x[89]);
  assign t[282] = (x[91] & x[92]);
  assign t[283] = (x[94] & x[95]);
  assign t[284] = (x[97] & x[98]);
  assign t[285] = (x[100] & x[101]);
  assign t[286] = (x[105] & x[106]);
  assign t[287] = (x[108] & x[109]);
  assign t[288] = (x[111] & x[112]);
  assign t[289] = (x[116] & x[117]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[119] & x[120]);
  assign t[291] = (x[122] & x[123]);
  assign t[292] = (x[125] & x[126]);
  assign t[293] = (x[128] & x[129]);
  assign t[294] = (x[131] & x[132]);
  assign t[295] = (x[134] & x[135]);
  assign t[296] = (x[137] & x[138]);
  assign t[297] = (x[140] & x[141]);
  assign t[298] = (x[143] & x[144]);
  assign t[299] = (x[146] & x[147]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[149] & x[150]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[216] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[44] ^ t[62]);
  assign t[38] = ~(t[63] | t[64]);
  assign t[39] = ~(t[38] ^ t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[66] | t[67]);
  assign t[41] = ~(t[217] | t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[47] = ~(t[79] ^ t[80]);
  assign t[48] = ~(t[214]);
  assign t[49] = ~(t[81] | t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81] | t[83]);
  assign t[51] = t[84] | t[85];
  assign t[52] = ~(t[86] & t[87]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[220] | t[92]);
  assign t[58] = t[214] ? x[36] : x[35];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[221] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[100] | t[101]);
  assign t[64] = ~(t[222] | t[102]);
  assign t[65] = ~(t[103] ^ t[104]);
  assign t[66] = ~(t[223]);
  assign t[67] = ~(t[224]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[225] | t[109]);
  assign t[71] = t[29] ? x[53] : x[52];
  assign t[72] = ~(t[110] & t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[226] | t[114]);
  assign t[75] = ~(t[115] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[227] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[212] ? t[128] : t[127];
  assign t[83] = t[212] ? t[130] : t[129];
  assign t[84] = ~(t[131] & t[132]);
  assign t[85] = ~(t[81] | t[133]);
  assign t[86] = ~(t[134] | t[135]);
  assign t[87] = t[126] | t[136];
  assign t[88] = ~(t[228]);
  assign t[89] = ~(t[218] | t[219]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[229]);
  assign t[91] = ~(t[230]);
  assign t[92] = ~(t[137] | t[138]);
  assign t[93] = ~(t[139] | t[140]);
  assign t[94] = ~(t[141] | t[142]);
  assign t[95] = ~(t[231]);
  assign t[96] = ~(t[232]);
  assign t[97] = ~(t[143] | t[144]);
  assign t[98] = t[145] ? x[76] : x[75];
  assign t[99] = ~(t[146] & t[147]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[211];
endmodule

module R1ind166(x, y);
 input [106:0] x;
 output y;

 wire [142:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[76];
  assign t[101] = t[133] ^ x[79];
  assign t[102] = t[134] ^ x[82];
  assign t[103] = t[135] ^ x[85];
  assign t[104] = t[136] ^ x[88];
  assign t[105] = t[137] ^ x[91];
  assign t[106] = t[138] ^ x[94];
  assign t[107] = t[139] ^ x[97];
  assign t[108] = t[140] ^ x[100];
  assign t[109] = t[141] ^ x[103];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[106];
  assign t[111] = (x[0] & x[1]);
  assign t[112] = (x[8] & x[9]);
  assign t[113] = (x[11] & x[12]);
  assign t[114] = (x[14] & x[15]);
  assign t[115] = (x[17] & x[18]);
  assign t[116] = (x[20] & x[21]);
  assign t[117] = (x[23] & x[24]);
  assign t[118] = (x[28] & x[29]);
  assign t[119] = (x[31] & x[32]);
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = (x[34] & x[35]);
  assign t[121] = (x[39] & x[40]);
  assign t[122] = (x[44] & x[45]);
  assign t[123] = (x[47] & x[48]);
  assign t[124] = (x[50] & x[51]);
  assign t[125] = (x[53] & x[54]);
  assign t[126] = (x[56] & x[57]);
  assign t[127] = (x[59] & x[60]);
  assign t[128] = (x[62] & x[63]);
  assign t[129] = (x[65] & x[66]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[68] & x[69]);
  assign t[131] = (x[71] & x[72]);
  assign t[132] = (x[74] & x[75]);
  assign t[133] = (x[77] & x[78]);
  assign t[134] = (x[80] & x[81]);
  assign t[135] = (x[83] & x[84]);
  assign t[136] = (x[86] & x[87]);
  assign t[137] = (x[89] & x[90]);
  assign t[138] = (x[92] & x[93]);
  assign t[139] = (x[95] & x[96]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[98] & x[99]);
  assign t[141] = (x[101] & x[102]);
  assign t[142] = (x[104] & x[105]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[80] & t[81]);
  assign t[16] = ~(t[82] & t[83]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[82]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = t[38] | t[84];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] | t[85];
  assign t[34] = t[17] ? x[27] : x[26];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[86]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[52] | t[36]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[88];
  assign t[41] = t[17] ? x[38] : x[37];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = t[60] | t[89];
  assign t[45] = t[61] ? x[43] : x[42];
  assign t[46] = ~(t[62] & t[63]);
  assign t[47] = ~(t[79]);
  assign t[48] = ~(t[90]);
  assign t[49] = ~(t[64] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[65] & t[66]);
  assign t[51] = t[67] | t[91];
  assign t[52] = ~(t[92]);
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[68] | t[53]);
  assign t[56] = ~(t[69] & t[70]);
  assign t[57] = t[71] | t[95];
  assign t[58] = ~(t[96]);
  assign t[59] = ~(t[97]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[72] | t[58]);
  assign t[61] = ~(t[23]);
  assign t[62] = ~(t[73] & t[74]);
  assign t[63] = t[75] | t[98];
  assign t[64] = ~(t[99]);
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[76] | t[65]);
  assign t[68] = ~(t[102]);
  assign t[69] = ~(t[103]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[77] | t[69]);
  assign t[72] = ~(t[105]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[78] | t[73]);
  assign t[76] = ~(t[108]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = t[111] ^ x[2];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[112] ^ x[10];
  assign t[81] = t[113] ^ x[13];
  assign t[82] = t[114] ^ x[16];
  assign t[83] = t[115] ^ x[19];
  assign t[84] = t[116] ^ x[22];
  assign t[85] = t[117] ^ x[25];
  assign t[86] = t[118] ^ x[30];
  assign t[87] = t[119] ^ x[33];
  assign t[88] = t[120] ^ x[36];
  assign t[89] = t[121] ^ x[41];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[46];
  assign t[91] = t[123] ^ x[49];
  assign t[92] = t[124] ^ x[52];
  assign t[93] = t[125] ^ x[55];
  assign t[94] = t[126] ^ x[58];
  assign t[95] = t[127] ^ x[61];
  assign t[96] = t[128] ^ x[64];
  assign t[97] = t[129] ^ x[67];
  assign t[98] = t[130] ^ x[70];
  assign t[99] = t[131] ^ x[73];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[79];
endmodule

module R1ind167(x, y);
 input [106:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[55];
  assign t[101] = t[133] ^ x[58];
  assign t[102] = t[134] ^ x[61];
  assign t[103] = t[135] ^ x[64];
  assign t[104] = t[136] ^ x[67];
  assign t[105] = t[137] ^ x[70];
  assign t[106] = t[138] ^ x[73];
  assign t[107] = t[139] ^ x[76];
  assign t[108] = t[140] ^ x[79];
  assign t[109] = t[141] ^ x[82];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[85];
  assign t[111] = t[143] ^ x[88];
  assign t[112] = t[144] ^ x[91];
  assign t[113] = t[145] ^ x[94];
  assign t[114] = t[146] ^ x[97];
  assign t[115] = t[147] ^ x[100];
  assign t[116] = t[148] ^ x[103];
  assign t[117] = t[149] ^ x[106];
  assign t[118] = (x[0] & x[1]);
  assign t[119] = (x[8] & x[9]);
  assign t[11] = t[87] ? x[6] : x[7];
  assign t[120] = (x[11] & x[12]);
  assign t[121] = (x[14] & x[15]);
  assign t[122] = (x[17] & x[18]);
  assign t[123] = (x[20] & x[21]);
  assign t[124] = (x[23] & x[24]);
  assign t[125] = (x[28] & x[29]);
  assign t[126] = (x[31] & x[32]);
  assign t[127] = (x[34] & x[35]);
  assign t[128] = (x[39] & x[40]);
  assign t[129] = (x[44] & x[45]);
  assign t[12] = ~(t[17] ^ t[14]);
  assign t[130] = (x[47] & x[48]);
  assign t[131] = (x[50] & x[51]);
  assign t[132] = (x[53] & x[54]);
  assign t[133] = (x[56] & x[57]);
  assign t[134] = (x[59] & x[60]);
  assign t[135] = (x[62] & x[63]);
  assign t[136] = (x[65] & x[66]);
  assign t[137] = (x[68] & x[69]);
  assign t[138] = (x[71] & x[72]);
  assign t[139] = (x[74] & x[75]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[77] & x[78]);
  assign t[141] = (x[80] & x[81]);
  assign t[142] = (x[83] & x[84]);
  assign t[143] = (x[86] & x[87]);
  assign t[144] = (x[89] & x[90]);
  assign t[145] = (x[92] & x[93]);
  assign t[146] = (x[95] & x[96]);
  assign t[147] = (x[98] & x[99]);
  assign t[148] = (x[101] & x[102]);
  assign t[149] = (x[104] & x[105]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[15] = ~(t[88] & t[89]);
  assign t[16] = ~(t[87] & t[90]);
  assign t[17] = x[4] ? t[23] : t[22];
  assign t[18] = ~(t[24] & t[25]);
  assign t[19] = t[11] ^ t[22];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[27] : t[26];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] ^ t[33];
  assign t[24] = ~(t[34] & t[35]);
  assign t[25] = ~(t[36] & t[91]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[27] = t[39] ^ t[40];
  assign t[28] = ~(t[41] & t[42]);
  assign t[29] = t[43] ^ t[44];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[31] = ~(t[47] & t[92]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[93]);
  assign t[35] = ~(t[94]);
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[53] & t[54]);
  assign t[38] = ~(t[55] & t[95]);
  assign t[39] = t[48] ? x[38] : x[37];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[57]);
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = ~(t[60] & t[96]);
  assign t[43] = t[61] ? x[43] : x[42];
  assign t[44] = ~(t[62] & t[63]);
  assign t[45] = ~(t[97]);
  assign t[46] = ~(t[98]);
  assign t[47] = ~(t[64] & t[65]);
  assign t[48] = ~(t[66]);
  assign t[49] = ~(t[67] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[69] & t[99]);
  assign t[51] = ~(t[94] & t[93]);
  assign t[52] = ~(t[100]);
  assign t[53] = ~(t[101]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(t[70] & t[71]);
  assign t[56] = ~(t[72] & t[73]);
  assign t[57] = ~(t[74] & t[103]);
  assign t[58] = ~(t[104]);
  assign t[59] = ~(t[105]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[75] & t[76]);
  assign t[61] = ~(t[66]);
  assign t[62] = ~(t[77] & t[78]);
  assign t[63] = ~(t[79] & t[106]);
  assign t[64] = ~(t[98] & t[97]);
  assign t[65] = ~(t[86]);
  assign t[66] = ~(t[87]);
  assign t[67] = ~(t[107]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[80] & t[81]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[102] & t[101]);
  assign t[71] = ~(t[109]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[82] & t[83]);
  assign t[75] = ~(t[105] & t[104]);
  assign t[76] = ~(t[112]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[84] & t[85]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[108] & t[107]);
  assign t[81] = ~(t[115]);
  assign t[82] = ~(t[111] & t[110]);
  assign t[83] = ~(t[116]);
  assign t[84] = ~(t[114] & t[113]);
  assign t[85] = ~(t[117]);
  assign t[86] = t[118] ^ x[2];
  assign t[87] = t[119] ^ x[10];
  assign t[88] = t[120] ^ x[13];
  assign t[89] = t[121] ^ x[16];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[19];
  assign t[91] = t[123] ^ x[22];
  assign t[92] = t[124] ^ x[25];
  assign t[93] = t[125] ^ x[30];
  assign t[94] = t[126] ^ x[33];
  assign t[95] = t[127] ^ x[36];
  assign t[96] = t[128] ^ x[41];
  assign t[97] = t[129] ^ x[46];
  assign t[98] = t[130] ^ x[49];
  assign t[99] = t[131] ^ x[52];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[86];
endmodule

module R1ind168(x, y);
 input [88:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[8] & x[9]);
  assign t[101] = (x[11] & x[12]);
  assign t[102] = (x[14] & x[15]);
  assign t[103] = (x[17] & x[18]);
  assign t[104] = (x[20] & x[21]);
  assign t[105] = (x[23] & x[24]);
  assign t[106] = (x[26] & x[27]);
  assign t[107] = (x[29] & x[30]);
  assign t[108] = (x[34] & x[35]);
  assign t[109] = (x[37] & x[38]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[40] & x[41]);
  assign t[111] = (x[45] & x[46]);
  assign t[112] = (x[48] & x[49]);
  assign t[113] = (x[53] & x[54]);
  assign t[114] = (x[56] & x[57]);
  assign t[115] = (x[59] & x[60]);
  assign t[116] = (x[62] & x[63]);
  assign t[117] = (x[65] & x[66]);
  assign t[118] = (x[68] & x[69]);
  assign t[119] = (x[71] & x[72]);
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = (x[74] & x[75]);
  assign t[121] = (x[77] & x[78]);
  assign t[122] = (x[80] & x[81]);
  assign t[123] = (x[83] & x[84]);
  assign t[124] = (x[86] & x[87]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[74] & t[75]);
  assign t[16] = ~(t[76] & t[77]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[76]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[78] & t[36]);
  assign t[27] = ~(t[79] & t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[80] & t[46]);
  assign t[33] = ~(t[81] & t[47]);
  assign t[34] = t[48] ? x[33] : x[32];
  assign t[35] = ~(t[49] & t[50]);
  assign t[36] = ~(t[82]);
  assign t[37] = ~(t[82] & t[51]);
  assign t[38] = ~(t[83] & t[52]);
  assign t[39] = ~(t[84] & t[53]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[54] ? x[44] : x[43];
  assign t[41] = ~(t[55] & t[56]);
  assign t[42] = ~(t[85] & t[57]);
  assign t[43] = ~(t[86] & t[58]);
  assign t[44] = t[48] ? x[52] : x[51];
  assign t[45] = ~(t[59] & t[60]);
  assign t[46] = ~(t[87]);
  assign t[47] = ~(t[87] & t[61]);
  assign t[48] = ~(t[23]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[78]);
  assign t[52] = ~(t[90]);
  assign t[53] = ~(t[90] & t[64]);
  assign t[54] = ~(t[23]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[80]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[96] & t[70]);
  assign t[64] = ~(t[83]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[97] & t[71]);
  assign t[67] = ~(t[85]);
  assign t[68] = ~(t[98]);
  assign t[69] = ~(t[98] & t[72]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[88]);
  assign t[71] = ~(t[91]);
  assign t[72] = ~(t[94]);
  assign t[73] = t[99] ^ x[2];
  assign t[74] = t[100] ^ x[10];
  assign t[75] = t[101] ^ x[13];
  assign t[76] = t[102] ^ x[16];
  assign t[77] = t[103] ^ x[19];
  assign t[78] = t[104] ^ x[22];
  assign t[79] = t[105] ^ x[25];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] ^ x[28];
  assign t[81] = t[107] ^ x[31];
  assign t[82] = t[108] ^ x[36];
  assign t[83] = t[109] ^ x[39];
  assign t[84] = t[110] ^ x[42];
  assign t[85] = t[111] ^ x[47];
  assign t[86] = t[112] ^ x[50];
  assign t[87] = t[113] ^ x[55];
  assign t[88] = t[114] ^ x[58];
  assign t[89] = t[115] ^ x[61];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[116] ^ x[64];
  assign t[91] = t[117] ^ x[67];
  assign t[92] = t[118] ^ x[70];
  assign t[93] = t[119] ^ x[73];
  assign t[94] = t[120] ^ x[76];
  assign t[95] = t[121] ^ x[79];
  assign t[96] = t[122] ^ x[82];
  assign t[97] = t[123] ^ x[85];
  assign t[98] = t[124] ^ x[88];
  assign t[99] = (x[0] & x[1]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[73];
endmodule

module R1ind169(x, y);
 input [106:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[184]);
  assign t[101] = ~(t[176] | t[177]);
  assign t[102] = ~(t[185]);
  assign t[103] = ~(t[186]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[42] | t[127]);
  assign t[106] = ~(t[41] | t[128]);
  assign t[107] = ~(t[187]);
  assign t[108] = ~(t[179] | t[180]);
  assign t[109] = ~(t[188]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[189]);
  assign t[111] = ~(t[129] | t[130]);
  assign t[112] = ~(t[131] | t[132]);
  assign t[113] = ~(t[116] | t[133]);
  assign t[114] = ~(t[190]);
  assign t[115] = ~(t[182] | t[183]);
  assign t[116] = ~(t[62] | t[134]);
  assign t[117] = ~(t[62] | t[135]);
  assign t[118] = t[43] | t[136];
  assign t[119] = ~(t[137] & t[138]);
  assign t[11] = ~(t[17] ^ t[14]);
  assign t[120] = x[4] & t[163];
  assign t[121] = ~(x[4] | t[163]);
  assign t[122] = ~(t[165]);
  assign t[123] = t[162] ? t[94] : t[93];
  assign t[124] = t[162] ? t[140] : t[139];
  assign t[125] = ~(t[191]);
  assign t[126] = ~(t[185] | t[186]);
  assign t[127] = ~(t[62] | t[141]);
  assign t[128] = ~(t[113] & t[138]);
  assign t[129] = ~(t[192]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[188] | t[189]);
  assign t[131] = ~(t[105] & t[142]);
  assign t[132] = ~(t[143] & t[138]);
  assign t[133] = ~(t[62] | t[144]);
  assign t[134] = t[162] ? t[92] : t[93];
  assign t[135] = t[162] ? t[139] : t[145];
  assign t[136] = ~(t[62] | t[146]);
  assign t[137] = ~(t[147] | t[148]);
  assign t[138] = t[65] | t[149];
  assign t[139] = ~(x[4] & t[150]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = ~(t[151] & t[122]);
  assign t[141] = t[162] ? t[140] : t[152];
  assign t[142] = ~(t[65] & t[153]);
  assign t[143] = ~(t[154] & t[155]);
  assign t[144] = t[162] ? t[94] : t[95];
  assign t[145] = ~(t[165] & t[151]);
  assign t[146] = t[162] ? t[145] : t[139];
  assign t[147] = ~(t[156]);
  assign t[148] = ~(t[62] | t[157]);
  assign t[149] = t[162] ? t[139] : t[140];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = ~(t[163] | t[165]);
  assign t[151] = ~(x[4] | t[158]);
  assign t[152] = ~(x[4] & t[98]);
  assign t[153] = ~(t[139] & t[145]);
  assign t[154] = t[165] & t[159];
  assign t[155] = t[121] | t[120];
  assign t[156] = ~(t[159] & t[160]);
  assign t[157] = t[162] ? t[152] : t[140];
  assign t[158] = ~(t[163]);
  assign t[159] = ~(t[65] | t[162]);
  assign t[15] = ~(t[162] & t[163]);
  assign t[160] = ~(t[145] & t[152]);
  assign t[161] = t[193] ^ x[2];
  assign t[162] = t[194] ^ x[10];
  assign t[163] = t[195] ^ x[13];
  assign t[164] = t[196] ^ x[16];
  assign t[165] = t[197] ^ x[19];
  assign t[166] = t[198] ^ x[22];
  assign t[167] = t[199] ^ x[25];
  assign t[168] = t[200] ^ x[28];
  assign t[169] = t[201] ^ x[31];
  assign t[16] = ~(t[164] & t[165]);
  assign t[170] = t[202] ^ x[34];
  assign t[171] = t[203] ^ x[37];
  assign t[172] = t[204] ^ x[40];
  assign t[173] = t[205] ^ x[43];
  assign t[174] = t[206] ^ x[46];
  assign t[175] = t[207] ^ x[51];
  assign t[176] = t[208] ^ x[54];
  assign t[177] = t[209] ^ x[57];
  assign t[178] = t[210] ^ x[60];
  assign t[179] = t[211] ^ x[65];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[212] ^ x[68];
  assign t[181] = t[213] ^ x[71];
  assign t[182] = t[214] ^ x[76];
  assign t[183] = t[215] ^ x[79];
  assign t[184] = t[216] ^ x[82];
  assign t[185] = t[217] ^ x[85];
  assign t[186] = t[218] ^ x[88];
  assign t[187] = t[219] ^ x[91];
  assign t[188] = t[220] ^ x[94];
  assign t[189] = t[221] ^ x[97];
  assign t[18] = t[26] ? x[6] : x[7];
  assign t[190] = t[222] ^ x[100];
  assign t[191] = t[223] ^ x[103];
  assign t[192] = t[224] ^ x[106];
  assign t[193] = (x[0] & x[1]);
  assign t[194] = (x[8] & x[9]);
  assign t[195] = (x[11] & x[12]);
  assign t[196] = (x[14] & x[15]);
  assign t[197] = (x[17] & x[18]);
  assign t[198] = (x[20] & x[21]);
  assign t[199] = (x[23] & x[24]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[26] & x[27]);
  assign t[201] = (x[29] & x[30]);
  assign t[202] = (x[32] & x[33]);
  assign t[203] = (x[35] & x[36]);
  assign t[204] = (x[38] & x[39]);
  assign t[205] = (x[41] & x[42]);
  assign t[206] = (x[44] & x[45]);
  assign t[207] = (x[49] & x[50]);
  assign t[208] = (x[52] & x[53]);
  assign t[209] = (x[55] & x[56]);
  assign t[20] = ~(t[29] | t[30]);
  assign t[210] = (x[58] & x[59]);
  assign t[211] = (x[63] & x[64]);
  assign t[212] = (x[66] & x[67]);
  assign t[213] = (x[69] & x[70]);
  assign t[214] = (x[74] & x[75]);
  assign t[215] = (x[77] & x[78]);
  assign t[216] = (x[80] & x[81]);
  assign t[217] = (x[83] & x[84]);
  assign t[218] = (x[86] & x[87]);
  assign t[219] = (x[89] & x[90]);
  assign t[21] = ~(t[24] ^ t[12]);
  assign t[220] = (x[92] & x[93]);
  assign t[221] = (x[95] & x[96]);
  assign t[222] = (x[98] & x[99]);
  assign t[223] = (x[101] & x[102]);
  assign t[224] = (x[104] & x[105]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[40] | t[41]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[29] = ~(t[44] | t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[166] | t[46]);
  assign t[31] = ~(t[47] | t[48]);
  assign t[32] = ~(t[49] ^ t[50]);
  assign t[33] = ~(t[51] | t[52]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[167] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] ^ t[61]);
  assign t[39] = ~(t[164]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] | t[63]);
  assign t[41] = ~(t[62] | t[64]);
  assign t[42] = ~(t[65] | t[66]);
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = ~(t[168]);
  assign t[45] = ~(t[169]);
  assign t[46] = ~(t[69] | t[70]);
  assign t[47] = ~(t[71] | t[72]);
  assign t[48] = ~(t[170] | t[73]);
  assign t[49] = ~(t[74] | t[75]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[76] ^ t[77]);
  assign t[51] = ~(t[78] | t[79]);
  assign t[52] = ~(t[171] | t[80]);
  assign t[53] = ~(t[81] | t[82]);
  assign t[54] = ~(t[83] ^ t[84]);
  assign t[55] = ~(t[172]);
  assign t[56] = ~(t[173]);
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[87] | t[88]);
  assign t[59] = ~(t[174] | t[89]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[26] ? x[48] : x[47];
  assign t[61] = ~(t[90] & t[91]);
  assign t[62] = ~(t[65]);
  assign t[63] = t[162] ? t[93] : t[92];
  assign t[64] = t[162] ? t[95] : t[94];
  assign t[65] = ~(t[164]);
  assign t[66] = t[162] ? t[93] : t[94];
  assign t[67] = ~(t[96] | t[97]);
  assign t[68] = ~(t[98] & t[99]);
  assign t[69] = ~(t[175]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[168] | t[169]);
  assign t[71] = ~(t[176]);
  assign t[72] = ~(t[177]);
  assign t[73] = ~(t[100] | t[101]);
  assign t[74] = ~(t[102] | t[103]);
  assign t[75] = ~(t[178] | t[104]);
  assign t[76] = t[26] ? x[62] : x[61];
  assign t[77] = ~(t[105] & t[106]);
  assign t[78] = ~(t[179]);
  assign t[79] = ~(t[180]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[107] | t[108]);
  assign t[81] = ~(t[109] | t[110]);
  assign t[82] = ~(t[181] | t[111]);
  assign t[83] = t[26] ? x[73] : x[72];
  assign t[84] = ~(t[112] & t[113]);
  assign t[85] = ~(t[161]);
  assign t[86] = ~(t[172] | t[173]);
  assign t[87] = ~(t[182]);
  assign t[88] = ~(t[183]);
  assign t[89] = ~(t[114] | t[115]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[116] | t[117]);
  assign t[91] = ~(t[118] | t[119]);
  assign t[92] = ~(t[120] & t[165]);
  assign t[93] = ~(t[121] & t[122]);
  assign t[94] = ~(t[120] & t[122]);
  assign t[95] = ~(t[121] & t[165]);
  assign t[96] = ~(t[65] | t[123]);
  assign t[97] = ~(t[65] | t[124]);
  assign t[98] = ~(t[163] | t[122]);
  assign t[99] = t[62] & t[162];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[161];
endmodule

module R1ind170(x, y);
 input [139:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = t[143] ^ x[2];
  assign t[103] = t[144] ^ x[10];
  assign t[104] = t[145] ^ x[13];
  assign t[105] = t[146] ^ x[16];
  assign t[106] = t[147] ^ x[19];
  assign t[107] = t[148] ^ x[22];
  assign t[108] = t[149] ^ x[27];
  assign t[109] = t[150] ^ x[32];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[35];
  assign t[111] = t[152] ^ x[38];
  assign t[112] = t[153] ^ x[43];
  assign t[113] = t[154] ^ x[48];
  assign t[114] = t[155] ^ x[51];
  assign t[115] = t[156] ^ x[54];
  assign t[116] = t[157] ^ x[57];
  assign t[117] = t[158] ^ x[62];
  assign t[118] = t[159] ^ x[67];
  assign t[119] = t[160] ^ x[70];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[73];
  assign t[121] = t[162] ^ x[76];
  assign t[122] = t[163] ^ x[79];
  assign t[123] = t[164] ^ x[82];
  assign t[124] = t[165] ^ x[85];
  assign t[125] = t[166] ^ x[88];
  assign t[126] = t[167] ^ x[91];
  assign t[127] = t[168] ^ x[94];
  assign t[128] = t[169] ^ x[97];
  assign t[129] = t[170] ^ x[100];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[103];
  assign t[131] = t[172] ^ x[106];
  assign t[132] = t[173] ^ x[109];
  assign t[133] = t[174] ^ x[112];
  assign t[134] = t[175] ^ x[115];
  assign t[135] = t[176] ^ x[118];
  assign t[136] = t[177] ^ x[121];
  assign t[137] = t[178] ^ x[124];
  assign t[138] = t[179] ^ x[127];
  assign t[139] = t[180] ^ x[130];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[133];
  assign t[141] = t[182] ^ x[136];
  assign t[142] = t[183] ^ x[139];
  assign t[143] = (x[0] & x[1]);
  assign t[144] = (x[8] & x[9]);
  assign t[145] = (x[11] & x[12]);
  assign t[146] = (x[14] & x[15]);
  assign t[147] = (x[17] & x[18]);
  assign t[148] = (x[20] & x[21]);
  assign t[149] = (x[25] & x[26]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[30] & x[31]);
  assign t[151] = (x[33] & x[34]);
  assign t[152] = (x[36] & x[37]);
  assign t[153] = (x[41] & x[42]);
  assign t[154] = (x[46] & x[47]);
  assign t[155] = (x[49] & x[50]);
  assign t[156] = (x[52] & x[53]);
  assign t[157] = (x[55] & x[56]);
  assign t[158] = (x[60] & x[61]);
  assign t[159] = (x[65] & x[66]);
  assign t[15] = ~(t[103] & t[104]);
  assign t[160] = (x[68] & x[69]);
  assign t[161] = (x[71] & x[72]);
  assign t[162] = (x[74] & x[75]);
  assign t[163] = (x[77] & x[78]);
  assign t[164] = (x[80] & x[81]);
  assign t[165] = (x[83] & x[84]);
  assign t[166] = (x[86] & x[87]);
  assign t[167] = (x[89] & x[90]);
  assign t[168] = (x[92] & x[93]);
  assign t[169] = (x[95] & x[96]);
  assign t[16] = ~(t[105] & t[106]);
  assign t[170] = (x[98] & x[99]);
  assign t[171] = (x[101] & x[102]);
  assign t[172] = (x[104] & x[105]);
  assign t[173] = (x[107] & x[108]);
  assign t[174] = (x[110] & x[111]);
  assign t[175] = (x[113] & x[114]);
  assign t[176] = (x[116] & x[117]);
  assign t[177] = (x[119] & x[120]);
  assign t[178] = (x[122] & x[123]);
  assign t[179] = (x[125] & x[126]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[128] & x[129]);
  assign t[181] = (x[131] & x[132]);
  assign t[182] = (x[134] & x[135]);
  assign t[183] = (x[137] & x[138]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[105]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[107];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[42];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[108];
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[63];
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[40];
  assign t[44] = ~(t[109]);
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[70] | t[111];
  assign t[49] = t[71] ? x[40] : x[39];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[112];
  assign t[52] = t[17] ? x[45] : x[44];
  assign t[53] = ~(t[75] & t[76]);
  assign t[54] = ~(t[113]);
  assign t[55] = ~(t[114]);
  assign t[56] = ~(t[77] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = t[80] | t[115];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[116];
  assign t[62] = t[57] ? x[59] : x[58];
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = t[88] | t[117];
  assign t[66] = t[57] ? x[64] : x[63];
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[24]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[90] | t[72]);
  assign t[75] = ~(t[91] & t[92]);
  assign t[76] = t[93] | t[123];
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[96] & t[97]);
  assign t[85] = t[98] | t[129];
  assign t[86] = ~(t[130]);
  assign t[87] = ~(t[131]);
  assign t[88] = ~(t[99] | t[86]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[100] | t[91]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[101] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[102];
endmodule

module R1ind171(x, y);
 input [139:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[109] & t[110]);
  assign t[105] = ~(t[140] & t[139]);
  assign t[106] = ~(t[149]);
  assign t[107] = ~(t[144] & t[143]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[148] & t[147]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[151]);
  assign t[111] = t[152] ^ x[2];
  assign t[112] = t[153] ^ x[10];
  assign t[113] = t[154] ^ x[13];
  assign t[114] = t[155] ^ x[16];
  assign t[115] = t[156] ^ x[19];
  assign t[116] = t[157] ^ x[22];
  assign t[117] = t[158] ^ x[27];
  assign t[118] = t[159] ^ x[32];
  assign t[119] = t[160] ^ x[35];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[38];
  assign t[121] = t[162] ^ x[43];
  assign t[122] = t[163] ^ x[48];
  assign t[123] = t[164] ^ x[51];
  assign t[124] = t[165] ^ x[54];
  assign t[125] = t[166] ^ x[57];
  assign t[126] = t[167] ^ x[62];
  assign t[127] = t[168] ^ x[67];
  assign t[128] = t[169] ^ x[70];
  assign t[129] = t[170] ^ x[73];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[76];
  assign t[131] = t[172] ^ x[79];
  assign t[132] = t[173] ^ x[82];
  assign t[133] = t[174] ^ x[85];
  assign t[134] = t[175] ^ x[88];
  assign t[135] = t[176] ^ x[91];
  assign t[136] = t[177] ^ x[94];
  assign t[137] = t[178] ^ x[97];
  assign t[138] = t[179] ^ x[100];
  assign t[139] = t[180] ^ x[103];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[106];
  assign t[141] = t[182] ^ x[109];
  assign t[142] = t[183] ^ x[112];
  assign t[143] = t[184] ^ x[115];
  assign t[144] = t[185] ^ x[118];
  assign t[145] = t[186] ^ x[121];
  assign t[146] = t[187] ^ x[124];
  assign t[147] = t[188] ^ x[127];
  assign t[148] = t[189] ^ x[130];
  assign t[149] = t[190] ^ x[133];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[136];
  assign t[151] = t[192] ^ x[139];
  assign t[152] = (x[0] & x[1]);
  assign t[153] = (x[8] & x[9]);
  assign t[154] = (x[11] & x[12]);
  assign t[155] = (x[14] & x[15]);
  assign t[156] = (x[17] & x[18]);
  assign t[157] = (x[20] & x[21]);
  assign t[158] = (x[25] & x[26]);
  assign t[159] = (x[30] & x[31]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[33] & x[34]);
  assign t[161] = (x[36] & x[37]);
  assign t[162] = (x[41] & x[42]);
  assign t[163] = (x[46] & x[47]);
  assign t[164] = (x[49] & x[50]);
  assign t[165] = (x[52] & x[53]);
  assign t[166] = (x[55] & x[56]);
  assign t[167] = (x[60] & x[61]);
  assign t[168] = (x[65] & x[66]);
  assign t[169] = (x[68] & x[69]);
  assign t[16] = ~(t[114] & t[115]);
  assign t[170] = (x[71] & x[72]);
  assign t[171] = (x[74] & x[75]);
  assign t[172] = (x[77] & x[78]);
  assign t[173] = (x[80] & x[81]);
  assign t[174] = (x[83] & x[84]);
  assign t[175] = (x[86] & x[87]);
  assign t[176] = (x[89] & x[90]);
  assign t[177] = (x[92] & x[93]);
  assign t[178] = (x[95] & x[96]);
  assign t[179] = (x[98] & x[99]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[101] & x[102]);
  assign t[181] = (x[104] & x[105]);
  assign t[182] = (x[107] & x[108]);
  assign t[183] = (x[110] & x[111]);
  assign t[184] = (x[113] & x[114]);
  assign t[185] = (x[116] & x[117]);
  assign t[186] = (x[119] & x[120]);
  assign t[187] = (x[122] & x[123]);
  assign t[188] = (x[125] & x[126]);
  assign t[189] = (x[128] & x[129]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[131] & x[132]);
  assign t[191] = (x[134] & x[135]);
  assign t[192] = (x[137] & x[138]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[114]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[116]);
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = t[50] ^ t[42];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = ~(t[57] & t[117]);
  assign t[38] = t[58] ? x[29] : x[28];
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[40];
  assign t[44] = ~(t[118]);
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[120]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[17] ? x[40] : x[39];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[121]);
  assign t[53] = t[47] ? x[45] : x[44];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] & t[124]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = ~(t[85] & t[125]);
  assign t[63] = t[58] ? x[59] : x[58];
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = ~(t[90] & t[126]);
  assign t[67] = t[114] ? x[64] : x[63];
  assign t[68] = ~(t[119] & t[118]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[93] & t[94]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[97] & t[132]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[103]);
  assign t[87] = ~(t[104] & t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[107] & t[108]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[111];
endmodule

module R1ind172(x, y);
 input [112:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[30];
  assign t[101] = t[133] ^ x[33];
  assign t[102] = t[134] ^ x[38];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[44];
  assign t[105] = t[137] ^ x[49];
  assign t[106] = t[138] ^ x[52];
  assign t[107] = t[139] ^ x[57];
  assign t[108] = t[140] ^ x[60];
  assign t[109] = t[141] ^ x[63];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[66];
  assign t[111] = t[143] ^ x[69];
  assign t[112] = t[144] ^ x[74];
  assign t[113] = t[145] ^ x[77];
  assign t[114] = t[146] ^ x[82];
  assign t[115] = t[147] ^ x[85];
  assign t[116] = t[148] ^ x[88];
  assign t[117] = t[149] ^ x[91];
  assign t[118] = t[150] ^ x[94];
  assign t[119] = t[151] ^ x[97];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[152] ^ x[100];
  assign t[121] = t[153] ^ x[103];
  assign t[122] = t[154] ^ x[106];
  assign t[123] = t[155] ^ x[109];
  assign t[124] = t[156] ^ x[112];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[23] & x[24]);
  assign t[132] = (x[28] & x[29]);
  assign t[133] = (x[31] & x[32]);
  assign t[134] = (x[36] & x[37]);
  assign t[135] = (x[39] & x[40]);
  assign t[136] = (x[42] & x[43]);
  assign t[137] = (x[47] & x[48]);
  assign t[138] = (x[50] & x[51]);
  assign t[139] = (x[55] & x[56]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[58] & x[59]);
  assign t[141] = (x[61] & x[62]);
  assign t[142] = (x[64] & x[65]);
  assign t[143] = (x[67] & x[68]);
  assign t[144] = (x[72] & x[73]);
  assign t[145] = (x[75] & x[76]);
  assign t[146] = (x[80] & x[81]);
  assign t[147] = (x[83] & x[84]);
  assign t[148] = (x[86] & x[87]);
  assign t[149] = (x[89] & x[90]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[92] & x[93]);
  assign t[151] = (x[95] & x[96]);
  assign t[152] = (x[98] & x[99]);
  assign t[153] = (x[101] & x[102]);
  assign t[154] = (x[104] & x[105]);
  assign t[155] = (x[107] & x[108]);
  assign t[156] = (x[110] & x[111]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[46] ? x[27] : x[26];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[40];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[100] & t[54]);
  assign t[37] = ~(t[101] & t[55]);
  assign t[38] = t[46] ? x[35] : x[34];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[42];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[65]);
  assign t[46] = ~(t[24]);
  assign t[47] = ~(t[103] & t[66]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = t[68] ? x[46] : x[45];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[46] ? x[54] : x[53];
  assign t[53] = ~(t[71] & t[72]);
  assign t[54] = ~(t[107]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = ~(t[109] & t[75]);
  assign t[58] = ~(t[110] & t[76]);
  assign t[59] = ~(t[111] & t[77]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[68] ? x[71] : x[70];
  assign t[61] = ~(t[112] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = t[17] ? x[79] : x[78];
  assign t[64] = ~(t[80] & t[81]);
  assign t[65] = ~(t[98]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[24]);
  assign t[69] = ~(t[115]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[118]);
  assign t[75] = ~(t[118] & t[86]);
  assign t[76] = ~(t[119]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[123]);
  assign t[85] = ~(t[123] & t[91]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[124]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[124] & t[92]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[121]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[25];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind173(x, y);
 input [139:0] x;
 output y;

 wire [285:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[140] ? x[78] : x[77];
  assign t[101] = ~(t[141] & t[142]);
  assign t[102] = ~(t[226]);
  assign t[103] = ~(t[215] | t[216]);
  assign t[104] = ~(t[227]);
  assign t[105] = ~(t[228]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[145] | t[146]);
  assign t[108] = ~(t[229]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[147] | t[148]);
  assign t[111] = ~(t[149] | t[150]);
  assign t[112] = ~(t[231] | t[151]);
  assign t[113] = t[29] ? x[98] : x[97];
  assign t[114] = ~(t[152] & t[153]);
  assign t[115] = ~(t[232]);
  assign t[116] = ~(t[233]);
  assign t[117] = ~(t[154] | t[155]);
  assign t[118] = t[29] ? x[106] : x[105];
  assign t[119] = ~(t[156] & t[157]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[158] & t[159]);
  assign t[121] = ~(t[160] & t[159]);
  assign t[122] = ~(x[4] & t[161]);
  assign t[123] = ~(t[162] & t[159]);
  assign t[124] = ~(t[160] & t[208]);
  assign t[125] = ~(t[80] | t[163]);
  assign t[126] = ~(t[80] | t[164]);
  assign t[127] = t[205] ? t[165] : t[123];
  assign t[128] = ~(t[78] | t[166]);
  assign t[129] = ~(t[167]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[80] | t[168]);
  assign t[131] = ~(t[234]);
  assign t[132] = ~(t[221] | t[222]);
  assign t[133] = ~(t[235]);
  assign t[134] = ~(t[236]);
  assign t[135] = ~(t[169] | t[170]);
  assign t[136] = ~(t[171] | t[126]);
  assign t[137] = ~(t[172] | t[173]);
  assign t[138] = ~(t[237]);
  assign t[139] = ~(t[224] | t[225]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[47]);
  assign t[141] = ~(t[174] | t[175]);
  assign t[142] = ~(t[176]);
  assign t[143] = ~(t[238]);
  assign t[144] = ~(t[227] | t[228]);
  assign t[145] = ~(t[30] & t[177]);
  assign t[146] = ~(t[178] & t[84]);
  assign t[147] = ~(t[239]);
  assign t[148] = ~(t[229] | t[230]);
  assign t[149] = ~(t[240]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[241]);
  assign t[151] = ~(t[179] | t[180]);
  assign t[152] = ~(t[125] | t[171]);
  assign t[153] = ~(t[181] | t[182]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[232] | t[233]);
  assign t[156] = ~(t[176] | t[50]);
  assign t[157] = ~(t[48] | t[183]);
  assign t[158] = x[4] & t[206];
  assign t[159] = ~(t[208]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(x[4] | t[206]);
  assign t[161] = ~(t[206] | t[159]);
  assign t[162] = ~(x[4] | t[184]);
  assign t[163] = t[205] ? t[185] : t[121];
  assign t[164] = t[205] ? t[120] : t[124];
  assign t[165] = ~(x[4] & t[186]);
  assign t[166] = t[205] ? t[123] : t[165];
  assign t[167] = ~(t[174] | t[126]);
  assign t[168] = t[205] ? t[187] : t[165];
  assign t[169] = ~(t[243]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = ~(t[235] | t[236]);
  assign t[171] = ~(t[80] | t[188]);
  assign t[172] = t[208] & t[189];
  assign t[173] = ~(t[190]);
  assign t[174] = ~(t[80] | t[191]);
  assign t[175] = ~(t[192] & t[190]);
  assign t[176] = ~(t[80] | t[193]);
  assign t[177] = ~(t[78] & t[194]);
  assign t[178] = ~(t[172] & t[195]);
  assign t[179] = ~(t[244]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[240] | t[241]);
  assign t[181] = t[183] | t[130];
  assign t[182] = ~(t[196] & t[84]);
  assign t[183] = ~(t[190] & t[197]);
  assign t[184] = ~(t[206]);
  assign t[185] = ~(t[158] & t[208]);
  assign t[186] = ~(t[206] | t[208]);
  assign t[187] = ~(t[208] & t[162]);
  assign t[188] = t[205] ? t[165] : t[187];
  assign t[189] = ~(t[78] | t[205]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[198] | t[128]);
  assign t[191] = t[205] ? t[122] : t[123];
  assign t[192] = ~(t[125] | t[145]);
  assign t[193] = t[205] ? t[121] : t[185];
  assign t[194] = ~(t[165] & t[187]);
  assign t[195] = t[160] | t[158];
  assign t[196] = ~(t[199] | t[174]);
  assign t[197] = ~(t[161] & t[200]);
  assign t[198] = ~(t[78] | t[201]);
  assign t[199] = ~(t[202]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[80] & t[205];
  assign t[201] = t[205] ? t[120] : t[121];
  assign t[202] = ~(t[189] & t[203]);
  assign t[203] = ~(t[187] & t[122]);
  assign t[204] = t[245] ^ x[2];
  assign t[205] = t[246] ^ x[10];
  assign t[206] = t[247] ^ x[13];
  assign t[207] = t[248] ^ x[16];
  assign t[208] = t[249] ^ x[19];
  assign t[209] = t[250] ^ x[22];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[25];
  assign t[211] = t[252] ^ x[28];
  assign t[212] = t[253] ^ x[31];
  assign t[213] = t[254] ^ x[36];
  assign t[214] = t[255] ^ x[39];
  assign t[215] = t[256] ^ x[42];
  assign t[216] = t[257] ^ x[45];
  assign t[217] = t[258] ^ x[48];
  assign t[218] = t[259] ^ x[53];
  assign t[219] = t[260] ^ x[56];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[59];
  assign t[221] = t[262] ^ x[62];
  assign t[222] = t[263] ^ x[65];
  assign t[223] = t[264] ^ x[68];
  assign t[224] = t[265] ^ x[73];
  assign t[225] = t[266] ^ x[76];
  assign t[226] = t[267] ^ x[81];
  assign t[227] = t[268] ^ x[84];
  assign t[228] = t[269] ^ x[87];
  assign t[229] = t[270] ^ x[90];
  assign t[22] = ~(t[21] ^ t[34]);
  assign t[230] = t[271] ^ x[93];
  assign t[231] = t[272] ^ x[96];
  assign t[232] = t[273] ^ x[101];
  assign t[233] = t[274] ^ x[104];
  assign t[234] = t[275] ^ x[109];
  assign t[235] = t[276] ^ x[112];
  assign t[236] = t[277] ^ x[115];
  assign t[237] = t[278] ^ x[118];
  assign t[238] = t[279] ^ x[121];
  assign t[239] = t[280] ^ x[124];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[281] ^ x[127];
  assign t[241] = t[282] ^ x[130];
  assign t[242] = t[283] ^ x[133];
  assign t[243] = t[284] ^ x[136];
  assign t[244] = t[285] ^ x[139];
  assign t[245] = (x[0] & x[1]);
  assign t[246] = (x[8] & x[9]);
  assign t[247] = (x[11] & x[12]);
  assign t[248] = (x[14] & x[15]);
  assign t[249] = (x[17] & x[18]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[20] & x[21]);
  assign t[251] = (x[23] & x[24]);
  assign t[252] = (x[26] & x[27]);
  assign t[253] = (x[29] & x[30]);
  assign t[254] = (x[34] & x[35]);
  assign t[255] = (x[37] & x[38]);
  assign t[256] = (x[40] & x[41]);
  assign t[257] = (x[43] & x[44]);
  assign t[258] = (x[46] & x[47]);
  assign t[259] = (x[51] & x[52]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[54] & x[55]);
  assign t[261] = (x[57] & x[58]);
  assign t[262] = (x[60] & x[61]);
  assign t[263] = (x[63] & x[64]);
  assign t[264] = (x[66] & x[67]);
  assign t[265] = (x[71] & x[72]);
  assign t[266] = (x[74] & x[75]);
  assign t[267] = (x[79] & x[80]);
  assign t[268] = (x[82] & x[83]);
  assign t[269] = (x[85] & x[86]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[88] & x[89]);
  assign t[271] = (x[91] & x[92]);
  assign t[272] = (x[94] & x[95]);
  assign t[273] = (x[99] & x[100]);
  assign t[274] = (x[102] & x[103]);
  assign t[275] = (x[107] & x[108]);
  assign t[276] = (x[110] & x[111]);
  assign t[277] = (x[113] & x[114]);
  assign t[278] = (x[116] & x[117]);
  assign t[279] = (x[119] & x[120]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[122] & x[123]);
  assign t[281] = (x[125] & x[126]);
  assign t[282] = (x[128] & x[129]);
  assign t[283] = (x[131] & x[132]);
  assign t[284] = (x[134] & x[135]);
  assign t[285] = (x[137] & x[138]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[209] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[37] = ~(t[61] | t[62]);
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[210] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[46] = ~(t[43] ^ t[77]);
  assign t[47] = ~(t[207]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[80] | t[82]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = ~(t[211]);
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = t[87] ? x[33] : x[32];
  assign t[56] = ~(t[88] & t[89]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[58] = ~(t[213] | t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] ^ t[96]);
  assign t[61] = ~(t[97] | t[98]);
  assign t[62] = ~(t[214] | t[99]);
  assign t[63] = ~(t[100] ^ t[101]);
  assign t[64] = ~(t[215]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[104] | t[105]);
  assign t[68] = ~(t[217] | t[106]);
  assign t[69] = t[29] ? x[50] : x[49];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[107] & t[83]);
  assign t[71] = ~(t[108] | t[109]);
  assign t[72] = ~(t[218] | t[110]);
  assign t[73] = ~(t[111] | t[112]);
  assign t[74] = ~(t[113] ^ t[114]);
  assign t[75] = ~(t[115] | t[116]);
  assign t[76] = ~(t[219] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[207]);
  assign t[79] = t[205] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[78]);
  assign t[81] = t[205] ? t[123] : t[122];
  assign t[82] = t[205] ? t[124] : t[120];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[78] | t[127];
  assign t[85] = ~(t[220]);
  assign t[86] = ~(t[211] | t[212]);
  assign t[87] = ~(t[47]);
  assign t[88] = ~(t[48] | t[128]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[221]);
  assign t[91] = ~(t[222]);
  assign t[92] = ~(t[131] | t[132]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[223] | t[135]);
  assign t[95] = t[87] ? x[70] : x[69];
  assign t[96] = ~(t[136] & t[137]);
  assign t[97] = ~(t[224]);
  assign t[98] = ~(t[225]);
  assign t[99] = ~(t[138] | t[139]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind174(x, y);
 input [151:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[107] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[108] | t[103]);
  assign t[106] = ~(t[151]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[32];
  assign t[117] = t[162] ^ x[35];
  assign t[118] = t[163] ^ x[38];
  assign t[119] = t[164] ^ x[41];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[46];
  assign t[121] = t[166] ^ x[51];
  assign t[122] = t[167] ^ x[54];
  assign t[123] = t[168] ^ x[57];
  assign t[124] = t[169] ^ x[60];
  assign t[125] = t[170] ^ x[65];
  assign t[126] = t[171] ^ x[70];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[76];
  assign t[129] = t[174] ^ x[79];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[82];
  assign t[131] = t[176] ^ x[85];
  assign t[132] = t[177] ^ x[88];
  assign t[133] = t[178] ^ x[91];
  assign t[134] = t[179] ^ x[94];
  assign t[135] = t[180] ^ x[97];
  assign t[136] = t[181] ^ x[100];
  assign t[137] = t[182] ^ x[103];
  assign t[138] = t[183] ^ x[106];
  assign t[139] = t[184] ^ x[109];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[112];
  assign t[141] = t[186] ^ x[115];
  assign t[142] = t[187] ^ x[118];
  assign t[143] = t[188] ^ x[121];
  assign t[144] = t[189] ^ x[124];
  assign t[145] = t[190] ^ x[127];
  assign t[146] = t[191] ^ x[130];
  assign t[147] = t[192] ^ x[133];
  assign t[148] = t[193] ^ x[136];
  assign t[149] = t[194] ^ x[139];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[142];
  assign t[151] = t[196] ^ x[145];
  assign t[152] = t[197] ^ x[148];
  assign t[153] = t[198] ^ x[151];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[30] & x[31]);
  assign t[162] = (x[33] & x[34]);
  assign t[163] = (x[36] & x[37]);
  assign t[164] = (x[39] & x[40]);
  assign t[165] = (x[44] & x[45]);
  assign t[166] = (x[49] & x[50]);
  assign t[167] = (x[52] & x[53]);
  assign t[168] = (x[55] & x[56]);
  assign t[169] = (x[58] & x[59]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[63] & x[64]);
  assign t[171] = (x[68] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[74] & x[75]);
  assign t[174] = (x[77] & x[78]);
  assign t[175] = (x[80] & x[81]);
  assign t[176] = (x[83] & x[84]);
  assign t[177] = (x[86] & x[87]);
  assign t[178] = (x[89] & x[90]);
  assign t[179] = (x[92] & x[93]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[95] & x[96]);
  assign t[181] = (x[98] & x[99]);
  assign t[182] = (x[101] & x[102]);
  assign t[183] = (x[104] & x[105]);
  assign t[184] = (x[107] & x[108]);
  assign t[185] = (x[110] & x[111]);
  assign t[186] = (x[113] & x[114]);
  assign t[187] = (x[116] & x[117]);
  assign t[188] = (x[119] & x[120]);
  assign t[189] = (x[122] & x[123]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[125] & x[126]);
  assign t[191] = (x[128] & x[129]);
  assign t[192] = (x[131] & x[132]);
  assign t[193] = (x[134] & x[135]);
  assign t[194] = (x[137] & x[138]);
  assign t[195] = (x[140] & x[141]);
  assign t[196] = (x[143] & x[144]);
  assign t[197] = (x[146] & x[147]);
  assign t[198] = (x[149] & x[150]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[56];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = t[59] | t[115];
  assign t[39] = t[60] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[41];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = t[73] | t[118];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = t[76] | t[119];
  assign t[52] = t[77] ? x[43] : x[42];
  assign t[53] = ~(t[78] & t[79]);
  assign t[54] = t[80] | t[120];
  assign t[55] = t[77] ? x[48] : x[47];
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[121]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[83] | t[57]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[24]);
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = t[86] | t[123];
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = t[89] | t[124];
  assign t[65] = t[17] ? x[62] : x[61];
  assign t[66] = ~(t[90] & t[91]);
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = t[94] | t[125];
  assign t[69] = t[17] ? x[67] : x[66];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[24]);
  assign t[78] = ~(t[131]);
  assign t[79] = ~(t[132]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[97] | t[78]);
  assign t[81] = ~(t[98] & t[99]);
  assign t[82] = t[100] | t[133];
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[101] | t[84]);
  assign t[87] = ~(t[137]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[102] | t[87]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[103] & t[104]);
  assign t[91] = t[105] | t[139];
  assign t[92] = ~(t[140]);
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[106] | t[92]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind175(x, y);
 input [151:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[155]);
  assign t[104] = ~(t[114] & t[115]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[116] & t[117]);
  assign t[112] = ~(t[150] & t[149]);
  assign t[113] = ~(t[160]);
  assign t[114] = ~(t[155] & t[154]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[159] & t[158]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[32];
  assign t[126] = t[171] ^ x[35];
  assign t[127] = t[172] ^ x[38];
  assign t[128] = t[173] ^ x[41];
  assign t[129] = t[174] ^ x[46];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[51];
  assign t[131] = t[176] ^ x[54];
  assign t[132] = t[177] ^ x[57];
  assign t[133] = t[178] ^ x[60];
  assign t[134] = t[179] ^ x[65];
  assign t[135] = t[180] ^ x[70];
  assign t[136] = t[181] ^ x[73];
  assign t[137] = t[182] ^ x[76];
  assign t[138] = t[183] ^ x[79];
  assign t[139] = t[184] ^ x[82];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[85];
  assign t[141] = t[186] ^ x[88];
  assign t[142] = t[187] ^ x[91];
  assign t[143] = t[188] ^ x[94];
  assign t[144] = t[189] ^ x[97];
  assign t[145] = t[190] ^ x[100];
  assign t[146] = t[191] ^ x[103];
  assign t[147] = t[192] ^ x[106];
  assign t[148] = t[193] ^ x[109];
  assign t[149] = t[194] ^ x[112];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[118];
  assign t[152] = t[197] ^ x[121];
  assign t[153] = t[198] ^ x[124];
  assign t[154] = t[199] ^ x[127];
  assign t[155] = t[200] ^ x[130];
  assign t[156] = t[201] ^ x[133];
  assign t[157] = t[202] ^ x[136];
  assign t[158] = t[203] ^ x[139];
  assign t[159] = t[204] ^ x[142];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[145];
  assign t[161] = t[206] ^ x[148];
  assign t[162] = t[207] ^ x[151];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[30] & x[31]);
  assign t[171] = (x[33] & x[34]);
  assign t[172] = (x[36] & x[37]);
  assign t[173] = (x[39] & x[40]);
  assign t[174] = (x[44] & x[45]);
  assign t[175] = (x[49] & x[50]);
  assign t[176] = (x[52] & x[53]);
  assign t[177] = (x[55] & x[56]);
  assign t[178] = (x[58] & x[59]);
  assign t[179] = (x[63] & x[64]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[68] & x[69]);
  assign t[181] = (x[71] & x[72]);
  assign t[182] = (x[74] & x[75]);
  assign t[183] = (x[77] & x[78]);
  assign t[184] = (x[80] & x[81]);
  assign t[185] = (x[83] & x[84]);
  assign t[186] = (x[86] & x[87]);
  assign t[187] = (x[89] & x[90]);
  assign t[188] = (x[92] & x[93]);
  assign t[189] = (x[95] & x[96]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[98] & x[99]);
  assign t[191] = (x[101] & x[102]);
  assign t[192] = (x[104] & x[105]);
  assign t[193] = (x[107] & x[108]);
  assign t[194] = (x[110] & x[111]);
  assign t[195] = (x[113] & x[114]);
  assign t[196] = (x[116] & x[117]);
  assign t[197] = (x[119] & x[120]);
  assign t[198] = (x[122] & x[123]);
  assign t[199] = (x[125] & x[126]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[128] & x[129]);
  assign t[201] = (x[131] & x[132]);
  assign t[202] = (x[134] & x[135]);
  assign t[203] = (x[137] & x[138]);
  assign t[204] = (x[140] & x[141]);
  assign t[205] = (x[143] & x[144]);
  assign t[206] = (x[146] & x[147]);
  assign t[207] = (x[149] & x[150]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[56];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = ~(t[59] & t[124]);
  assign t[39] = t[60] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[41];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[74] & t[127]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[75] & t[76]);
  assign t[51] = ~(t[77] & t[128]);
  assign t[52] = t[60] ? x[43] : x[42];
  assign t[53] = ~(t[78] & t[79]);
  assign t[54] = ~(t[80] & t[129]);
  assign t[55] = t[60] ? x[48] : x[47];
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[130]);
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[83] & t[84]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[24]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[132]);
  assign t[63] = ~(t[88] & t[89]);
  assign t[64] = ~(t[90] & t[133]);
  assign t[65] = t[17] ? x[62] : x[61];
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[94]);
  assign t[68] = ~(t[95] & t[134]);
  assign t[69] = t[121] ? x[67] : x[66];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126] & t[125]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[96] & t[97]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[98] & t[99]);
  assign t[78] = ~(t[140]);
  assign t[79] = ~(t[141]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[100] & t[101]);
  assign t[81] = ~(t[102] & t[103]);
  assign t[82] = ~(t[104] & t[142]);
  assign t[83] = ~(t[131] & t[130]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[105] & t[106]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[107] & t[108]);
  assign t[91] = ~(t[109] & t[110]);
  assign t[92] = ~(t[111] & t[148]);
  assign t[93] = ~(t[149]);
  assign t[94] = ~(t[150]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind176(x, y);
 input [121:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[25];
  assign t[106] = t[141] ^ x[30];
  assign t[107] = t[142] ^ x[33];
  assign t[108] = t[143] ^ x[38];
  assign t[109] = t[144] ^ x[41];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[44];
  assign t[111] = t[146] ^ x[47];
  assign t[112] = t[147] ^ x[50];
  assign t[113] = t[148] ^ x[55];
  assign t[114] = t[149] ^ x[58];
  assign t[115] = t[150] ^ x[63];
  assign t[116] = t[151] ^ x[66];
  assign t[117] = t[152] ^ x[69];
  assign t[118] = t[153] ^ x[72];
  assign t[119] = t[154] ^ x[75];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[155] ^ x[80];
  assign t[121] = t[156] ^ x[83];
  assign t[122] = t[157] ^ x[88];
  assign t[123] = t[158] ^ x[91];
  assign t[124] = t[159] ^ x[94];
  assign t[125] = t[160] ^ x[97];
  assign t[126] = t[161] ^ x[100];
  assign t[127] = t[162] ^ x[103];
  assign t[128] = t[163] ^ x[106];
  assign t[129] = t[164] ^ x[109];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[112];
  assign t[131] = t[166] ^ x[115];
  assign t[132] = t[167] ^ x[118];
  assign t[133] = t[168] ^ x[121];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[23] & x[24]);
  assign t[141] = (x[28] & x[29]);
  assign t[142] = (x[31] & x[32]);
  assign t[143] = (x[36] & x[37]);
  assign t[144] = (x[39] & x[40]);
  assign t[145] = (x[42] & x[43]);
  assign t[146] = (x[45] & x[46]);
  assign t[147] = (x[48] & x[49]);
  assign t[148] = (x[53] & x[54]);
  assign t[149] = (x[56] & x[57]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[61] & x[62]);
  assign t[151] = (x[64] & x[65]);
  assign t[152] = (x[67] & x[68]);
  assign t[153] = (x[70] & x[71]);
  assign t[154] = (x[73] & x[74]);
  assign t[155] = (x[78] & x[79]);
  assign t[156] = (x[81] & x[82]);
  assign t[157] = (x[86] & x[87]);
  assign t[158] = (x[89] & x[90]);
  assign t[159] = (x[92] & x[93]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[95] & x[96]);
  assign t[161] = (x[98] & x[99]);
  assign t[162] = (x[101] & x[102]);
  assign t[163] = (x[104] & x[105]);
  assign t[164] = (x[107] & x[108]);
  assign t[165] = (x[110] & x[111]);
  assign t[166] = (x[113] & x[114]);
  assign t[167] = (x[116] & x[117]);
  assign t[168] = (x[119] & x[120]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[27] : x[26];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[33];
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = t[47] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[43];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[68]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[73] ? x[52] : x[51];
  assign t[53] = ~(t[74] & t[75]);
  assign t[54] = ~(t[113] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = t[73] ? x[60] : x[59];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[73] ? x[77] : x[76];
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = ~(t[121] & t[84]);
  assign t[66] = t[47] ? x[85] : x[84];
  assign t[67] = ~(t[85] & t[86]);
  assign t[68] = ~(t[104]);
  assign t[69] = ~(t[122]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[24]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[132] & t[97]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[120]);
  assign t[95] = ~(t[133]);
  assign t[96] = ~(t[133] & t[98]);
  assign t[97] = ~(t[124]);
  assign t[98] = ~(t[130]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind177(x, y);
 input [151:0] x;
 output y;

 wire [293:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[226]);
  assign t[101] = ~(t[227]);
  assign t[102] = ~(t[145] | t[146]);
  assign t[103] = ~(t[147] | t[148]);
  assign t[104] = ~(t[228] | t[149]);
  assign t[105] = t[142] ? x[87] : x[86];
  assign t[106] = ~(t[150] & t[151]);
  assign t[107] = ~(t[229]);
  assign t[108] = ~(t[216] | t[217]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[152] | t[153]);
  assign t[112] = ~(t[154] | t[155]);
  assign t[113] = ~(t[232]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[156] | t[157]);
  assign t[116] = ~(t[158] | t[159]);
  assign t[117] = ~(t[234] | t[160]);
  assign t[118] = t[29] ? x[107] : x[106];
  assign t[119] = ~(t[161] & t[162]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[235]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[163] | t[164]);
  assign t[123] = t[29] ? x[115] : x[114];
  assign t[124] = ~(t[165] & t[166]);
  assign t[125] = ~(t[127] | t[167]);
  assign t[126] = ~(t[85] | t[168]);
  assign t[127] = ~(t[207]);
  assign t[128] = ~(t[169] & t[170]);
  assign t[129] = t[208] & t[171];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[172] | t[173];
  assign t[131] = t[205] ? t[169] : t[174];
  assign t[132] = ~(t[172] & t[175]);
  assign t[133] = ~(t[173] & t[208]);
  assign t[134] = ~(t[172] & t[208]);
  assign t[135] = ~(t[173] & t[175]);
  assign t[136] = ~(t[237]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[206] | t[175]);
  assign t[139] = t[85] & t[205];
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[238]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[48]);
  assign t[143] = ~(t[176] & t[94]);
  assign t[144] = ~(t[85] | t[177]);
  assign t[145] = ~(t[239]);
  assign t[146] = ~(t[226] | t[227]);
  assign t[147] = ~(t[240]);
  assign t[148] = ~(t[241]);
  assign t[149] = ~(t[178] | t[179]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[51]);
  assign t[151] = ~(t[180] | t[144]);
  assign t[152] = ~(t[242]);
  assign t[153] = ~(t[230] | t[231]);
  assign t[154] = ~(t[85] | t[181]);
  assign t[155] = ~(t[31] & t[84]);
  assign t[156] = ~(t[243]);
  assign t[157] = ~(t[232] | t[233]);
  assign t[158] = ~(t[244]);
  assign t[159] = ~(t[245]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(t[182] | t[183]);
  assign t[161] = ~(t[51] | t[184]);
  assign t[162] = ~(t[99] | t[185]);
  assign t[163] = ~(t[246]);
  assign t[164] = ~(t[235] | t[236]);
  assign t[165] = ~(t[186] | t[154]);
  assign t[166] = ~(t[125] | t[143]);
  assign t[167] = t[205] ? t[132] : t[135];
  assign t[168] = t[205] ? t[174] : t[187];
  assign t[169] = ~(x[4] & t[188]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = ~(t[208] & t[189]);
  assign t[171] = ~(t[127] | t[205]);
  assign t[172] = ~(x[4] | t[206]);
  assign t[173] = x[4] & t[206];
  assign t[174] = ~(t[189] & t[175]);
  assign t[175] = ~(t[208]);
  assign t[176] = ~(t[190] | t[191]);
  assign t[177] = t[205] ? t[170] : t[169];
  assign t[178] = ~(t[247]);
  assign t[179] = ~(t[240] | t[241]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[192]);
  assign t[181] = t[205] ? t[134] : t[135];
  assign t[182] = ~(t[248]);
  assign t[183] = ~(t[244] | t[245]);
  assign t[184] = ~(t[85] | t[193]);
  assign t[185] = ~(t[194] & t[84]);
  assign t[186] = ~(t[85] | t[195]);
  assign t[187] = ~(x[4] & t[138]);
  assign t[188] = ~(t[206] | t[208]);
  assign t[189] = ~(x[4] | t[196]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[127] | t[197]);
  assign t[191] = ~(t[127] | t[198]);
  assign t[192] = ~(t[199] | t[52]);
  assign t[193] = t[205] ? t[169] : t[170];
  assign t[194] = ~(t[200] | t[199]);
  assign t[195] = t[205] ? t[132] : t[133];
  assign t[196] = ~(t[206]);
  assign t[197] = t[205] ? t[135] : t[132];
  assign t[198] = t[205] ? t[174] : t[169];
  assign t[199] = ~(t[85] | t[201]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[202]);
  assign t[201] = t[205] ? t[187] : t[174];
  assign t[202] = ~(t[171] & t[203]);
  assign t[203] = ~(t[170] & t[187]);
  assign t[204] = t[249] ^ x[2];
  assign t[205] = t[250] ^ x[10];
  assign t[206] = t[251] ^ x[13];
  assign t[207] = t[252] ^ x[16];
  assign t[208] = t[253] ^ x[19];
  assign t[209] = t[254] ^ x[22];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[25];
  assign t[211] = t[256] ^ x[28];
  assign t[212] = t[257] ^ x[31];
  assign t[213] = t[258] ^ x[34];
  assign t[214] = t[259] ^ x[39];
  assign t[215] = t[260] ^ x[42];
  assign t[216] = t[261] ^ x[45];
  assign t[217] = t[262] ^ x[48];
  assign t[218] = t[263] ^ x[51];
  assign t[219] = t[264] ^ x[56];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[59];
  assign t[221] = t[266] ^ x[62];
  assign t[222] = t[267] ^ x[65];
  assign t[223] = t[268] ^ x[68];
  assign t[224] = t[269] ^ x[71];
  assign t[225] = t[270] ^ x[74];
  assign t[226] = t[271] ^ x[79];
  assign t[227] = t[272] ^ x[82];
  assign t[228] = t[273] ^ x[85];
  assign t[229] = t[274] ^ x[90];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[93];
  assign t[231] = t[276] ^ x[96];
  assign t[232] = t[277] ^ x[99];
  assign t[233] = t[278] ^ x[102];
  assign t[234] = t[279] ^ x[105];
  assign t[235] = t[280] ^ x[110];
  assign t[236] = t[281] ^ x[113];
  assign t[237] = t[282] ^ x[118];
  assign t[238] = t[283] ^ x[121];
  assign t[239] = t[284] ^ x[124];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[127];
  assign t[241] = t[286] ^ x[130];
  assign t[242] = t[287] ^ x[133];
  assign t[243] = t[288] ^ x[136];
  assign t[244] = t[289] ^ x[139];
  assign t[245] = t[290] ^ x[142];
  assign t[246] = t[291] ^ x[145];
  assign t[247] = t[292] ^ x[148];
  assign t[248] = t[293] ^ x[151];
  assign t[249] = (x[0] & x[1]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[8] & x[9]);
  assign t[251] = (x[11] & x[12]);
  assign t[252] = (x[14] & x[15]);
  assign t[253] = (x[17] & x[18]);
  assign t[254] = (x[20] & x[21]);
  assign t[255] = (x[23] & x[24]);
  assign t[256] = (x[26] & x[27]);
  assign t[257] = (x[29] & x[30]);
  assign t[258] = (x[32] & x[33]);
  assign t[259] = (x[37] & x[38]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[40] & x[41]);
  assign t[261] = (x[43] & x[44]);
  assign t[262] = (x[46] & x[47]);
  assign t[263] = (x[49] & x[50]);
  assign t[264] = (x[54] & x[55]);
  assign t[265] = (x[57] & x[58]);
  assign t[266] = (x[60] & x[61]);
  assign t[267] = (x[63] & x[64]);
  assign t[268] = (x[66] & x[67]);
  assign t[269] = (x[69] & x[70]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[72] & x[73]);
  assign t[271] = (x[77] & x[78]);
  assign t[272] = (x[80] & x[81]);
  assign t[273] = (x[83] & x[84]);
  assign t[274] = (x[88] & x[89]);
  assign t[275] = (x[91] & x[92]);
  assign t[276] = (x[94] & x[95]);
  assign t[277] = (x[97] & x[98]);
  assign t[278] = (x[100] & x[101]);
  assign t[279] = (x[103] & x[104]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[108] & x[109]);
  assign t[281] = (x[111] & x[112]);
  assign t[282] = (x[116] & x[117]);
  assign t[283] = (x[119] & x[120]);
  assign t[284] = (x[122] & x[123]);
  assign t[285] = (x[125] & x[126]);
  assign t[286] = (x[128] & x[129]);
  assign t[287] = (x[131] & x[132]);
  assign t[288] = (x[134] & x[135]);
  assign t[289] = (x[137] & x[138]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[140] & x[141]);
  assign t[291] = (x[143] & x[144]);
  assign t[292] = (x[146] & x[147]);
  assign t[293] = (x[149] & x[150]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[209] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[38] ^ t[62]);
  assign t[38] = ~(t[63] | t[64]);
  assign t[39] = ~(t[65] ^ t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[67] | t[68]);
  assign t[41] = ~(t[210] | t[69]);
  assign t[42] = ~(t[70] | t[71]);
  assign t[43] = ~(t[72] ^ t[73]);
  assign t[44] = ~(t[74] | t[75]);
  assign t[45] = ~(t[76] ^ t[77]);
  assign t[46] = ~(t[78] | t[79]);
  assign t[47] = ~(t[44] ^ t[80]);
  assign t[48] = ~(t[207]);
  assign t[49] = ~(t[81] & t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[83] & t[84]);
  assign t[51] = ~(t[85] | t[86]);
  assign t[52] = ~(t[85] | t[87]);
  assign t[53] = ~(t[211]);
  assign t[54] = ~(t[212]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[213] | t[92]);
  assign t[58] = t[29] ? x[36] : x[35];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[214] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[100] | t[101]);
  assign t[64] = ~(t[215] | t[102]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[66] = ~(t[105] ^ t[106]);
  assign t[67] = ~(t[216]);
  assign t[68] = ~(t[217]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[109] | t[110]);
  assign t[71] = ~(t[218] | t[111]);
  assign t[72] = t[29] ? x[53] : x[52];
  assign t[73] = ~(t[81] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[219] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[220] | t[122]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[123] ^ t[124]);
  assign t[81] = ~(t[125] | t[126]);
  assign t[82] = ~(t[127] & t[128]);
  assign t[83] = ~(t[129] & t[130]);
  assign t[84] = t[127] | t[131];
  assign t[85] = ~(t[127]);
  assign t[86] = t[205] ? t[133] : t[132];
  assign t[87] = t[205] ? t[135] : t[134];
  assign t[88] = ~(t[221]);
  assign t[89] = ~(t[211] | t[212]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[222]);
  assign t[91] = ~(t[223]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[51] | t[49]);
  assign t[94] = ~(t[138] & t[139]);
  assign t[95] = ~(t[224]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[140] | t[141]);
  assign t[98] = t[142] ? x[76] : x[75];
  assign t[99] = t[143] | t[144];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind178(x, y);
 input [139:0] x;
 output y;

 wire [180:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[141] ^ x[8];
  assign t[101] = t[142] ^ x[11];
  assign t[102] = t[143] ^ x[14];
  assign t[103] = t[144] ^ x[17];
  assign t[104] = t[145] ^ x[22];
  assign t[105] = t[146] ^ x[27];
  assign t[106] = t[147] ^ x[32];
  assign t[107] = t[148] ^ x[35];
  assign t[108] = t[149] ^ x[38];
  assign t[109] = t[150] ^ x[41];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[46];
  assign t[111] = t[152] ^ x[51];
  assign t[112] = t[153] ^ x[54];
  assign t[113] = t[154] ^ x[57];
  assign t[114] = t[155] ^ x[62];
  assign t[115] = t[156] ^ x[67];
  assign t[116] = t[157] ^ x[70];
  assign t[117] = t[158] ^ x[73];
  assign t[118] = t[159] ^ x[76];
  assign t[119] = t[160] ^ x[79];
  assign t[11] = t[102] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[82];
  assign t[121] = t[162] ^ x[85];
  assign t[122] = t[163] ^ x[88];
  assign t[123] = t[164] ^ x[91];
  assign t[124] = t[165] ^ x[94];
  assign t[125] = t[166] ^ x[97];
  assign t[126] = t[167] ^ x[100];
  assign t[127] = t[168] ^ x[103];
  assign t[128] = t[169] ^ x[106];
  assign t[129] = t[170] ^ x[109];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[112];
  assign t[131] = t[172] ^ x[115];
  assign t[132] = t[173] ^ x[118];
  assign t[133] = t[174] ^ x[121];
  assign t[134] = t[175] ^ x[124];
  assign t[135] = t[176] ^ x[127];
  assign t[136] = t[177] ^ x[130];
  assign t[137] = t[178] ^ x[133];
  assign t[138] = t[179] ^ x[136];
  assign t[139] = t[180] ^ x[139];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[0] & x[1]);
  assign t[141] = (x[6] & x[7]);
  assign t[142] = (x[9] & x[10]);
  assign t[143] = (x[12] & x[13]);
  assign t[144] = (x[15] & x[16]);
  assign t[145] = (x[20] & x[21]);
  assign t[146] = (x[25] & x[26]);
  assign t[147] = (x[30] & x[31]);
  assign t[148] = (x[33] & x[34]);
  assign t[149] = (x[36] & x[37]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[39] & x[40]);
  assign t[151] = (x[44] & x[45]);
  assign t[152] = (x[49] & x[50]);
  assign t[153] = (x[52] & x[53]);
  assign t[154] = (x[55] & x[56]);
  assign t[155] = (x[60] & x[61]);
  assign t[156] = (x[65] & x[66]);
  assign t[157] = (x[68] & x[69]);
  assign t[158] = (x[71] & x[72]);
  assign t[159] = (x[74] & x[75]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[77] & x[78]);
  assign t[161] = (x[80] & x[81]);
  assign t[162] = (x[83] & x[84]);
  assign t[163] = (x[86] & x[87]);
  assign t[164] = (x[89] & x[90]);
  assign t[165] = (x[92] & x[93]);
  assign t[166] = (x[95] & x[96]);
  assign t[167] = (x[98] & x[99]);
  assign t[168] = (x[101] & x[102]);
  assign t[169] = (x[104] & x[105]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[107] & x[108]);
  assign t[171] = (x[110] & x[111]);
  assign t[172] = (x[113] & x[114]);
  assign t[173] = (x[116] & x[117]);
  assign t[174] = (x[119] & x[120]);
  assign t[175] = (x[122] & x[123]);
  assign t[176] = (x[125] & x[126]);
  assign t[177] = (x[128] & x[129]);
  assign t[178] = (x[131] & x[132]);
  assign t[179] = (x[134] & x[135]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[137] & x[138]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = t[42] | t[104];
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = ~(t[46] & t[47]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[48] ^ t[36];
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[29];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = t[54] | t[105];
  assign t[35] = t[102] ? x[29] : x[28];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[106]);
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[63] | t[40]);
  assign t[43] = ~(t[64]);
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] | t[108];
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = t[70] | t[109];
  assign t[48] = t[43] ? x[43] : x[42];
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[73] | t[110];
  assign t[51] = t[43] ? x[48] : x[47];
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[74] | t[52]);
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = t[77] | t[113];
  assign t[57] = t[102] ? x[59] : x[58];
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = t[82] | t[114];
  assign t[61] = t[83] ? x[64] : x[63];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[115]);
  assign t[64] = ~(t[102]);
  assign t[65] = ~(t[116]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[86] | t[65]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = ~(t[100] & t[101]);
  assign t[70] = ~(t[87] | t[68]);
  assign t[71] = ~(t[120]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[88] | t[71]);
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[89] | t[75]);
  assign t[78] = ~(t[90] & t[91]);
  assign t[79] = t[92] | t[125];
  assign t[7] = ~(t[102] & t[103]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[93] | t[80]);
  assign t[83] = ~(t[64]);
  assign t[84] = ~(t[94] & t[95]);
  assign t[85] = t[96] | t[128];
  assign t[86] = ~(t[129]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[97] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[98] | t[94]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = t[140] ^ x[2];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind179(x, y);
 input [139:0] x;
 output y;

 wire [188:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[144]);
  assign t[101] = ~(t[145]);
  assign t[102] = ~(t[105] & t[106]);
  assign t[103] = ~(t[142] & t[141]);
  assign t[104] = ~(t[146]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[147]);
  assign t[107] = t[148] ^ x[2];
  assign t[108] = t[149] ^ x[8];
  assign t[109] = t[150] ^ x[11];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[14];
  assign t[111] = t[152] ^ x[17];
  assign t[112] = t[153] ^ x[22];
  assign t[113] = t[154] ^ x[27];
  assign t[114] = t[155] ^ x[32];
  assign t[115] = t[156] ^ x[35];
  assign t[116] = t[157] ^ x[38];
  assign t[117] = t[158] ^ x[41];
  assign t[118] = t[159] ^ x[46];
  assign t[119] = t[160] ^ x[51];
  assign t[11] = t[110] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[54];
  assign t[121] = t[162] ^ x[57];
  assign t[122] = t[163] ^ x[62];
  assign t[123] = t[164] ^ x[67];
  assign t[124] = t[165] ^ x[70];
  assign t[125] = t[166] ^ x[73];
  assign t[126] = t[167] ^ x[76];
  assign t[127] = t[168] ^ x[79];
  assign t[128] = t[169] ^ x[82];
  assign t[129] = t[170] ^ x[85];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[88];
  assign t[131] = t[172] ^ x[91];
  assign t[132] = t[173] ^ x[94];
  assign t[133] = t[174] ^ x[97];
  assign t[134] = t[175] ^ x[100];
  assign t[135] = t[176] ^ x[103];
  assign t[136] = t[177] ^ x[106];
  assign t[137] = t[178] ^ x[109];
  assign t[138] = t[179] ^ x[112];
  assign t[139] = t[180] ^ x[115];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = t[181] ^ x[118];
  assign t[141] = t[182] ^ x[121];
  assign t[142] = t[183] ^ x[124];
  assign t[143] = t[184] ^ x[127];
  assign t[144] = t[185] ^ x[130];
  assign t[145] = t[186] ^ x[133];
  assign t[146] = t[187] ^ x[136];
  assign t[147] = t[188] ^ x[139];
  assign t[148] = (x[0] & x[1]);
  assign t[149] = (x[6] & x[7]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[9] & x[10]);
  assign t[151] = (x[12] & x[13]);
  assign t[152] = (x[15] & x[16]);
  assign t[153] = (x[20] & x[21]);
  assign t[154] = (x[25] & x[26]);
  assign t[155] = (x[30] & x[31]);
  assign t[156] = (x[33] & x[34]);
  assign t[157] = (x[36] & x[37]);
  assign t[158] = (x[39] & x[40]);
  assign t[159] = (x[44] & x[45]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[49] & x[50]);
  assign t[161] = (x[52] & x[53]);
  assign t[162] = (x[55] & x[56]);
  assign t[163] = (x[60] & x[61]);
  assign t[164] = (x[65] & x[66]);
  assign t[165] = (x[68] & x[69]);
  assign t[166] = (x[71] & x[72]);
  assign t[167] = (x[74] & x[75]);
  assign t[168] = (x[77] & x[78]);
  assign t[169] = (x[80] & x[81]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[83] & x[84]);
  assign t[171] = (x[86] & x[87]);
  assign t[172] = (x[89] & x[90]);
  assign t[173] = (x[92] & x[93]);
  assign t[174] = (x[95] & x[96]);
  assign t[175] = (x[98] & x[99]);
  assign t[176] = (x[101] & x[102]);
  assign t[177] = (x[104] & x[105]);
  assign t[178] = (x[107] & x[108]);
  assign t[179] = (x[110] & x[111]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[113] & x[114]);
  assign t[181] = (x[116] & x[117]);
  assign t[182] = (x[119] & x[120]);
  assign t[183] = (x[122] & x[123]);
  assign t[184] = (x[125] & x[126]);
  assign t[185] = (x[128] & x[129]);
  assign t[186] = (x[131] & x[132]);
  assign t[187] = (x[134] & x[135]);
  assign t[188] = (x[137] & x[138]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = ~(t[42] & t[112]);
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = ~(t[46] & t[47]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[48] ^ t[36];
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[29];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = ~(t[54] & t[113]);
  assign t[35] = t[110] ? x[29] : x[28];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[114]);
  assign t[41] = ~(t[115]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = ~(t[65]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = ~(t[68] & t[116]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[117]);
  assign t[48] = t[43] ? x[43] : x[42];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[74] & t[118]);
  assign t[51] = t[110] ? x[48] : x[47];
  assign t[52] = ~(t[119]);
  assign t[53] = ~(t[120]);
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[79] & t[121]);
  assign t[57] = t[110] ? x[59] : x[58];
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[84] & t[122]);
  assign t[61] = t[43] ? x[64] : x[63];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[115] & t[114]);
  assign t[64] = ~(t[123]);
  assign t[65] = ~(t[110]);
  assign t[66] = ~(t[124]);
  assign t[67] = ~(t[125]);
  assign t[68] = ~(t[87] & t[88]);
  assign t[69] = ~(t[126]);
  assign t[6] = ~(t[108] & t[109]);
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[89] & t[90]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[91] & t[92]);
  assign t[75] = ~(t[120] & t[119]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[93] & t[94]);
  assign t[7] = ~(t[110] & t[111]);
  assign t[80] = ~(t[95] & t[96]);
  assign t[81] = ~(t[97] & t[133]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[98] & t[99]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[136]);
  assign t[87] = ~(t[125] & t[124]);
  assign t[88] = ~(t[137]);
  assign t[89] = ~(t[127] & t[126]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[139]);
  assign t[93] = ~(t[132] & t[131]);
  assign t[94] = ~(t[140]);
  assign t[95] = ~(t[141]);
  assign t[96] = ~(t[142]);
  assign t[97] = ~(t[103] & t[104]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[143]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[107];
endmodule

module R1ind180(x, y);
 input [112:0] x;
 output y;

 wire [154:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[132] ^ x[38];
  assign t[101] = t[133] ^ x[41];
  assign t[102] = t[134] ^ x[44];
  assign t[103] = t[135] ^ x[47];
  assign t[104] = t[136] ^ x[50];
  assign t[105] = t[137] ^ x[55];
  assign t[106] = t[138] ^ x[58];
  assign t[107] = t[139] ^ x[63];
  assign t[108] = t[140] ^ x[66];
  assign t[109] = t[141] ^ x[69];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[142] ^ x[74];
  assign t[111] = t[143] ^ x[77];
  assign t[112] = t[144] ^ x[82];
  assign t[113] = t[145] ^ x[85];
  assign t[114] = t[146] ^ x[88];
  assign t[115] = t[147] ^ x[91];
  assign t[116] = t[148] ^ x[94];
  assign t[117] = t[149] ^ x[97];
  assign t[118] = t[150] ^ x[100];
  assign t[119] = t[151] ^ x[103];
  assign t[11] = t[94] ? x[18] : x[19];
  assign t[120] = t[152] ^ x[106];
  assign t[121] = t[153] ^ x[109];
  assign t[122] = t[154] ^ x[112];
  assign t[123] = (x[0] & x[1]);
  assign t[124] = (x[6] & x[7]);
  assign t[125] = (x[9] & x[10]);
  assign t[126] = (x[12] & x[13]);
  assign t[127] = (x[15] & x[16]);
  assign t[128] = (x[20] & x[21]);
  assign t[129] = (x[23] & x[24]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = (x[28] & x[29]);
  assign t[131] = (x[31] & x[32]);
  assign t[132] = (x[36] & x[37]);
  assign t[133] = (x[39] & x[40]);
  assign t[134] = (x[42] & x[43]);
  assign t[135] = (x[45] & x[46]);
  assign t[136] = (x[48] & x[49]);
  assign t[137] = (x[53] & x[54]);
  assign t[138] = (x[56] & x[57]);
  assign t[139] = (x[61] & x[62]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[64] & x[65]);
  assign t[141] = (x[67] & x[68]);
  assign t[142] = (x[72] & x[73]);
  assign t[143] = (x[75] & x[76]);
  assign t[144] = (x[80] & x[81]);
  assign t[145] = (x[83] & x[84]);
  assign t[146] = (x[86] & x[87]);
  assign t[147] = (x[89] & x[90]);
  assign t[148] = (x[92] & x[93]);
  assign t[149] = (x[95] & x[96]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[98] & x[99]);
  assign t[151] = (x[101] & x[102]);
  assign t[152] = (x[104] & x[105]);
  assign t[153] = (x[107] & x[108]);
  assign t[154] = (x[110] & x[111]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[96] & t[40]);
  assign t[26] = ~(t[97] & t[41]);
  assign t[27] = t[42] ? x[27] : x[26];
  assign t[28] = ~(t[43] & t[44]);
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[47] ^ t[31];
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[36];
  assign t[33] = ~(t[98] & t[51]);
  assign t[34] = ~(t[99] & t[52]);
  assign t[35] = t[94] ? x[35] : x[34];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[56];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[100]);
  assign t[41] = ~(t[100] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[101] & t[63]);
  assign t[44] = ~(t[102] & t[64]);
  assign t[45] = ~(t[103] & t[65]);
  assign t[46] = ~(t[104] & t[66]);
  assign t[47] = t[67] ? x[52] : x[51];
  assign t[48] = ~(t[105] & t[68]);
  assign t[49] = ~(t[106] & t[69]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[70] ? x[60] : x[59];
  assign t[51] = ~(t[107]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = t[94] ? x[71] : x[70];
  assign t[56] = ~(t[74] & t[75]);
  assign t[57] = ~(t[110] & t[76]);
  assign t[58] = ~(t[111] & t[77]);
  assign t[59] = t[42] ? x[79] : x[78];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[78] & t[79]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[94]);
  assign t[63] = ~(t[112]);
  assign t[64] = ~(t[112] & t[80]);
  assign t[65] = ~(t[113]);
  assign t[66] = ~(t[113] & t[81]);
  assign t[67] = ~(t[62]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = ~(t[92] & t[93]);
  assign t[70] = ~(t[62]);
  assign t[71] = ~(t[98]);
  assign t[72] = ~(t[115]);
  assign t[73] = ~(t[115] & t[83]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[94] & t[95]);
  assign t[80] = ~(t[101]);
  assign t[81] = ~(t[103]);
  assign t[82] = ~(t[105]);
  assign t[83] = ~(t[108]);
  assign t[84] = ~(t[121]);
  assign t[85] = ~(t[121] & t[89]);
  assign t[86] = ~(t[110]);
  assign t[87] = ~(t[122]);
  assign t[88] = ~(t[122] & t[90]);
  assign t[89] = ~(t[116]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[119]);
  assign t[91] = t[123] ^ x[2];
  assign t[92] = t[124] ^ x[8];
  assign t[93] = t[125] ^ x[11];
  assign t[94] = t[126] ^ x[14];
  assign t[95] = t[127] ^ x[17];
  assign t[96] = t[128] ^ x[22];
  assign t[97] = t[129] ^ x[25];
  assign t[98] = t[130] ^ x[30];
  assign t[99] = t[131] ^ x[33];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[91];
endmodule

module R1ind181(x, y);
 input [139:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[212] | t[213]);
  assign t[101] = ~(t[137] & t[139]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[142] | t[143]);
  assign t[106] = ~(t[226] | t[144]);
  assign t[107] = t[203] ? x[95] : x[94];
  assign t[108] = ~(t[145] & t[146]);
  assign t[109] = ~(t[227]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[228]);
  assign t[111] = ~(t[147] | t[148]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[229] | t[151]);
  assign t[114] = t[203] ? x[106] : x[105];
  assign t[115] = ~(t[145] & t[152]);
  assign t[116] = ~(t[121] | t[201]);
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = ~(t[202] | t[155]);
  assign t[119] = t[79] & t[201];
  assign t[11] = ~(t[15] ^ t[16]);
  assign t[120] = ~(t[121] | t[156]);
  assign t[121] = ~(t[203]);
  assign t[122] = t[201] ? t[158] : t[157];
  assign t[123] = ~(t[159] & t[204]);
  assign t[124] = ~(t[160] & t[155]);
  assign t[125] = ~(t[230]);
  assign t[126] = ~(t[217] | t[218]);
  assign t[127] = ~(t[161] & t[162]);
  assign t[128] = ~(t[163] & t[78]);
  assign t[129] = ~(t[79] | t[164]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(t[79] | t[165]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[219] | t[220]);
  assign t[133] = ~(t[129] | t[166]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[232]);
  assign t[136] = ~(t[221] | t[222]);
  assign t[137] = ~(t[48] | t[169]);
  assign t[138] = ~(t[170] | t[171]);
  assign t[139] = ~(t[166] | t[130]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = ~(t[233]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[234]);
  assign t[143] = ~(t[235]);
  assign t[144] = ~(t[172] | t[173]);
  assign t[145] = ~(t[48] | t[174]);
  assign t[146] = ~(t[120] | t[175]);
  assign t[147] = ~(t[236]);
  assign t[148] = ~(t[227] | t[228]);
  assign t[149] = ~(t[237]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = ~(t[238]);
  assign t[151] = ~(t[176] | t[177]);
  assign t[152] = ~(t[178] | t[130]);
  assign t[153] = ~(t[204] & t[179]);
  assign t[154] = ~(x[4] & t[118]);
  assign t[155] = ~(t[204]);
  assign t[156] = t[201] ? t[157] : t[158];
  assign t[157] = ~(t[179] & t[155]);
  assign t[158] = ~(x[4] & t[180]);
  assign t[159] = x[4] & t[202];
  assign t[15] = x[4] ? t[24] : t[23];
  assign t[160] = ~(x[4] | t[202]);
  assign t[161] = ~(t[170] | t[181]);
  assign t[162] = ~(t[121] & t[182]);
  assign t[163] = ~(t[183] & t[184]);
  assign t[164] = t[201] ? t[123] : t[124];
  assign t[165] = t[201] ? t[186] : t[185];
  assign t[166] = ~(t[79] | t[187]);
  assign t[167] = t[171] | t[188];
  assign t[168] = ~(t[189] & t[78]);
  assign t[169] = ~(t[79] | t[190]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[121] | t[191]);
  assign t[171] = ~(t[192] & t[76]);
  assign t[172] = ~(t[239]);
  assign t[173] = ~(t[234] | t[235]);
  assign t[174] = ~(t[133] & t[163]);
  assign t[175] = t[169] | t[193];
  assign t[176] = ~(t[240]);
  assign t[177] = ~(t[237] | t[238]);
  assign t[178] = ~(t[79] | t[194]);
  assign t[179] = ~(x[4] | t[195]);
  assign t[17] = t[27] ? x[18] : x[19];
  assign t[180] = ~(t[202] | t[204]);
  assign t[181] = ~(t[79] | t[196]);
  assign t[182] = ~(t[158] & t[153]);
  assign t[183] = t[204] & t[116];
  assign t[184] = t[160] | t[159];
  assign t[185] = ~(t[160] & t[204]);
  assign t[186] = ~(t[159] & t[155]);
  assign t[187] = t[201] ? t[158] : t[153];
  assign t[188] = ~(t[79] | t[197]);
  assign t[189] = ~(t[193] | t[178]);
  assign t[18] = ~(t[28] & t[29]);
  assign t[190] = t[201] ? t[185] : t[186];
  assign t[191] = t[201] ? t[124] : t[186];
  assign t[192] = ~(t[198] | t[120]);
  assign t[193] = ~(t[75]);
  assign t[194] = t[201] ? t[154] : t[157];
  assign t[195] = ~(t[202]);
  assign t[196] = t[201] ? t[157] : t[154];
  assign t[197] = t[201] ? t[153] : t[158];
  assign t[198] = ~(t[121] | t[199]);
  assign t[199] = t[201] ? t[186] : t[124];
  assign t[19] = ~(t[30] | t[31]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[8];
  assign t[202] = t[243] ^ x[11];
  assign t[203] = t[244] ^ x[14];
  assign t[204] = t[245] ^ x[17];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[28];
  assign t[208] = t[249] ^ x[31];
  assign t[209] = t[250] ^ x[34];
  assign t[20] = ~(t[32] ^ t[33]);
  assign t[210] = t[251] ^ x[39];
  assign t[211] = t[252] ^ x[42];
  assign t[212] = t[253] ^ x[45];
  assign t[213] = t[254] ^ x[48];
  assign t[214] = t[255] ^ x[53];
  assign t[215] = t[256] ^ x[56];
  assign t[216] = t[257] ^ x[59];
  assign t[217] = t[258] ^ x[62];
  assign t[218] = t[259] ^ x[65];
  assign t[219] = t[260] ^ x[68];
  assign t[21] = x[4] ? t[35] : t[34];
  assign t[220] = t[261] ^ x[71];
  assign t[221] = t[262] ^ x[76];
  assign t[222] = t[263] ^ x[79];
  assign t[223] = t[264] ^ x[84];
  assign t[224] = t[265] ^ x[87];
  assign t[225] = t[266] ^ x[90];
  assign t[226] = t[267] ^ x[93];
  assign t[227] = t[268] ^ x[98];
  assign t[228] = t[269] ^ x[101];
  assign t[229] = t[270] ^ x[104];
  assign t[22] = x[4] ? t[37] : t[36];
  assign t[230] = t[271] ^ x[109];
  assign t[231] = t[272] ^ x[112];
  assign t[232] = t[273] ^ x[115];
  assign t[233] = t[274] ^ x[118];
  assign t[234] = t[275] ^ x[121];
  assign t[235] = t[276] ^ x[124];
  assign t[236] = t[277] ^ x[127];
  assign t[237] = t[278] ^ x[130];
  assign t[238] = t[279] ^ x[133];
  assign t[239] = t[280] ^ x[136];
  assign t[23] = ~(t[38] | t[39]);
  assign t[240] = t[281] ^ x[139];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[6] & x[7]);
  assign t[243] = (x[9] & x[10]);
  assign t[244] = (x[12] & x[13]);
  assign t[245] = (x[15] & x[16]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[26] & x[27]);
  assign t[249] = (x[29] & x[30]);
  assign t[24] = ~(t[23] ^ t[40]);
  assign t[250] = (x[32] & x[33]);
  assign t[251] = (x[37] & x[38]);
  assign t[252] = (x[40] & x[41]);
  assign t[253] = (x[43] & x[44]);
  assign t[254] = (x[46] & x[47]);
  assign t[255] = (x[51] & x[52]);
  assign t[256] = (x[54] & x[55]);
  assign t[257] = (x[57] & x[58]);
  assign t[258] = (x[60] & x[61]);
  assign t[259] = (x[63] & x[64]);
  assign t[25] = x[4] ? t[42] : t[41];
  assign t[260] = (x[66] & x[67]);
  assign t[261] = (x[69] & x[70]);
  assign t[262] = (x[74] & x[75]);
  assign t[263] = (x[77] & x[78]);
  assign t[264] = (x[82] & x[83]);
  assign t[265] = (x[85] & x[86]);
  assign t[266] = (x[88] & x[89]);
  assign t[267] = (x[91] & x[92]);
  assign t[268] = (x[96] & x[97]);
  assign t[269] = (x[99] & x[100]);
  assign t[26] = x[4] ? t[44] : t[43];
  assign t[270] = (x[102] & x[103]);
  assign t[271] = (x[107] & x[108]);
  assign t[272] = (x[110] & x[111]);
  assign t[273] = (x[113] & x[114]);
  assign t[274] = (x[116] & x[117]);
  assign t[275] = (x[119] & x[120]);
  assign t[276] = (x[122] & x[123]);
  assign t[277] = (x[125] & x[126]);
  assign t[278] = (x[128] & x[129]);
  assign t[279] = (x[131] & x[132]);
  assign t[27] = ~(t[45]);
  assign t[280] = (x[134] & x[135]);
  assign t[281] = (x[137] & x[138]);
  assign t[28] = ~(t[46] | t[47]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[205] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[54] ^ t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[43] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[34] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[206] | t[64]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[45] = ~(t[203]);
  assign t[46] = ~(t[75] & t[76]);
  assign t[47] = ~(t[77] & t[78]);
  assign t[48] = ~(t[79] | t[80]);
  assign t[49] = ~(t[207]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[208]);
  assign t[51] = ~(t[81] | t[82]);
  assign t[52] = ~(t[83] | t[84]);
  assign t[53] = ~(t[209] | t[85]);
  assign t[54] = t[86] ? x[36] : x[35];
  assign t[55] = ~(t[87] & t[88]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[210] | t[91]);
  assign t[58] = ~(t[92] ^ t[93]);
  assign t[59] = ~(t[94] | t[95]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[211] | t[96]);
  assign t[61] = ~(t[97] ^ t[98]);
  assign t[62] = ~(t[212]);
  assign t[63] = ~(t[213]);
  assign t[64] = ~(t[99] | t[100]);
  assign t[65] = t[203] ? x[50] : x[49];
  assign t[66] = t[46] | t[101];
  assign t[67] = ~(t[102] | t[103]);
  assign t[68] = ~(t[214] | t[104]);
  assign t[69] = ~(t[105] | t[106]);
  assign t[6] = ~(t[201] & t[202]);
  assign t[70] = ~(t[107] ^ t[108]);
  assign t[71] = ~(t[109] | t[110]);
  assign t[72] = ~(t[215] | t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[114] ^ t[115]);
  assign t[75] = ~(t[116] & t[117]);
  assign t[76] = ~(t[118] & t[119]);
  assign t[77] = ~(t[120]);
  assign t[78] = t[121] | t[122];
  assign t[79] = ~(t[121]);
  assign t[7] = ~(t[203] & t[204]);
  assign t[80] = t[201] ? t[124] : t[123];
  assign t[81] = ~(t[216]);
  assign t[82] = ~(t[207] | t[208]);
  assign t[83] = ~(t[217]);
  assign t[84] = ~(t[218]);
  assign t[85] = ~(t[125] | t[126]);
  assign t[86] = ~(t[45]);
  assign t[87] = ~(t[127] | t[128]);
  assign t[88] = ~(t[129] | t[130]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[11] ^ t[12]);
  assign t[90] = ~(t[220]);
  assign t[91] = ~(t[131] | t[132]);
  assign t[92] = t[86] ? x[73] : x[72];
  assign t[93] = ~(t[133] & t[134]);
  assign t[94] = ~(t[221]);
  assign t[95] = ~(t[222]);
  assign t[96] = ~(t[135] | t[136]);
  assign t[97] = t[86] ? x[81] : x[80];
  assign t[98] = ~(t[137] & t[138]);
  assign t[99] = ~(t[223]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind182(x, y);
 input [97:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = (x[20] & x[21]);
  assign t[101] = (x[25] & x[26]);
  assign t[102] = (x[28] & x[29]);
  assign t[103] = (x[31] & x[32]);
  assign t[104] = (x[34] & x[35]);
  assign t[105] = (x[39] & x[40]);
  assign t[106] = (x[44] & x[45]);
  assign t[107] = (x[47] & x[48]);
  assign t[108] = (x[50] & x[51]);
  assign t[109] = (x[53] & x[54]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = (x[56] & x[57]);
  assign t[111] = (x[59] & x[60]);
  assign t[112] = (x[62] & x[63]);
  assign t[113] = (x[65] & x[66]);
  assign t[114] = (x[68] & x[69]);
  assign t[115] = (x[71] & x[72]);
  assign t[116] = (x[74] & x[75]);
  assign t[117] = (x[77] & x[78]);
  assign t[118] = (x[80] & x[81]);
  assign t[119] = (x[83] & x[84]);
  assign t[11] = t[69] ? x[18] : x[19];
  assign t[120] = (x[86] & x[87]);
  assign t[121] = (x[89] & x[90]);
  assign t[122] = (x[92] & x[93]);
  assign t[123] = (x[95] & x[96]);
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[71];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[69] ? x[24] : x[23];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = t[33] ^ t[34];
  assign t[24] = ~(t[35] & t[36]);
  assign t[25] = t[37] ^ t[38];
  assign t[26] = ~(t[72]);
  assign t[27] = ~(t[73]);
  assign t[28] = ~(t[39] | t[26]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[42] | t[74];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] | t[75];
  assign t[33] = t[69] ? x[38] : x[37];
  assign t[34] = ~(t[46] & t[47]);
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = t[50] | t[76];
  assign t[37] = t[51] ? x[43] : x[42];
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[77]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[78]);
  assign t[41] = ~(t[79]);
  assign t[42] = ~(t[54] | t[40]);
  assign t[43] = ~(t[80]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[55] | t[43]);
  assign t[46] = ~(t[56] & t[57]);
  assign t[47] = t[58] | t[82];
  assign t[48] = ~(t[83]);
  assign t[49] = ~(t[84]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[59] | t[48]);
  assign t[51] = ~(t[60]);
  assign t[52] = ~(t[61] & t[62]);
  assign t[53] = t[63] | t[85];
  assign t[54] = ~(t[86]);
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[89]);
  assign t[58] = ~(t[64] | t[56]);
  assign t[59] = ~(t[90]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[69]);
  assign t[61] = ~(t[91]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[65] | t[61]);
  assign t[64] = ~(t[93]);
  assign t[65] = ~(t[94]);
  assign t[66] = t[95] ^ x[2];
  assign t[67] = t[96] ^ x[8];
  assign t[68] = t[97] ^ x[11];
  assign t[69] = t[98] ^ x[14];
  assign t[6] = ~(t[67] & t[68]);
  assign t[70] = t[99] ^ x[17];
  assign t[71] = t[100] ^ x[22];
  assign t[72] = t[101] ^ x[27];
  assign t[73] = t[102] ^ x[30];
  assign t[74] = t[103] ^ x[33];
  assign t[75] = t[104] ^ x[36];
  assign t[76] = t[105] ^ x[41];
  assign t[77] = t[106] ^ x[46];
  assign t[78] = t[107] ^ x[49];
  assign t[79] = t[108] ^ x[52];
  assign t[7] = ~(t[69] & t[70]);
  assign t[80] = t[109] ^ x[55];
  assign t[81] = t[110] ^ x[58];
  assign t[82] = t[111] ^ x[61];
  assign t[83] = t[112] ^ x[64];
  assign t[84] = t[113] ^ x[67];
  assign t[85] = t[114] ^ x[70];
  assign t[86] = t[115] ^ x[73];
  assign t[87] = t[116] ^ x[76];
  assign t[88] = t[117] ^ x[79];
  assign t[89] = t[118] ^ x[82];
  assign t[8] = t[11] ^ t[9];
  assign t[90] = t[119] ^ x[85];
  assign t[91] = t[120] ^ x[88];
  assign t[92] = t[121] ^ x[91];
  assign t[93] = t[122] ^ x[94];
  assign t[94] = t[123] ^ x[97];
  assign t[95] = (x[0] & x[1]);
  assign t[96] = (x[6] & x[7]);
  assign t[97] = (x[9] & x[10]);
  assign t[98] = (x[12] & x[13]);
  assign t[99] = (x[15] & x[16]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[66];
endmodule

module R1ind183(x, y);
 input [97:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[129] ^ x[97];
  assign t[101] = (x[0] & x[1]);
  assign t[102] = (x[6] & x[7]);
  assign t[103] = (x[9] & x[10]);
  assign t[104] = (x[12] & x[13]);
  assign t[105] = (x[15] & x[16]);
  assign t[106] = (x[20] & x[21]);
  assign t[107] = (x[25] & x[26]);
  assign t[108] = (x[28] & x[29]);
  assign t[109] = (x[31] & x[32]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = (x[34] & x[35]);
  assign t[111] = (x[39] & x[40]);
  assign t[112] = (x[44] & x[45]);
  assign t[113] = (x[47] & x[48]);
  assign t[114] = (x[50] & x[51]);
  assign t[115] = (x[53] & x[54]);
  assign t[116] = (x[56] & x[57]);
  assign t[117] = (x[59] & x[60]);
  assign t[118] = (x[62] & x[63]);
  assign t[119] = (x[65] & x[66]);
  assign t[11] = t[75] ? x[18] : x[19];
  assign t[120] = (x[68] & x[69]);
  assign t[121] = (x[71] & x[72]);
  assign t[122] = (x[74] & x[75]);
  assign t[123] = (x[77] & x[78]);
  assign t[124] = (x[80] & x[81]);
  assign t[125] = (x[83] & x[84]);
  assign t[126] = (x[86] & x[87]);
  assign t[127] = (x[89] & x[90]);
  assign t[128] = (x[92] & x[93]);
  assign t[129] = (x[95] & x[96]);
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[77]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[75] ? x[24] : x[23];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = t[33] ^ t[34];
  assign t[24] = ~(t[35] & t[36]);
  assign t[25] = t[37] ^ t[38];
  assign t[26] = ~(t[78]);
  assign t[27] = ~(t[79]);
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = ~(t[41] & t[42]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[43] & t[80]);
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[46] & t[81]);
  assign t[33] = t[75] ? x[38] : x[37];
  assign t[34] = ~(t[47] & t[48]);
  assign t[35] = ~(t[49] & t[50]);
  assign t[36] = ~(t[51] & t[82]);
  assign t[37] = t[52] ? x[43] : x[42];
  assign t[38] = ~(t[53] & t[54]);
  assign t[39] = ~(t[79] & t[78]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[83]);
  assign t[41] = ~(t[84]);
  assign t[42] = ~(t[85]);
  assign t[43] = ~(t[55] & t[56]);
  assign t[44] = ~(t[86]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[57] & t[58]);
  assign t[47] = ~(t[59] & t[60]);
  assign t[48] = ~(t[61] & t[88]);
  assign t[49] = ~(t[89]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[90]);
  assign t[51] = ~(t[62] & t[63]);
  assign t[52] = ~(t[64]);
  assign t[53] = ~(t[65] & t[66]);
  assign t[54] = ~(t[67] & t[91]);
  assign t[55] = ~(t[85] & t[84]);
  assign t[56] = ~(t[92]);
  assign t[57] = ~(t[87] & t[86]);
  assign t[58] = ~(t[93]);
  assign t[59] = ~(t[94]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[68] & t[69]);
  assign t[62] = ~(t[90] & t[89]);
  assign t[63] = ~(t[96]);
  assign t[64] = ~(t[75]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[70] & t[71]);
  assign t[68] = ~(t[95] & t[94]);
  assign t[69] = ~(t[99]);
  assign t[6] = ~(t[73] & t[74]);
  assign t[70] = ~(t[98] & t[97]);
  assign t[71] = ~(t[100]);
  assign t[72] = t[101] ^ x[2];
  assign t[73] = t[102] ^ x[8];
  assign t[74] = t[103] ^ x[11];
  assign t[75] = t[104] ^ x[14];
  assign t[76] = t[105] ^ x[17];
  assign t[77] = t[106] ^ x[22];
  assign t[78] = t[107] ^ x[27];
  assign t[79] = t[108] ^ x[30];
  assign t[7] = ~(t[75] & t[76]);
  assign t[80] = t[109] ^ x[33];
  assign t[81] = t[110] ^ x[36];
  assign t[82] = t[111] ^ x[41];
  assign t[83] = t[112] ^ x[46];
  assign t[84] = t[113] ^ x[49];
  assign t[85] = t[114] ^ x[52];
  assign t[86] = t[115] ^ x[55];
  assign t[87] = t[116] ^ x[58];
  assign t[88] = t[117] ^ x[61];
  assign t[89] = t[118] ^ x[64];
  assign t[8] = t[11] ^ t[9];
  assign t[90] = t[119] ^ x[67];
  assign t[91] = t[120] ^ x[70];
  assign t[92] = t[121] ^ x[73];
  assign t[93] = t[122] ^ x[76];
  assign t[94] = t[123] ^ x[79];
  assign t[95] = t[124] ^ x[82];
  assign t[96] = t[125] ^ x[85];
  assign t[97] = t[126] ^ x[88];
  assign t[98] = t[127] ^ x[91];
  assign t[99] = t[128] ^ x[94];
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[72];
endmodule

module R1ind184(x, y);
 input [79:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = (x[62] & x[63]);
  assign t[101] = (x[65] & x[66]);
  assign t[102] = (x[68] & x[69]);
  assign t[103] = (x[71] & x[72]);
  assign t[104] = (x[74] & x[75]);
  assign t[105] = (x[77] & x[78]);
  assign t[10] = x[18] ^ x[19];
  assign t[11] = t[63] ? x[19] : x[18];
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[65] & t[26]);
  assign t[19] = ~(t[66] & t[27]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[63] ? x[27] : x[26];
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] ^ t[33];
  assign t[24] = ~(t[34] & t[35]);
  assign t[25] = t[36] ^ t[37];
  assign t[26] = ~(t[67]);
  assign t[27] = ~(t[67] & t[38]);
  assign t[28] = ~(t[68] & t[39]);
  assign t[29] = ~(t[69] & t[40]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[70] & t[41]);
  assign t[31] = ~(t[71] & t[42]);
  assign t[32] = t[63] ? x[44] : x[43];
  assign t[33] = ~(t[43] & t[44]);
  assign t[34] = ~(t[72] & t[45]);
  assign t[35] = ~(t[73] & t[46]);
  assign t[36] = t[47] ? x[52] : x[51];
  assign t[37] = ~(t[48] & t[49]);
  assign t[38] = ~(t[65]);
  assign t[39] = ~(t[74]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[74] & t[50]);
  assign t[41] = ~(t[75]);
  assign t[42] = ~(t[75] & t[51]);
  assign t[43] = ~(t[76] & t[52]);
  assign t[44] = ~(t[77] & t[53]);
  assign t[45] = ~(t[78]);
  assign t[46] = ~(t[78] & t[54]);
  assign t[47] = ~(t[55]);
  assign t[48] = ~(t[79] & t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[68]);
  assign t[51] = ~(t[70]);
  assign t[52] = ~(t[81]);
  assign t[53] = ~(t[81] & t[58]);
  assign t[54] = ~(t[72]);
  assign t[55] = ~(t[63]);
  assign t[56] = ~(t[82]);
  assign t[57] = ~(t[82] & t[59]);
  assign t[58] = ~(t[76]);
  assign t[59] = ~(t[79]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = t[83] ^ x[2];
  assign t[61] = t[84] ^ x[8];
  assign t[62] = t[85] ^ x[11];
  assign t[63] = t[86] ^ x[14];
  assign t[64] = t[87] ^ x[17];
  assign t[65] = t[88] ^ x[22];
  assign t[66] = t[89] ^ x[25];
  assign t[67] = t[90] ^ x[30];
  assign t[68] = t[91] ^ x[33];
  assign t[69] = t[92] ^ x[36];
  assign t[6] = ~(t[61] & t[62]);
  assign t[70] = t[93] ^ x[39];
  assign t[71] = t[94] ^ x[42];
  assign t[72] = t[95] ^ x[47];
  assign t[73] = t[96] ^ x[50];
  assign t[74] = t[97] ^ x[55];
  assign t[75] = t[98] ^ x[58];
  assign t[76] = t[99] ^ x[61];
  assign t[77] = t[100] ^ x[64];
  assign t[78] = t[101] ^ x[67];
  assign t[79] = t[102] ^ x[70];
  assign t[7] = ~(t[63] & t[64]);
  assign t[80] = t[103] ^ x[73];
  assign t[81] = t[104] ^ x[76];
  assign t[82] = t[105] ^ x[79];
  assign t[83] = (x[0] & x[1]);
  assign t[84] = (x[6] & x[7]);
  assign t[85] = (x[9] & x[10]);
  assign t[86] = (x[12] & x[13]);
  assign t[87] = (x[15] & x[16]);
  assign t[88] = (x[20] & x[21]);
  assign t[89] = (x[23] & x[24]);
  assign t[8] = t[11] ^ t[9];
  assign t[90] = (x[28] & x[29]);
  assign t[91] = (x[31] & x[32]);
  assign t[92] = (x[34] & x[35]);
  assign t[93] = (x[37] & x[38]);
  assign t[94] = (x[40] & x[41]);
  assign t[95] = (x[45] & x[46]);
  assign t[96] = (x[48] & x[49]);
  assign t[97] = (x[53] & x[54]);
  assign t[98] = (x[56] & x[57]);
  assign t[99] = (x[59] & x[60]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[60];
endmodule

module R1ind185(x, y);
 input [97:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[153] | t[154]);
  assign t[101] = ~(t[161]);
  assign t[102] = ~(t[162]);
  assign t[103] = ~(t[118] | t[119]);
  assign t[104] = ~(t[120] | t[56]);
  assign t[105] = ~(x[4] | t[121]);
  assign t[106] = ~(t[122] & t[140]);
  assign t[107] = ~(t[123] & t[82]);
  assign t[108] = ~(t[122] & t[82]);
  assign t[109] = ~(t[123] & t[140]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(x[4] & t[124]);
  assign t[111] = ~(t[116]);
  assign t[112] = t[79] | t[125];
  assign t[113] = ~(t[163]);
  assign t[114] = ~(t[158] | t[159]);
  assign t[115] = ~(t[126] & t[127]);
  assign t[116] = ~(t[79] | t[128]);
  assign t[117] = t[54] | t[129];
  assign t[118] = ~(t[164]);
  assign t[119] = ~(t[161] | t[162]);
  assign t[11] = ~(t[14] ^ t[15]);
  assign t[120] = ~(t[83] | t[130]);
  assign t[121] = ~(t[138]);
  assign t[122] = x[4] & t[138];
  assign t[123] = ~(x[4] | t[138]);
  assign t[124] = ~(t[138] | t[140]);
  assign t[125] = t[137] ? t[110] : t[131];
  assign t[126] = ~(t[132] | t[55]);
  assign t[127] = ~(t[133] & t[134]);
  assign t[128] = t[137] ? t[131] : t[110];
  assign t[129] = ~(t[30]);
  assign t[12] = x[4] ? t[17] : t[16];
  assign t[130] = t[137] ? t[81] : t[131];
  assign t[131] = ~(t[105] & t[82]);
  assign t[132] = ~(t[83] | t[135]);
  assign t[133] = t[140] & t[49];
  assign t[134] = t[123] | t[122];
  assign t[135] = t[137] ? t[106] : t[107];
  assign t[136] = t[165] ^ x[2];
  assign t[137] = t[166] ^ x[8];
  assign t[138] = t[167] ^ x[11];
  assign t[139] = t[168] ^ x[14];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[169] ^ x[17];
  assign t[141] = t[170] ^ x[22];
  assign t[142] = t[171] ^ x[25];
  assign t[143] = t[172] ^ x[28];
  assign t[144] = t[173] ^ x[31];
  assign t[145] = t[174] ^ x[36];
  assign t[146] = t[175] ^ x[39];
  assign t[147] = t[176] ^ x[42];
  assign t[148] = t[177] ^ x[45];
  assign t[149] = t[178] ^ x[48];
  assign t[14] = t[139] ? x[19] : x[18];
  assign t[150] = t[179] ^ x[51];
  assign t[151] = t[180] ^ x[54];
  assign t[152] = t[181] ^ x[57];
  assign t[153] = t[182] ^ x[62];
  assign t[154] = t[183] ^ x[65];
  assign t[155] = t[184] ^ x[68];
  assign t[156] = t[185] ^ x[73];
  assign t[157] = t[186] ^ x[76];
  assign t[158] = t[187] ^ x[79];
  assign t[159] = t[188] ^ x[82];
  assign t[15] = t[20] | t[21];
  assign t[160] = t[189] ^ x[85];
  assign t[161] = t[190] ^ x[88];
  assign t[162] = t[191] ^ x[91];
  assign t[163] = t[192] ^ x[94];
  assign t[164] = t[193] ^ x[97];
  assign t[165] = (x[0] & x[1]);
  assign t[166] = (x[6] & x[7]);
  assign t[167] = (x[9] & x[10]);
  assign t[168] = (x[12] & x[13]);
  assign t[169] = (x[15] & x[16]);
  assign t[16] = ~(t[22] | t[23]);
  assign t[170] = (x[20] & x[21]);
  assign t[171] = (x[23] & x[24]);
  assign t[172] = (x[26] & x[27]);
  assign t[173] = (x[29] & x[30]);
  assign t[174] = (x[34] & x[35]);
  assign t[175] = (x[37] & x[38]);
  assign t[176] = (x[40] & x[41]);
  assign t[177] = (x[43] & x[44]);
  assign t[178] = (x[46] & x[47]);
  assign t[179] = (x[49] & x[50]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (x[52] & x[53]);
  assign t[181] = (x[55] & x[56]);
  assign t[182] = (x[60] & x[61]);
  assign t[183] = (x[63] & x[64]);
  assign t[184] = (x[66] & x[67]);
  assign t[185] = (x[71] & x[72]);
  assign t[186] = (x[74] & x[75]);
  assign t[187] = (x[77] & x[78]);
  assign t[188] = (x[80] & x[81]);
  assign t[189] = (x[83] & x[84]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = (x[86] & x[87]);
  assign t[191] = (x[89] & x[90]);
  assign t[192] = (x[92] & x[93]);
  assign t[193] = (x[95] & x[96]);
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = ~(t[30] & t[31]);
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[141] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[28] = ~(t[45] | t[46]);
  assign t[29] = ~(t[47] ^ t[48]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[49] & t[50]);
  assign t[31] = ~(t[51] & t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[55] | t[56]);
  assign t[34] = ~(t[142]);
  assign t[35] = ~(t[143]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[59] | t[60]);
  assign t[38] = ~(t[144] | t[61]);
  assign t[39] = t[62] ? x[33] : x[32];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[63] & t[64]);
  assign t[41] = ~(t[65] | t[66]);
  assign t[42] = ~(t[145] | t[67]);
  assign t[43] = ~(t[68] | t[69]);
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = ~(t[72] | t[73]);
  assign t[46] = ~(t[146] | t[74]);
  assign t[47] = ~(t[75] | t[76]);
  assign t[48] = ~(t[77] ^ t[78]);
  assign t[49] = ~(t[79] | t[137]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[80] & t[81]);
  assign t[51] = ~(t[138] | t[82]);
  assign t[52] = t[83] & t[137];
  assign t[53] = ~(t[83] | t[84]);
  assign t[54] = ~(t[83] | t[85]);
  assign t[55] = ~(t[83] | t[86]);
  assign t[56] = ~(t[83] | t[87]);
  assign t[57] = ~(t[147]);
  assign t[58] = ~(t[142] | t[143]);
  assign t[59] = ~(t[148]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[149]);
  assign t[61] = ~(t[88] | t[89]);
  assign t[62] = ~(t[90]);
  assign t[63] = ~(t[20] | t[91]);
  assign t[64] = ~(t[53]);
  assign t[65] = ~(t[150]);
  assign t[66] = ~(t[151]);
  assign t[67] = ~(t[92] | t[93]);
  assign t[68] = ~(t[94] | t[95]);
  assign t[69] = ~(t[152] | t[96]);
  assign t[6] = ~(t[137] & t[138]);
  assign t[70] = t[139] ? x[59] : x[58];
  assign t[71] = ~(t[97] & t[98]);
  assign t[72] = ~(t[153]);
  assign t[73] = ~(t[154]);
  assign t[74] = ~(t[99] | t[100]);
  assign t[75] = ~(t[101] | t[102]);
  assign t[76] = ~(t[155] | t[103]);
  assign t[77] = t[139] ? x[70] : x[69];
  assign t[78] = ~(t[97] & t[104]);
  assign t[79] = ~(t[139]);
  assign t[7] = ~(t[139] & t[140]);
  assign t[80] = ~(t[140] & t[105]);
  assign t[81] = ~(x[4] & t[51]);
  assign t[82] = ~(t[140]);
  assign t[83] = ~(t[79]);
  assign t[84] = t[137] ? t[107] : t[106];
  assign t[85] = t[137] ? t[109] : t[108];
  assign t[86] = t[137] ? t[110] : t[80];
  assign t[87] = t[137] ? t[108] : t[109];
  assign t[88] = ~(t[156]);
  assign t[89] = ~(t[148] | t[149]);
  assign t[8] = ~(t[9] ^ t[11]);
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[111] & t[112]);
  assign t[92] = ~(t[157]);
  assign t[93] = ~(t[150] | t[151]);
  assign t[94] = ~(t[158]);
  assign t[95] = ~(t[159]);
  assign t[96] = ~(t[113] | t[114]);
  assign t[97] = ~(t[53] | t[115]);
  assign t[98] = ~(t[116] | t[117]);
  assign t[99] = ~(t[160]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[136];
endmodule

module R1ind186(x, y);
 input [151:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[105] | t[100]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[150]);
  assign t[106] = t[151] ^ x[2];
  assign t[107] = t[152] ^ x[8];
  assign t[108] = t[153] ^ x[11];
  assign t[109] = t[154] ^ x[14];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[155] ^ x[17];
  assign t[111] = t[156] ^ x[22];
  assign t[112] = t[157] ^ x[27];
  assign t[113] = t[158] ^ x[32];
  assign t[114] = t[159] ^ x[35];
  assign t[115] = t[160] ^ x[38];
  assign t[116] = t[161] ^ x[41];
  assign t[117] = t[162] ^ x[46];
  assign t[118] = t[163] ^ x[51];
  assign t[119] = t[164] ^ x[54];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[165] ^ x[57];
  assign t[121] = t[166] ^ x[60];
  assign t[122] = t[167] ^ x[65];
  assign t[123] = t[168] ^ x[70];
  assign t[124] = t[169] ^ x[73];
  assign t[125] = t[170] ^ x[76];
  assign t[126] = t[171] ^ x[79];
  assign t[127] = t[172] ^ x[82];
  assign t[128] = t[173] ^ x[85];
  assign t[129] = t[174] ^ x[88];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[91];
  assign t[131] = t[176] ^ x[94];
  assign t[132] = t[177] ^ x[97];
  assign t[133] = t[178] ^ x[100];
  assign t[134] = t[179] ^ x[103];
  assign t[135] = t[180] ^ x[106];
  assign t[136] = t[181] ^ x[109];
  assign t[137] = t[182] ^ x[112];
  assign t[138] = t[183] ^ x[115];
  assign t[139] = t[184] ^ x[118];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[121];
  assign t[141] = t[186] ^ x[124];
  assign t[142] = t[187] ^ x[127];
  assign t[143] = t[188] ^ x[130];
  assign t[144] = t[189] ^ x[133];
  assign t[145] = t[190] ^ x[136];
  assign t[146] = t[191] ^ x[139];
  assign t[147] = t[192] ^ x[142];
  assign t[148] = t[193] ^ x[145];
  assign t[149] = t[194] ^ x[148];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[151];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[6] & x[7]);
  assign t[153] = (x[9] & x[10]);
  assign t[154] = (x[12] & x[13]);
  assign t[155] = (x[15] & x[16]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[30] & x[31]);
  assign t[159] = (x[33] & x[34]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[36] & x[37]);
  assign t[161] = (x[39] & x[40]);
  assign t[162] = (x[44] & x[45]);
  assign t[163] = (x[49] & x[50]);
  assign t[164] = (x[52] & x[53]);
  assign t[165] = (x[55] & x[56]);
  assign t[166] = (x[58] & x[59]);
  assign t[167] = (x[63] & x[64]);
  assign t[168] = (x[68] & x[69]);
  assign t[169] = (x[71] & x[72]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[74] & x[75]);
  assign t[171] = (x[77] & x[78]);
  assign t[172] = (x[80] & x[81]);
  assign t[173] = (x[83] & x[84]);
  assign t[174] = (x[86] & x[87]);
  assign t[175] = (x[89] & x[90]);
  assign t[176] = (x[92] & x[93]);
  assign t[177] = (x[95] & x[96]);
  assign t[178] = (x[98] & x[99]);
  assign t[179] = (x[101] & x[102]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[104] & x[105]);
  assign t[181] = (x[107] & x[108]);
  assign t[182] = (x[110] & x[111]);
  assign t[183] = (x[113] & x[114]);
  assign t[184] = (x[116] & x[117]);
  assign t[185] = (x[119] & x[120]);
  assign t[186] = (x[122] & x[123]);
  assign t[187] = (x[125] & x[126]);
  assign t[188] = (x[128] & x[129]);
  assign t[189] = (x[131] & x[132]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[134] & x[135]);
  assign t[191] = (x[137] & x[138]);
  assign t[192] = (x[140] & x[141]);
  assign t[193] = (x[143] & x[144]);
  assign t[194] = (x[146] & x[147]);
  assign t[195] = (x[149] & x[150]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[109]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = t[45] | t[111];
  assign t[29] = t[15] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[39];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] | t[112];
  assign t[37] = t[109] ? x[29] : x[28];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[113]);
  assign t[44] = ~(t[114]);
  assign t[45] = ~(t[67] | t[43]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = t[70] | t[115];
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = t[73] | t[116];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[74] ? x[43] : x[42];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[117];
  assign t[53] = t[74] ? x[48] : x[47];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[118]);
  assign t[56] = ~(t[119]);
  assign t[57] = ~(t[80] | t[55]);
  assign t[58] = ~(t[81] & t[82]);
  assign t[59] = t[83] | t[120];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = t[86] | t[121];
  assign t[62] = t[109] ? x[62] : x[61];
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = t[91] | t[122];
  assign t[66] = t[109] ? x[67] : x[66];
  assign t[67] = ~(t[123]);
  assign t[68] = ~(t[124]);
  assign t[69] = ~(t[125]);
  assign t[6] = ~(t[107] & t[108]);
  assign t[70] = ~(t[92] | t[68]);
  assign t[71] = ~(t[126]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[93] | t[71]);
  assign t[74] = ~(t[22]);
  assign t[75] = ~(t[128]);
  assign t[76] = ~(t[129]);
  assign t[77] = ~(t[94] | t[75]);
  assign t[78] = ~(t[95] & t[96]);
  assign t[79] = t[97] | t[130];
  assign t[7] = ~(t[109] & t[110]);
  assign t[80] = ~(t[131]);
  assign t[81] = ~(t[132]);
  assign t[82] = ~(t[133]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[134]);
  assign t[85] = ~(t[135]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[100] & t[101]);
  assign t[88] = t[102] | t[136];
  assign t[89] = ~(t[137]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[103] | t[89]);
  assign t[92] = ~(t[139]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[141]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[104] | t[95]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[106];
endmodule

module R1ind187(x, y);
 input [151:0] x;
 output y;

 wire [205:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[112] & t[113]);
  assign t[103] = ~(t[143] & t[142]);
  assign t[104] = ~(t[154]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[155]);
  assign t[107] = ~(t[156]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[114] & t[115]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[148] & t[147]);
  assign t[111] = ~(t[158]);
  assign t[112] = ~(t[153] & t[152]);
  assign t[113] = ~(t[159]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[160]);
  assign t[116] = t[161] ^ x[2];
  assign t[117] = t[162] ^ x[8];
  assign t[118] = t[163] ^ x[11];
  assign t[119] = t[164] ^ x[14];
  assign t[11] = t[15] ? x[18] : x[19];
  assign t[120] = t[165] ^ x[17];
  assign t[121] = t[166] ^ x[22];
  assign t[122] = t[167] ^ x[27];
  assign t[123] = t[168] ^ x[32];
  assign t[124] = t[169] ^ x[35];
  assign t[125] = t[170] ^ x[38];
  assign t[126] = t[171] ^ x[41];
  assign t[127] = t[172] ^ x[46];
  assign t[128] = t[173] ^ x[51];
  assign t[129] = t[174] ^ x[54];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[57];
  assign t[131] = t[176] ^ x[60];
  assign t[132] = t[177] ^ x[65];
  assign t[133] = t[178] ^ x[70];
  assign t[134] = t[179] ^ x[73];
  assign t[135] = t[180] ^ x[76];
  assign t[136] = t[181] ^ x[79];
  assign t[137] = t[182] ^ x[82];
  assign t[138] = t[183] ^ x[85];
  assign t[139] = t[184] ^ x[88];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[91];
  assign t[141] = t[186] ^ x[94];
  assign t[142] = t[187] ^ x[97];
  assign t[143] = t[188] ^ x[100];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[106];
  assign t[146] = t[191] ^ x[109];
  assign t[147] = t[192] ^ x[112];
  assign t[148] = t[193] ^ x[115];
  assign t[149] = t[194] ^ x[118];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[121];
  assign t[151] = t[196] ^ x[124];
  assign t[152] = t[197] ^ x[127];
  assign t[153] = t[198] ^ x[130];
  assign t[154] = t[199] ^ x[133];
  assign t[155] = t[200] ^ x[136];
  assign t[156] = t[201] ^ x[139];
  assign t[157] = t[202] ^ x[142];
  assign t[158] = t[203] ^ x[145];
  assign t[159] = t[204] ^ x[148];
  assign t[15] = ~(t[22]);
  assign t[160] = t[205] ^ x[151];
  assign t[161] = (x[0] & x[1]);
  assign t[162] = (x[6] & x[7]);
  assign t[163] = (x[9] & x[10]);
  assign t[164] = (x[12] & x[13]);
  assign t[165] = (x[15] & x[16]);
  assign t[166] = (x[20] & x[21]);
  assign t[167] = (x[25] & x[26]);
  assign t[168] = (x[30] & x[31]);
  assign t[169] = (x[33] & x[34]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[36] & x[37]);
  assign t[171] = (x[39] & x[40]);
  assign t[172] = (x[44] & x[45]);
  assign t[173] = (x[49] & x[50]);
  assign t[174] = (x[52] & x[53]);
  assign t[175] = (x[55] & x[56]);
  assign t[176] = (x[58] & x[59]);
  assign t[177] = (x[63] & x[64]);
  assign t[178] = (x[68] & x[69]);
  assign t[179] = (x[71] & x[72]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[74] & x[75]);
  assign t[181] = (x[77] & x[78]);
  assign t[182] = (x[80] & x[81]);
  assign t[183] = (x[83] & x[84]);
  assign t[184] = (x[86] & x[87]);
  assign t[185] = (x[89] & x[90]);
  assign t[186] = (x[92] & x[93]);
  assign t[187] = (x[95] & x[96]);
  assign t[188] = (x[98] & x[99]);
  assign t[189] = (x[101] & x[102]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[104] & x[105]);
  assign t[191] = (x[107] & x[108]);
  assign t[192] = (x[110] & x[111]);
  assign t[193] = (x[113] & x[114]);
  assign t[194] = (x[116] & x[117]);
  assign t[195] = (x[119] & x[120]);
  assign t[196] = (x[122] & x[123]);
  assign t[197] = (x[125] & x[126]);
  assign t[198] = (x[128] & x[129]);
  assign t[199] = (x[131] & x[132]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = (x[134] & x[135]);
  assign t[201] = (x[137] & x[138]);
  assign t[202] = (x[140] & x[141]);
  assign t[203] = (x[143] & x[144]);
  assign t[204] = (x[146] & x[147]);
  assign t[205] = (x[149] & x[150]);
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[119]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = ~(t[45] & t[121]);
  assign t[29] = t[46] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[39];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = ~(t[56] & t[57]);
  assign t[36] = ~(t[58] & t[122]);
  assign t[37] = t[119] ? x[29] : x[28];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = ~(t[61] & t[62]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = ~(t[65] & t[66]);
  assign t[42] = t[67] ^ t[41];
  assign t[43] = ~(t[123]);
  assign t[44] = ~(t[124]);
  assign t[45] = ~(t[68] & t[69]);
  assign t[46] = ~(t[22]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[125]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[75] & t[126]);
  assign t[51] = t[15] ? x[43] : x[42];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = ~(t[78] & t[127]);
  assign t[54] = t[15] ? x[48] : x[47];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[128]);
  assign t[57] = ~(t[129]);
  assign t[58] = ~(t[81] & t[82]);
  assign t[59] = ~(t[83] & t[84]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[85] & t[130]);
  assign t[61] = ~(t[86] & t[87]);
  assign t[62] = ~(t[88] & t[131]);
  assign t[63] = t[119] ? x[62] : x[61];
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[92]);
  assign t[66] = ~(t[93] & t[132]);
  assign t[67] = t[119] ? x[67] : x[66];
  assign t[68] = ~(t[124] & t[123]);
  assign t[69] = ~(t[133]);
  assign t[6] = ~(t[117] & t[118]);
  assign t[70] = ~(t[134]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[94] & t[95]);
  assign t[73] = ~(t[136]);
  assign t[74] = ~(t[137]);
  assign t[75] = ~(t[96] & t[97]);
  assign t[76] = ~(t[138]);
  assign t[77] = ~(t[139]);
  assign t[78] = ~(t[98] & t[99]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[119] & t[120]);
  assign t[80] = ~(t[102] & t[140]);
  assign t[81] = ~(t[129] & t[128]);
  assign t[82] = ~(t[141]);
  assign t[83] = ~(t[142]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[103] & t[104]);
  assign t[86] = ~(t[144]);
  assign t[87] = ~(t[145]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[109] & t[146]);
  assign t[91] = ~(t[147]);
  assign t[92] = ~(t[148]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[135] & t[134]);
  assign t[95] = ~(t[149]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[150]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[151]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[116];
endmodule

module R1ind188(x, y);
 input [121:0] x;
 output y;

 wire [166:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[135] ^ x[14];
  assign t[101] = t[136] ^ x[17];
  assign t[102] = t[137] ^ x[22];
  assign t[103] = t[138] ^ x[25];
  assign t[104] = t[139] ^ x[30];
  assign t[105] = t[140] ^ x[33];
  assign t[106] = t[141] ^ x[38];
  assign t[107] = t[142] ^ x[41];
  assign t[108] = t[143] ^ x[44];
  assign t[109] = t[144] ^ x[47];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[145] ^ x[50];
  assign t[111] = t[146] ^ x[55];
  assign t[112] = t[147] ^ x[58];
  assign t[113] = t[148] ^ x[63];
  assign t[114] = t[149] ^ x[66];
  assign t[115] = t[150] ^ x[69];
  assign t[116] = t[151] ^ x[72];
  assign t[117] = t[152] ^ x[75];
  assign t[118] = t[153] ^ x[80];
  assign t[119] = t[154] ^ x[83];
  assign t[11] = t[15] ? x[18] : x[19];
  assign t[120] = t[155] ^ x[88];
  assign t[121] = t[156] ^ x[91];
  assign t[122] = t[157] ^ x[94];
  assign t[123] = t[158] ^ x[97];
  assign t[124] = t[159] ^ x[100];
  assign t[125] = t[160] ^ x[103];
  assign t[126] = t[161] ^ x[106];
  assign t[127] = t[162] ^ x[109];
  assign t[128] = t[163] ^ x[112];
  assign t[129] = t[164] ^ x[115];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[165] ^ x[118];
  assign t[131] = t[166] ^ x[121];
  assign t[132] = (x[0] & x[1]);
  assign t[133] = (x[6] & x[7]);
  assign t[134] = (x[9] & x[10]);
  assign t[135] = (x[12] & x[13]);
  assign t[136] = (x[15] & x[16]);
  assign t[137] = (x[20] & x[21]);
  assign t[138] = (x[23] & x[24]);
  assign t[139] = (x[28] & x[29]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[31] & x[32]);
  assign t[141] = (x[36] & x[37]);
  assign t[142] = (x[39] & x[40]);
  assign t[143] = (x[42] & x[43]);
  assign t[144] = (x[45] & x[46]);
  assign t[145] = (x[48] & x[49]);
  assign t[146] = (x[53] & x[54]);
  assign t[147] = (x[56] & x[57]);
  assign t[148] = (x[61] & x[62]);
  assign t[149] = (x[64] & x[65]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (x[67] & x[68]);
  assign t[151] = (x[70] & x[71]);
  assign t[152] = (x[73] & x[74]);
  assign t[153] = (x[78] & x[79]);
  assign t[154] = (x[81] & x[82]);
  assign t[155] = (x[86] & x[87]);
  assign t[156] = (x[89] & x[90]);
  assign t[157] = (x[92] & x[93]);
  assign t[158] = (x[95] & x[96]);
  assign t[159] = (x[98] & x[99]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[101] & x[102]);
  assign t[161] = (x[104] & x[105]);
  assign t[162] = (x[107] & x[108]);
  assign t[163] = (x[110] & x[111]);
  assign t[164] = (x[113] & x[114]);
  assign t[165] = (x[116] & x[117]);
  assign t[166] = (x[119] & x[120]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[100]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[102] & t[43]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[29] = t[45] ? x[27] : x[26];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[41];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[104] & t[55]);
  assign t[36] = ~(t[105] & t[56]);
  assign t[37] = t[100] ? x[35] : x[34];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[61] ^ t[39];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[106]);
  assign t[44] = ~(t[106] & t[66]);
  assign t[45] = ~(t[22]);
  assign t[46] = ~(t[107] & t[67]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[71] ? x[52] : x[51];
  assign t[51] = ~(t[111] & t[72]);
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = t[71] ? x[60] : x[59];
  assign t[54] = ~(t[74] & t[75]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[113] & t[76]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = t[100] ? x[77] : x[76];
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = t[100] ? x[85] : x[84];
  assign t[65] = ~(t[83] & t[84]);
  assign t[66] = ~(t[102]);
  assign t[67] = ~(t[120]);
  assign t[68] = ~(t[120] & t[85]);
  assign t[69] = ~(t[121]);
  assign t[6] = ~(t[98] & t[99]);
  assign t[70] = ~(t[121] & t[86]);
  assign t[71] = ~(t[22]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[122] & t[87]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[104]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[100] & t[101]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[127] & t[92]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[130]);
  assign t[89] = ~(t[130] & t[95]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[114]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[118]);
  assign t[93] = ~(t[131]);
  assign t[94] = ~(t[131] & t[96]);
  assign t[95] = ~(t[123]);
  assign t[96] = ~(t[128]);
  assign t[97] = t[132] ^ x[2];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[11];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[97];
endmodule

module R1ind189(x, y);
 input [151:0] x;
 output y;

 wire [293:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[145] ? x[79] : x[78];
  assign t[101] = ~(t[146] & t[82]);
  assign t[102] = ~(t[227]);
  assign t[103] = ~(t[228]);
  assign t[104] = ~(t[147] | t[148]);
  assign t[105] = t[145] ? x[87] : x[86];
  assign t[106] = ~(t[149] & t[150]);
  assign t[107] = ~(t[229]);
  assign t[108] = ~(t[216] | t[217]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[151] | t[152]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[232]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[155] | t[156]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[234] | t[159]);
  assign t[118] = t[92] ? x[107] : x[106];
  assign t[119] = ~(t[160] & t[161]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[235]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = t[207] ? x[115] : x[114];
  assign t[124] = t[164] | t[165];
  assign t[125] = ~(t[166] & t[208]);
  assign t[126] = ~(t[167] & t[168]);
  assign t[127] = ~(t[79] | t[169]);
  assign t[128] = ~(t[79] | t[170]);
  assign t[129] = t[208] & t[171];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[167] | t[166];
  assign t[131] = ~(x[4] & t[172]);
  assign t[132] = ~(t[173] & t[168]);
  assign t[133] = t[205] ? t[175] : t[174];
  assign t[134] = ~(t[171] & t[176]);
  assign t[135] = ~(t[237]);
  assign t[136] = ~(t[222] | t[223]);
  assign t[137] = ~(t[207]);
  assign t[138] = ~(t[112]);
  assign t[139] = ~(t[79] | t[177]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[238]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[239]);
  assign t[143] = ~(t[240]);
  assign t[144] = ~(t[178] | t[179]);
  assign t[145] = ~(t[137]);
  assign t[146] = ~(t[164] | t[180]);
  assign t[147] = ~(t[241]);
  assign t[148] = ~(t[227] | t[228]);
  assign t[149] = ~(t[127] | t[181]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[182] & t[183]);
  assign t[151] = ~(t[242]);
  assign t[152] = ~(t[230] | t[231]);
  assign t[153] = ~(t[79] | t[184]);
  assign t[154] = ~(t[79] | t[185]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[232] | t[233]);
  assign t[157] = ~(t[244]);
  assign t[158] = ~(t[245]);
  assign t[159] = ~(t[186] | t[187]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(t[164] | t[188]);
  assign t[161] = ~(t[47]);
  assign t[162] = ~(t[246]);
  assign t[163] = ~(t[235] | t[236]);
  assign t[164] = ~(t[134] & t[150]);
  assign t[165] = ~(t[189] & t[190]);
  assign t[166] = x[4] & t[206];
  assign t[167] = ~(x[4] | t[206]);
  assign t[168] = ~(t[208]);
  assign t[169] = t[205] ? t[125] : t[126];
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = t[205] ? t[131] : t[191];
  assign t[171] = ~(t[83] | t[205]);
  assign t[172] = ~(t[206] | t[208]);
  assign t[173] = ~(x[4] | t[192]);
  assign t[174] = ~(t[166] & t[168]);
  assign t[175] = ~(t[167] & t[208]);
  assign t[176] = ~(t[191] & t[193]);
  assign t[177] = t[205] ? t[191] : t[131];
  assign t[178] = ~(t[247]);
  assign t[179] = ~(t[239] | t[240]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = t[139] | t[85];
  assign t[181] = ~(t[194] & t[195]);
  assign t[182] = ~(t[206] | t[168]);
  assign t[183] = t[79] & t[205];
  assign t[184] = t[205] ? t[193] : t[132];
  assign t[185] = t[205] ? t[174] : t[175];
  assign t[186] = ~(t[248]);
  assign t[187] = ~(t[244] | t[245]);
  assign t[188] = ~(t[196] & t[197]);
  assign t[189] = ~(t[47] | t[85]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[128] | t[154]);
  assign t[191] = ~(t[208] & t[173]);
  assign t[192] = ~(t[206]);
  assign t[193] = ~(x[4] & t[182]);
  assign t[194] = ~(t[198] | t[199]);
  assign t[195] = ~(t[83] & t[200]);
  assign t[196] = ~(t[49]);
  assign t[197] = t[83] | t[201];
  assign t[198] = ~(t[83] | t[202]);
  assign t[199] = ~(t[79] | t[203]);
  assign t[19] = t[207] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[131] & t[191]);
  assign t[201] = t[205] ? t[131] : t[132];
  assign t[202] = t[205] ? t[126] : t[174];
  assign t[203] = t[205] ? t[132] : t[193];
  assign t[204] = t[249] ^ x[2];
  assign t[205] = t[250] ^ x[10];
  assign t[206] = t[251] ^ x[13];
  assign t[207] = t[252] ^ x[16];
  assign t[208] = t[253] ^ x[19];
  assign t[209] = t[254] ^ x[22];
  assign t[20] = ~(t[29] & t[30]);
  assign t[210] = t[255] ^ x[25];
  assign t[211] = t[256] ^ x[28];
  assign t[212] = t[257] ^ x[31];
  assign t[213] = t[258] ^ x[34];
  assign t[214] = t[259] ^ x[39];
  assign t[215] = t[260] ^ x[42];
  assign t[216] = t[261] ^ x[45];
  assign t[217] = t[262] ^ x[48];
  assign t[218] = t[263] ^ x[51];
  assign t[219] = t[264] ^ x[56];
  assign t[21] = ~(t[31] | t[32]);
  assign t[220] = t[265] ^ x[59];
  assign t[221] = t[266] ^ x[62];
  assign t[222] = t[267] ^ x[65];
  assign t[223] = t[268] ^ x[68];
  assign t[224] = t[269] ^ x[71];
  assign t[225] = t[270] ^ x[74];
  assign t[226] = t[271] ^ x[77];
  assign t[227] = t[272] ^ x[82];
  assign t[228] = t[273] ^ x[85];
  assign t[229] = t[274] ^ x[90];
  assign t[22] = ~(t[33] ^ t[34]);
  assign t[230] = t[275] ^ x[93];
  assign t[231] = t[276] ^ x[96];
  assign t[232] = t[277] ^ x[99];
  assign t[233] = t[278] ^ x[102];
  assign t[234] = t[279] ^ x[105];
  assign t[235] = t[280] ^ x[110];
  assign t[236] = t[281] ^ x[113];
  assign t[237] = t[282] ^ x[118];
  assign t[238] = t[283] ^ x[121];
  assign t[239] = t[284] ^ x[124];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[285] ^ x[127];
  assign t[241] = t[286] ^ x[130];
  assign t[242] = t[287] ^ x[133];
  assign t[243] = t[288] ^ x[136];
  assign t[244] = t[289] ^ x[139];
  assign t[245] = t[290] ^ x[142];
  assign t[246] = t[291] ^ x[145];
  assign t[247] = t[292] ^ x[148];
  assign t[248] = t[293] ^ x[151];
  assign t[249] = (x[0] & x[1]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[8] & x[9]);
  assign t[251] = (x[11] & x[12]);
  assign t[252] = (x[14] & x[15]);
  assign t[253] = (x[17] & x[18]);
  assign t[254] = (x[20] & x[21]);
  assign t[255] = (x[23] & x[24]);
  assign t[256] = (x[26] & x[27]);
  assign t[257] = (x[29] & x[30]);
  assign t[258] = (x[32] & x[33]);
  assign t[259] = (x[37] & x[38]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[40] & x[41]);
  assign t[261] = (x[43] & x[44]);
  assign t[262] = (x[46] & x[47]);
  assign t[263] = (x[49] & x[50]);
  assign t[264] = (x[54] & x[55]);
  assign t[265] = (x[57] & x[58]);
  assign t[266] = (x[60] & x[61]);
  assign t[267] = (x[63] & x[64]);
  assign t[268] = (x[66] & x[67]);
  assign t[269] = (x[69] & x[70]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[72] & x[73]);
  assign t[271] = (x[75] & x[76]);
  assign t[272] = (x[80] & x[81]);
  assign t[273] = (x[83] & x[84]);
  assign t[274] = (x[88] & x[89]);
  assign t[275] = (x[91] & x[92]);
  assign t[276] = (x[94] & x[95]);
  assign t[277] = (x[97] & x[98]);
  assign t[278] = (x[100] & x[101]);
  assign t[279] = (x[103] & x[104]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[108] & x[109]);
  assign t[281] = (x[111] & x[112]);
  assign t[282] = (x[116] & x[117]);
  assign t[283] = (x[119] & x[120]);
  assign t[284] = (x[122] & x[123]);
  assign t[285] = (x[125] & x[126]);
  assign t[286] = (x[128] & x[129]);
  assign t[287] = (x[131] & x[132]);
  assign t[288] = (x[134] & x[135]);
  assign t[289] = (x[137] & x[138]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = (x[140] & x[141]);
  assign t[291] = (x[143] & x[144]);
  assign t[292] = (x[146] & x[147]);
  assign t[293] = (x[149] & x[150]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[209] | t[53]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[34] = ~(t[56] ^ t[57]);
  assign t[35] = ~(t[58] | t[59]);
  assign t[36] = ~(t[60] ^ t[61]);
  assign t[37] = ~(t[62] | t[63]);
  assign t[38] = ~(t[43] ^ t[64]);
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[210] | t[67]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[42] = ~(t[70] ^ t[71]);
  assign t[43] = ~(t[72] | t[73]);
  assign t[44] = ~(t[74] ^ t[75]);
  assign t[45] = ~(t[76] | t[77]);
  assign t[46] = ~(t[45] ^ t[78]);
  assign t[47] = ~(t[79] | t[80]);
  assign t[48] = ~(t[81] & t[82]);
  assign t[49] = ~(t[83] | t[84]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[85] | t[86];
  assign t[51] = ~(t[211]);
  assign t[52] = ~(t[212]);
  assign t[53] = ~(t[87] | t[88]);
  assign t[54] = ~(t[89] | t[90]);
  assign t[55] = ~(t[213] | t[91]);
  assign t[56] = t[92] ? x[36] : x[35];
  assign t[57] = ~(t[93] & t[94]);
  assign t[58] = ~(t[95] | t[96]);
  assign t[59] = ~(t[214] | t[97]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[98] | t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = ~(t[102] | t[103]);
  assign t[63] = ~(t[215] | t[104]);
  assign t[64] = ~(t[105] ^ t[106]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[107] | t[108]);
  assign t[68] = ~(t[109] | t[110]);
  assign t[69] = ~(t[218] | t[111]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[207] ? x[53] : x[52];
  assign t[71] = ~(t[29] & t[112]);
  assign t[72] = ~(t[113] | t[114]);
  assign t[73] = ~(t[219] | t[115]);
  assign t[74] = ~(t[116] | t[117]);
  assign t[75] = ~(t[118] ^ t[119]);
  assign t[76] = ~(t[120] | t[121]);
  assign t[77] = ~(t[220] | t[122]);
  assign t[78] = ~(t[123] ^ t[124]);
  assign t[79] = ~(t[83]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[205] ? t[126] : t[125];
  assign t[81] = ~(t[127] | t[128]);
  assign t[82] = ~(t[129] & t[130]);
  assign t[83] = ~(t[207]);
  assign t[84] = t[205] ? t[132] : t[131];
  assign t[85] = ~(t[79] | t[133]);
  assign t[86] = ~(t[134]);
  assign t[87] = ~(t[221]);
  assign t[88] = ~(t[211] | t[212]);
  assign t[89] = ~(t[222]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[135] | t[136]);
  assign t[92] = ~(t[137]);
  assign t[93] = ~(t[127]);
  assign t[94] = ~(t[138] | t[139]);
  assign t[95] = ~(t[224]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[140] | t[141]);
  assign t[98] = ~(t[142] | t[143]);
  assign t[99] = ~(t[226] | t[144]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind190(x, y);
 input [139:0] x;
 output y;

 wire [180:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[141] ^ x[8];
  assign t[101] = t[142] ^ x[11];
  assign t[102] = t[143] ^ x[14];
  assign t[103] = t[144] ^ x[17];
  assign t[104] = t[145] ^ x[22];
  assign t[105] = t[146] ^ x[27];
  assign t[106] = t[147] ^ x[32];
  assign t[107] = t[148] ^ x[35];
  assign t[108] = t[149] ^ x[38];
  assign t[109] = t[150] ^ x[43];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[48];
  assign t[111] = t[152] ^ x[51];
  assign t[112] = t[153] ^ x[54];
  assign t[113] = t[154] ^ x[57];
  assign t[114] = t[155] ^ x[62];
  assign t[115] = t[156] ^ x[67];
  assign t[116] = t[157] ^ x[70];
  assign t[117] = t[158] ^ x[73];
  assign t[118] = t[159] ^ x[76];
  assign t[119] = t[160] ^ x[79];
  assign t[11] = t[102] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[82];
  assign t[121] = t[162] ^ x[85];
  assign t[122] = t[163] ^ x[88];
  assign t[123] = t[164] ^ x[91];
  assign t[124] = t[165] ^ x[94];
  assign t[125] = t[166] ^ x[97];
  assign t[126] = t[167] ^ x[100];
  assign t[127] = t[168] ^ x[103];
  assign t[128] = t[169] ^ x[106];
  assign t[129] = t[170] ^ x[109];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[112];
  assign t[131] = t[172] ^ x[115];
  assign t[132] = t[173] ^ x[118];
  assign t[133] = t[174] ^ x[121];
  assign t[134] = t[175] ^ x[124];
  assign t[135] = t[176] ^ x[127];
  assign t[136] = t[177] ^ x[130];
  assign t[137] = t[178] ^ x[133];
  assign t[138] = t[179] ^ x[136];
  assign t[139] = t[180] ^ x[139];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[0] & x[1]);
  assign t[141] = (x[6] & x[7]);
  assign t[142] = (x[9] & x[10]);
  assign t[143] = (x[12] & x[13]);
  assign t[144] = (x[15] & x[16]);
  assign t[145] = (x[20] & x[21]);
  assign t[146] = (x[25] & x[26]);
  assign t[147] = (x[30] & x[31]);
  assign t[148] = (x[33] & x[34]);
  assign t[149] = (x[36] & x[37]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[41] & x[42]);
  assign t[151] = (x[46] & x[47]);
  assign t[152] = (x[49] & x[50]);
  assign t[153] = (x[52] & x[53]);
  assign t[154] = (x[55] & x[56]);
  assign t[155] = (x[60] & x[61]);
  assign t[156] = (x[65] & x[66]);
  assign t[157] = (x[68] & x[69]);
  assign t[158] = (x[71] & x[72]);
  assign t[159] = (x[74] & x[75]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[77] & x[78]);
  assign t[161] = (x[80] & x[81]);
  assign t[162] = (x[83] & x[84]);
  assign t[163] = (x[86] & x[87]);
  assign t[164] = (x[89] & x[90]);
  assign t[165] = (x[92] & x[93]);
  assign t[166] = (x[95] & x[96]);
  assign t[167] = (x[98] & x[99]);
  assign t[168] = (x[101] & x[102]);
  assign t[169] = (x[104] & x[105]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[107] & x[108]);
  assign t[171] = (x[110] & x[111]);
  assign t[172] = (x[113] & x[114]);
  assign t[173] = (x[116] & x[117]);
  assign t[174] = (x[119] & x[120]);
  assign t[175] = (x[122] & x[123]);
  assign t[176] = (x[125] & x[126]);
  assign t[177] = (x[128] & x[129]);
  assign t[178] = (x[131] & x[132]);
  assign t[179] = (x[134] & x[135]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[137] & x[138]);
  assign t[18] = t[27] ^ t[21];
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = t[42] | t[104];
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = t[46] ^ t[28];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = t[49] ^ t[50];
  assign t[32] = ~(t[51] & t[52]);
  assign t[33] = t[53] | t[105];
  assign t[34] = t[54] ? x[29] : x[28];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = ~(t[57] & t[58]);
  assign t[37] = t[59] ^ t[60];
  assign t[38] = ~(t[61] & t[62]);
  assign t[39] = t[63] ^ t[38];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[106]);
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[64] | t[40]);
  assign t[43] = ~(t[65]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] | t[108];
  assign t[46] = t[43] ? x[40] : x[39];
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[109];
  assign t[49] = t[43] ? x[45] : x[44];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[110]);
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[74] | t[51]);
  assign t[54] = ~(t[65]);
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = t[77] | t[112];
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = t[80] | t[113];
  assign t[59] = t[102] ? x[59] : x[58];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = t[85] | t[114];
  assign t[63] = t[102] ? x[64] : x[63];
  assign t[64] = ~(t[115]);
  assign t[65] = ~(t[102]);
  assign t[66] = ~(t[116]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[86] | t[66]);
  assign t[69] = ~(t[118]);
  assign t[6] = ~(t[100] & t[101]);
  assign t[70] = ~(t[119]);
  assign t[71] = ~(t[87] | t[69]);
  assign t[72] = ~(t[88] & t[89]);
  assign t[73] = t[90] | t[120];
  assign t[74] = ~(t[121]);
  assign t[75] = ~(t[122]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[91] | t[75]);
  assign t[78] = ~(t[124]);
  assign t[79] = ~(t[125]);
  assign t[7] = ~(t[102] & t[103]);
  assign t[80] = ~(t[92] | t[78]);
  assign t[81] = ~(t[93] & t[94]);
  assign t[82] = t[95] | t[126];
  assign t[83] = ~(t[127]);
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[96] | t[83]);
  assign t[86] = ~(t[129]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[97] | t[88]);
  assign t[91] = ~(t[133]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[98] | t[93]);
  assign t[96] = ~(t[137]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = t[140] ^ x[2];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind191(x, y);
 input [139:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[108] & t[109]);
  assign t[104] = ~(t[139] & t[138]);
  assign t[105] = ~(t[148]);
  assign t[106] = ~(t[143] & t[142]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[147] & t[146]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[32];
  assign t[118] = t[159] ^ x[35];
  assign t[119] = t[160] ^ x[38];
  assign t[11] = t[111] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[43];
  assign t[121] = t[162] ^ x[48];
  assign t[122] = t[163] ^ x[51];
  assign t[123] = t[164] ^ x[54];
  assign t[124] = t[165] ^ x[57];
  assign t[125] = t[166] ^ x[62];
  assign t[126] = t[167] ^ x[67];
  assign t[127] = t[168] ^ x[70];
  assign t[128] = t[169] ^ x[73];
  assign t[129] = t[170] ^ x[76];
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = t[171] ^ x[79];
  assign t[131] = t[172] ^ x[82];
  assign t[132] = t[173] ^ x[85];
  assign t[133] = t[174] ^ x[88];
  assign t[134] = t[175] ^ x[91];
  assign t[135] = t[176] ^ x[94];
  assign t[136] = t[177] ^ x[97];
  assign t[137] = t[178] ^ x[100];
  assign t[138] = t[179] ^ x[103];
  assign t[139] = t[180] ^ x[106];
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = t[181] ^ x[109];
  assign t[141] = t[182] ^ x[112];
  assign t[142] = t[183] ^ x[115];
  assign t[143] = t[184] ^ x[118];
  assign t[144] = t[185] ^ x[121];
  assign t[145] = t[186] ^ x[124];
  assign t[146] = t[187] ^ x[127];
  assign t[147] = t[188] ^ x[130];
  assign t[148] = t[189] ^ x[133];
  assign t[149] = t[190] ^ x[136];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = t[191] ^ x[139];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[30] & x[31]);
  assign t[159] = (x[33] & x[34]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[36] & x[37]);
  assign t[161] = (x[41] & x[42]);
  assign t[162] = (x[46] & x[47]);
  assign t[163] = (x[49] & x[50]);
  assign t[164] = (x[52] & x[53]);
  assign t[165] = (x[55] & x[56]);
  assign t[166] = (x[60] & x[61]);
  assign t[167] = (x[65] & x[66]);
  assign t[168] = (x[68] & x[69]);
  assign t[169] = (x[71] & x[72]);
  assign t[16] = ~(t[111] & t[114]);
  assign t[170] = (x[74] & x[75]);
  assign t[171] = (x[77] & x[78]);
  assign t[172] = (x[80] & x[81]);
  assign t[173] = (x[83] & x[84]);
  assign t[174] = (x[86] & x[87]);
  assign t[175] = (x[89] & x[90]);
  assign t[176] = (x[92] & x[93]);
  assign t[177] = (x[95] & x[96]);
  assign t[178] = (x[98] & x[99]);
  assign t[179] = (x[101] & x[102]);
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = (x[104] & x[105]);
  assign t[181] = (x[107] & x[108]);
  assign t[182] = (x[110] & x[111]);
  assign t[183] = (x[113] & x[114]);
  assign t[184] = (x[116] & x[117]);
  assign t[185] = (x[119] & x[120]);
  assign t[186] = (x[122] & x[123]);
  assign t[187] = (x[125] & x[126]);
  assign t[188] = (x[128] & x[129]);
  assign t[189] = (x[131] & x[132]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = (x[134] & x[135]);
  assign t[191] = (x[137] & x[138]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ t[23];
  assign t[21] = x[4] ? t[31] : t[30];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = ~(t[34] & t[35]);
  assign t[24] = t[36] ^ t[37];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[27] = ~(t[42] & t[43]);
  assign t[28] = ~(t[44] & t[115]);
  assign t[29] = t[45] ? x[24] : x[23];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = t[48] ^ t[30];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = ~(t[53] & t[54]);
  assign t[35] = ~(t[55] & t[116]);
  assign t[36] = t[56] ? x[29] : x[28];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[63] & t[64]);
  assign t[41] = t[65] ^ t[40];
  assign t[42] = ~(t[117]);
  assign t[43] = ~(t[118]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = ~(t[68]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[119]);
  assign t[48] = t[45] ? x[40] : x[39];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[120]);
  assign t[51] = t[45] ? x[45] : x[44];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = ~(t[121]);
  assign t[54] = ~(t[122]);
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[68]);
  assign t[57] = ~(t[79] & t[80]);
  assign t[58] = ~(t[81] & t[123]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[124]);
  assign t[61] = t[111] ? x[59] : x[58];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[125]);
  assign t[65] = t[111] ? x[64] : x[63];
  assign t[66] = ~(t[118] & t[117]);
  assign t[67] = ~(t[126]);
  assign t[68] = ~(t[111]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = ~(t[129]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[92] & t[93]);
  assign t[75] = ~(t[94] & t[95]);
  assign t[76] = ~(t[96] & t[131]);
  assign t[77] = ~(t[122] & t[121]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[97] & t[98]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[101] & t[102]);
  assign t[86] = ~(t[103] & t[137]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[106] & t[107]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind192(x, y);
 input [112:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[132] ^ x[44];
  assign t[101] = t[133] ^ x[49];
  assign t[102] = t[134] ^ x[52];
  assign t[103] = t[135] ^ x[57];
  assign t[104] = t[136] ^ x[60];
  assign t[105] = t[137] ^ x[63];
  assign t[106] = t[138] ^ x[66];
  assign t[107] = t[139] ^ x[69];
  assign t[108] = t[140] ^ x[74];
  assign t[109] = t[141] ^ x[77];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[142] ^ x[82];
  assign t[111] = t[143] ^ x[85];
  assign t[112] = t[144] ^ x[88];
  assign t[113] = t[145] ^ x[91];
  assign t[114] = t[146] ^ x[94];
  assign t[115] = t[147] ^ x[97];
  assign t[116] = t[148] ^ x[100];
  assign t[117] = t[149] ^ x[103];
  assign t[118] = t[150] ^ x[106];
  assign t[119] = t[151] ^ x[109];
  assign t[11] = t[92] ? x[18] : x[19];
  assign t[120] = t[152] ^ x[112];
  assign t[121] = (x[0] & x[1]);
  assign t[122] = (x[6] & x[7]);
  assign t[123] = (x[9] & x[10]);
  assign t[124] = (x[12] & x[13]);
  assign t[125] = (x[15] & x[16]);
  assign t[126] = (x[20] & x[21]);
  assign t[127] = (x[23] & x[24]);
  assign t[128] = (x[28] & x[29]);
  assign t[129] = (x[31] & x[32]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = (x[36] & x[37]);
  assign t[131] = (x[39] & x[40]);
  assign t[132] = (x[42] & x[43]);
  assign t[133] = (x[47] & x[48]);
  assign t[134] = (x[50] & x[51]);
  assign t[135] = (x[55] & x[56]);
  assign t[136] = (x[58] & x[59]);
  assign t[137] = (x[61] & x[62]);
  assign t[138] = (x[64] & x[65]);
  assign t[139] = (x[67] & x[68]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[72] & x[73]);
  assign t[141] = (x[75] & x[76]);
  assign t[142] = (x[80] & x[81]);
  assign t[143] = (x[83] & x[84]);
  assign t[144] = (x[86] & x[87]);
  assign t[145] = (x[89] & x[90]);
  assign t[146] = (x[92] & x[93]);
  assign t[147] = (x[95] & x[96]);
  assign t[148] = (x[98] & x[99]);
  assign t[149] = (x[101] & x[102]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[104] & x[105]);
  assign t[151] = (x[107] & x[108]);
  assign t[152] = (x[110] & x[111]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] ^ t[21];
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[94] & t[40]);
  assign t[26] = ~(t[95] & t[41]);
  assign t[27] = t[42] ? x[27] : x[26];
  assign t[28] = ~(t[43] & t[44]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = t[49] ^ t[30];
  assign t[32] = ~(t[96] & t[50]);
  assign t[33] = ~(t[97] & t[51]);
  assign t[34] = t[42] ? x[35] : x[34];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[36];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[98]);
  assign t[41] = ~(t[98] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[99] & t[63]);
  assign t[44] = ~(t[100] & t[64]);
  assign t[45] = t[42] ? x[46] : x[45];
  assign t[46] = ~(t[65] & t[66]);
  assign t[47] = ~(t[101] & t[67]);
  assign t[48] = ~(t[102] & t[68]);
  assign t[49] = t[42] ? x[54] : x[53];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[103]);
  assign t[51] = ~(t[103] & t[69]);
  assign t[52] = ~(t[104] & t[70]);
  assign t[53] = ~(t[105] & t[71]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = t[92] ? x[71] : x[70];
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = t[92] ? x[79] : x[78];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[76] & t[77]);
  assign t[61] = ~(t[94]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[110]);
  assign t[64] = ~(t[110] & t[78]);
  assign t[65] = ~(t[111] & t[79]);
  assign t[66] = ~(t[112] & t[80]);
  assign t[67] = ~(t[113]);
  assign t[68] = ~(t[113] & t[81]);
  assign t[69] = ~(t[96]);
  assign t[6] = ~(t[90] & t[91]);
  assign t[70] = ~(t[114]);
  assign t[71] = ~(t[114] & t[82]);
  assign t[72] = ~(t[115]);
  assign t[73] = ~(t[115] & t[83]);
  assign t[74] = ~(t[116]);
  assign t[75] = ~(t[116] & t[84]);
  assign t[76] = ~(t[117] & t[85]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[99]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[92] & t[93]);
  assign t[80] = ~(t[119] & t[87]);
  assign t[81] = ~(t[101]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[106]);
  assign t[84] = ~(t[108]);
  assign t[85] = ~(t[120]);
  assign t[86] = ~(t[120] & t[88]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[117]);
  assign t[89] = t[121] ^ x[2];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[122] ^ x[8];
  assign t[91] = t[123] ^ x[11];
  assign t[92] = t[124] ^ x[14];
  assign t[93] = t[125] ^ x[17];
  assign t[94] = t[126] ^ x[22];
  assign t[95] = t[127] ^ x[25];
  assign t[96] = t[128] ^ x[30];
  assign t[97] = t[129] ^ x[33];
  assign t[98] = t[130] ^ x[38];
  assign t[99] = t[131] ^ x[41];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[89];
endmodule

module R1ind193(x, y);
 input [139:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[211] | t[212]);
  assign t[101] = ~(t[223]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[141] | t[142]);
  assign t[104] = ~(t[143] | t[144]);
  assign t[105] = ~(t[225]);
  assign t[106] = ~(t[226]);
  assign t[107] = ~(t[145] | t[146]);
  assign t[108] = ~(t[147] | t[148]);
  assign t[109] = ~(t[227] | t[149]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[150] ? x[98] : x[97];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = ~(t[228]);
  assign t[113] = ~(t[229]);
  assign t[114] = ~(t[153] | t[154]);
  assign t[115] = t[203] ? x[106] : x[105];
  assign t[116] = t[155] | t[156];
  assign t[117] = ~(t[203]);
  assign t[118] = ~(t[157] & t[204]);
  assign t[119] = ~(t[158] & t[159]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[76] | t[160]);
  assign t[121] = ~(t[76] | t[161]);
  assign t[122] = t[204] & t[162];
  assign t[123] = t[158] | t[157];
  assign t[124] = ~(t[163] & t[159]);
  assign t[125] = ~(x[4] & t[164]);
  assign t[126] = ~(t[158] & t[204]);
  assign t[127] = ~(t[157] & t[159]);
  assign t[128] = ~(t[203]);
  assign t[129] = ~(t[139]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[230]);
  assign t[131] = ~(t[217] | t[218]);
  assign t[132] = ~(t[165] | t[143]);
  assign t[133] = ~(t[166] | t[167]);
  assign t[134] = ~(t[231]);
  assign t[135] = ~(t[219] | t[220]);
  assign t[136] = ~(t[232]);
  assign t[137] = ~(t[233]);
  assign t[138] = ~(t[168] | t[169]);
  assign t[139] = ~(t[170] | t[143]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[171] | t[172]);
  assign t[141] = ~(t[234]);
  assign t[142] = ~(t[223] | t[224]);
  assign t[143] = ~(t[117] | t[173]);
  assign t[144] = t[174] | t[175];
  assign t[145] = ~(t[235]);
  assign t[146] = ~(t[225] | t[226]);
  assign t[147] = ~(t[236]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[128]);
  assign t[151] = ~(t[155] | t[178]);
  assign t[152] = ~(t[46]);
  assign t[153] = ~(t[238]);
  assign t[154] = ~(t[228] | t[229]);
  assign t[155] = ~(t[179] & t[180]);
  assign t[156] = ~(t[181] & t[85]);
  assign t[157] = x[4] & t[202];
  assign t[158] = ~(x[4] | t[202]);
  assign t[159] = ~(t[204]);
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = t[201] ? t[118] : t[119];
  assign t[161] = t[201] ? t[183] : t[182];
  assign t[162] = ~(t[117] | t[201]);
  assign t[163] = ~(x[4] | t[184]);
  assign t[164] = ~(t[202] | t[159]);
  assign t[165] = ~(t[117] | t[185]);
  assign t[166] = ~(t[30]);
  assign t[167] = ~(t[76] | t[186]);
  assign t[168] = ~(t[239]);
  assign t[169] = ~(t[232] | t[233]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[117] | t[187]);
  assign t[171] = ~(t[188] & t[189]);
  assign t[172] = ~(t[79] & t[190]);
  assign t[173] = t[201] ? t[124] : t[183];
  assign t[174] = ~(t[76] | t[191]);
  assign t[175] = ~(t[179]);
  assign t[176] = ~(t[240]);
  assign t[177] = ~(t[236] | t[237]);
  assign t[178] = ~(t[192] & t[190]);
  assign t[179] = ~(t[162] & t[193]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[164] & t[194]);
  assign t[181] = ~(t[46] | t[174]);
  assign t[182] = ~(t[204] & t[163]);
  assign t[183] = ~(x[4] & t[195]);
  assign t[184] = ~(t[202]);
  assign t[185] = t[201] ? t[119] : t[127];
  assign t[186] = t[201] ? t[182] : t[183];
  assign t[187] = t[201] ? t[127] : t[119];
  assign t[188] = ~(t[165] | t[196]);
  assign t[189] = ~(t[117] & t[197]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[117] | t[198];
  assign t[191] = t[201] ? t[126] : t[127];
  assign t[192] = ~(t[143]);
  assign t[193] = ~(t[182] & t[125]);
  assign t[194] = t[76] & t[201];
  assign t[195] = ~(t[202] | t[204]);
  assign t[196] = ~(t[76] | t[199]);
  assign t[197] = ~(t[183] & t[182]);
  assign t[198] = t[201] ? t[183] : t[124];
  assign t[199] = t[201] ? t[124] : t[125];
  assign t[19] = t[203] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[10];
  assign t[202] = t[243] ^ x[13];
  assign t[203] = t[244] ^ x[16];
  assign t[204] = t[245] ^ x[19];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[28];
  assign t[208] = t[249] ^ x[31];
  assign t[209] = t[250] ^ x[36];
  assign t[20] = ~(t[29] & t[30]);
  assign t[210] = t[251] ^ x[39];
  assign t[211] = t[252] ^ x[42];
  assign t[212] = t[253] ^ x[45];
  assign t[213] = t[254] ^ x[48];
  assign t[214] = t[255] ^ x[53];
  assign t[215] = t[256] ^ x[56];
  assign t[216] = t[257] ^ x[59];
  assign t[217] = t[258] ^ x[62];
  assign t[218] = t[259] ^ x[65];
  assign t[219] = t[260] ^ x[70];
  assign t[21] = ~(t[31] | t[32]);
  assign t[220] = t[261] ^ x[73];
  assign t[221] = t[262] ^ x[76];
  assign t[222] = t[263] ^ x[81];
  assign t[223] = t[264] ^ x[84];
  assign t[224] = t[265] ^ x[87];
  assign t[225] = t[266] ^ x[90];
  assign t[226] = t[267] ^ x[93];
  assign t[227] = t[268] ^ x[96];
  assign t[228] = t[269] ^ x[101];
  assign t[229] = t[270] ^ x[104];
  assign t[22] = ~(t[25] ^ t[33]);
  assign t[230] = t[271] ^ x[109];
  assign t[231] = t[272] ^ x[112];
  assign t[232] = t[273] ^ x[115];
  assign t[233] = t[274] ^ x[118];
  assign t[234] = t[275] ^ x[121];
  assign t[235] = t[276] ^ x[124];
  assign t[236] = t[277] ^ x[127];
  assign t[237] = t[278] ^ x[130];
  assign t[238] = t[279] ^ x[133];
  assign t[239] = t[280] ^ x[136];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[281] ^ x[139];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[8] & x[9]);
  assign t[243] = (x[11] & x[12]);
  assign t[244] = (x[14] & x[15]);
  assign t[245] = (x[17] & x[18]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[26] & x[27]);
  assign t[249] = (x[29] & x[30]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (x[34] & x[35]);
  assign t[251] = (x[37] & x[38]);
  assign t[252] = (x[40] & x[41]);
  assign t[253] = (x[43] & x[44]);
  assign t[254] = (x[46] & x[47]);
  assign t[255] = (x[51] & x[52]);
  assign t[256] = (x[54] & x[55]);
  assign t[257] = (x[57] & x[58]);
  assign t[258] = (x[60] & x[61]);
  assign t[259] = (x[63] & x[64]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = (x[68] & x[69]);
  assign t[261] = (x[71] & x[72]);
  assign t[262] = (x[74] & x[75]);
  assign t[263] = (x[79] & x[80]);
  assign t[264] = (x[82] & x[83]);
  assign t[265] = (x[85] & x[86]);
  assign t[266] = (x[88] & x[89]);
  assign t[267] = (x[91] & x[92]);
  assign t[268] = (x[94] & x[95]);
  assign t[269] = (x[99] & x[100]);
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = (x[102] & x[103]);
  assign t[271] = (x[107] & x[108]);
  assign t[272] = (x[110] & x[111]);
  assign t[273] = (x[113] & x[114]);
  assign t[274] = (x[116] & x[117]);
  assign t[275] = (x[119] & x[120]);
  assign t[276] = (x[122] & x[123]);
  assign t[277] = (x[125] & x[126]);
  assign t[278] = (x[128] & x[129]);
  assign t[279] = (x[131] & x[132]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[134] & x[135]);
  assign t[281] = (x[137] & x[138]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[205] | t[52]);
  assign t[33] = ~(t[53] ^ t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[34] ^ t[57]);
  assign t[36] = ~(t[58] | t[59]);
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[206] | t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[67] ^ t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[44] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] & t[79]);
  assign t[48] = ~(t[76] | t[80]);
  assign t[49] = ~(t[76] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[207]);
  assign t[51] = ~(t[208]);
  assign t[52] = ~(t[82] | t[83]);
  assign t[53] = t[84] ? x[33] : x[32];
  assign t[54] = ~(t[85] & t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[209] | t[89]);
  assign t[57] = ~(t[90] ^ t[91]);
  assign t[58] = ~(t[92] | t[93]);
  assign t[59] = ~(t[210] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[97] ^ t[98]);
  assign t[62] = ~(t[211]);
  assign t[63] = ~(t[212]);
  assign t[64] = ~(t[99] | t[100]);
  assign t[65] = ~(t[101] | t[102]);
  assign t[66] = ~(t[213] | t[103]);
  assign t[67] = t[203] ? x[50] : x[49];
  assign t[68] = ~(t[29] & t[104]);
  assign t[69] = ~(t[105] | t[106]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[214] | t[107]);
  assign t[71] = ~(t[108] | t[109]);
  assign t[72] = ~(t[110] ^ t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[215] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117]);
  assign t[77] = t[201] ? t[119] : t[118];
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[122] & t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[201] ? t[125] : t[124];
  assign t[81] = t[201] ? t[127] : t[126];
  assign t[82] = ~(t[216]);
  assign t[83] = ~(t[207] | t[208]);
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[121] | t[49]);
  assign t[86] = ~(t[122] | t[129]);
  assign t[87] = ~(t[217]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[84] ? x[67] : x[66];
  assign t[91] = ~(t[132] & t[133]);
  assign t[92] = ~(t[219]);
  assign t[93] = ~(t[220]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[136] | t[137]);
  assign t[96] = ~(t[221] | t[138]);
  assign t[97] = t[84] ? x[78] : x[77];
  assign t[98] = ~(t[139] & t[140]);
  assign t[99] = ~(t[222]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind194(x, y);
 input [12:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[10] ^ t[1];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = (x[1] & x[2]);
  assign t[15] = (x[4] & x[5]);
  assign t[16] = (x[7] & x[8]);
  assign t[17] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[11]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[5] & t[13]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = ~(t[13] & t[12]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind195(x, y);
 input [12:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[9] ^ t[1]);
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[9];
  assign t[12] = t[16] ^ x[12];
  assign t[13] = (x[1] & x[2]);
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[10] & x[11]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[10]);
  assign t[3] = ~(t[4] & t[11]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(x[0]);
  assign t[7] = ~(t[9] & t[12]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = t[13] ^ x[3];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind196(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = t[7] ^ t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[8] & t[7]);
  assign t[7] = t[11] ^ x[3];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[9];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind197(x, y);
 input [12:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[6] ^ t[1]);
  assign t[10] = (x[1] & x[2]);
  assign t[11] = (x[4] & x[5]);
  assign t[12] = (x[7] & x[8]);
  assign t[13] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[0]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[6] & t[9]);
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[6];
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[12];
  assign y = ~(x[0] | t[0]);
endmodule

module R1_ind(x, y);
 input [592:0] x;
 output [197:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[210], x[209]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[202], x[201], x[200], x[205], x[204], x[203], x[208], x[207], x[206], x[212], x[211]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[205], x[204], x[203], x[202], x[201], x[200], x[208], x[207], x[206], x[199], x[198], x[197], x[214], x[213]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[230], x[229]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[222], x[221], x[220], x[225], x[224], x[223], x[228], x[227], x[226], x[232], x[231]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[225], x[224], x[223], x[222], x[221], x[220], x[228], x[227], x[226], x[219], x[218], x[217], x[234], x[233]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[250], x[249]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[242], x[241], x[240], x[245], x[244], x[243], x[248], x[247], x[246], x[252], x[251]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[245], x[244], x[243], x[242], x[241], x[240], x[248], x[247], x[246], x[239], x[238], x[237], x[254], x[253]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[270], x[269]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[262], x[261], x[260], x[265], x[264], x[263], x[268], x[267], x[266], x[272], x[271]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[265], x[264], x[263], x[262], x[261], x[260], x[268], x[267], x[266], x[259], x[258], x[257], x[274], x[273]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[290], x[289]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[282], x[281], x[280], x[285], x[284], x[283], x[288], x[287], x[286], x[292], x[291]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[285], x[284], x[283], x[282], x[281], x[280], x[288], x[287], x[286], x[279], x[278], x[277], x[294], x[293]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[310], x[309]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[302], x[301], x[300], x[305], x[304], x[303], x[308], x[307], x[306], x[312], x[311]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[305], x[304], x[303], x[302], x[301], x[300], x[308], x[307], x[306], x[299], x[298], x[297], x[314], x[313]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[330], x[329]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[322], x[321], x[320], x[325], x[324], x[323], x[328], x[327], x[326], x[332], x[331]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[325], x[324], x[323], x[322], x[321], x[320], x[328], x[327], x[326], x[319], x[318], x[317], x[334], x[333]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[350], x[349]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[342], x[341], x[340], x[345], x[344], x[343], x[348], x[347], x[346], x[352], x[351]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[345], x[344], x[343], x[342], x[341], x[340], x[348], x[347], x[346], x[339], x[338], x[337], x[354], x[353]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[368], x[367], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[355]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[368], x[367], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[357], x[370], x[369]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[362], x[361], x[360], x[365], x[364], x[363], x[368], x[367], x[366], x[372], x[371]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[365], x[364], x[363], x[362], x[361], x[360], x[368], x[367], x[366], x[359], x[358], x[357], x[374], x[373]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[375]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[390], x[389]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[382], x[381], x[380], x[385], x[384], x[383], x[388], x[387], x[386], x[392], x[391]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[385], x[384], x[383], x[382], x[381], x[380], x[388], x[387], x[386], x[379], x[378], x[377], x[394], x[393]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[410], x[409]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[402], x[401], x[400], x[405], x[404], x[403], x[408], x[407], x[406], x[412], x[411]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[405], x[404], x[403], x[402], x[401], x[400], x[408], x[407], x[406], x[399], x[398], x[397], x[414], x[413]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[430], x[429]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[422], x[421], x[420], x[425], x[424], x[423], x[428], x[427], x[426], x[432], x[431]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[425], x[424], x[423], x[422], x[421], x[420], x[428], x[427], x[426], x[419], x[418], x[417], x[434], x[433]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[450], x[449]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[442], x[441], x[440], x[445], x[444], x[443], x[448], x[447], x[446], x[452], x[451]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[448], x[447], x[446], x[439], x[438], x[437], x[454], x[453]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[468], x[467], x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[456], x[455]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[468], x[467], x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[470], x[469]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[462], x[461], x[460], x[465], x[464], x[463], x[468], x[467], x[466], x[472], x[471]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[465], x[464], x[463], x[462], x[461], x[460], x[468], x[467], x[466], x[459], x[458], x[457], x[474], x[473]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[476], x[475]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[490], x[489]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[482], x[481], x[480], x[485], x[484], x[483], x[488], x[487], x[486], x[492], x[491]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[485], x[484], x[483], x[482], x[481], x[480], x[488], x[487], x[486], x[479], x[478], x[477], x[494], x[493]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[508], x[507], x[506], x[505], x[504], x[503], x[502], x[501], x[500], x[499], x[498], x[497], x[496], x[495]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[508], x[507], x[506], x[505], x[504], x[503], x[502], x[501], x[500], x[499], x[498], x[497], x[510], x[509]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[502], x[501], x[500], x[505], x[504], x[503], x[508], x[507], x[506], x[512], x[511]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[505], x[504], x[503], x[502], x[501], x[500], x[508], x[507], x[506], x[499], x[498], x[497], x[514], x[513]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[248], x[247], x[246], x[268], x[267], x[266], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[228], x[227], x[226], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[236], x[235], x[299], x[298], x[297], x[256], x[255], x[499], x[498], x[497], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[216], x[215], x[399], x[398], x[397], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[196], x[195], x[529], x[528], x[527], x[202], x[201], x[200]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[248], x[247], x[246], x[268], x[267], x[266], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[228], x[227], x[226], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[250], x[249], x[299], x[298], x[297], x[270], x[269], x[499], x[498], x[497], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[230], x[229], x[399], x[398], x[397], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[210], x[209], x[530], x[528], x[527], x[208], x[207], x[206]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[242], x[241], x[240], x[262], x[261], x[260], x[245], x[244], x[243], x[248], x[247], x[246], x[302], x[301], x[300], x[265], x[264], x[263], x[268], x[267], x[266], x[502], x[501], x[500], x[222], x[221], x[220], x[252], x[251], x[305], x[304], x[303], x[308], x[307], x[306], x[272], x[271], x[505], x[504], x[503], x[508], x[507], x[506], x[225], x[224], x[223], x[228], x[227], x[226], x[402], x[401], x[400], x[232], x[231], x[405], x[404], x[403], x[408], x[407], x[406], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[212], x[211], x[531], x[528], x[527], x[199], x[198], x[197]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[265], x[264], x[263], x[245], x[244], x[243], x[262], x[261], x[260], x[268], x[267], x[266], x[505], x[504], x[503], x[242], x[241], x[240], x[248], x[247], x[246], x[305], x[304], x[303], x[225], x[224], x[223], x[274], x[273], x[259], x[258], x[257], x[502], x[501], x[500], x[508], x[507], x[506], x[254], x[253], x[239], x[238], x[237], x[302], x[301], x[300], x[308], x[307], x[306], x[222], x[221], x[220], x[228], x[227], x[226], x[405], x[404], x[403], x[499], x[498], x[497], x[299], x[298], x[297], x[234], x[233], x[219], x[218], x[217], x[402], x[401], x[400], x[408], x[407], x[406], x[399], x[398], x[397], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[214], x[213], x[532], x[528], x[527], x[205], x[204], x[203]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[248], x[247], x[246], x[268], x[267], x[266], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[288], x[287], x[286], x[488], x[487], x[486], x[328], x[327], x[326], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[208], x[207], x[206], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[236], x[235], x[299], x[298], x[297], x[256], x[255], x[499], x[498], x[497], x[205], x[204], x[203], x[202], x[201], x[200], x[296], x[295], x[279], x[278], x[277], x[276], x[275], x[479], x[478], x[477], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[196], x[195], x[199], x[198], x[197], x[316], x[315], x[419], x[418], x[417], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[216], x[215], x[533], x[528], x[527], x[222], x[221], x[220]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[248], x[247], x[246], x[268], x[267], x[266], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[288], x[287], x[286], x[488], x[487], x[486], x[328], x[327], x[326], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[208], x[207], x[206], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[250], x[249], x[299], x[298], x[297], x[270], x[269], x[499], x[498], x[497], x[205], x[204], x[203], x[202], x[201], x[200], x[310], x[309], x[279], x[278], x[277], x[290], x[289], x[479], x[478], x[477], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[210], x[209], x[199], x[198], x[197], x[330], x[329], x[419], x[418], x[417], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[230], x[229], x[534], x[528], x[527], x[228], x[227], x[226]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[242], x[241], x[240], x[262], x[261], x[260], x[245], x[244], x[243], x[248], x[247], x[246], x[302], x[301], x[300], x[265], x[264], x[263], x[268], x[267], x[266], x[502], x[501], x[500], x[482], x[481], x[480], x[282], x[281], x[280], x[322], x[321], x[320], x[252], x[251], x[305], x[304], x[303], x[308], x[307], x[306], x[272], x[271], x[505], x[504], x[503], x[508], x[507], x[506], x[202], x[201], x[200], x[292], x[291], x[485], x[484], x[483], x[488], x[487], x[486], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[325], x[324], x[323], x[328], x[327], x[326], x[422], x[421], x[420], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[332], x[331], x[425], x[424], x[423], x[428], x[427], x[426], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[232], x[231], x[535], x[528], x[527], x[219], x[218], x[217]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[265], x[264], x[263], x[245], x[244], x[243], x[262], x[261], x[260], x[268], x[267], x[266], x[505], x[504], x[503], x[242], x[241], x[240], x[248], x[247], x[246], x[305], x[304], x[303], x[285], x[284], x[283], x[485], x[484], x[483], x[325], x[324], x[323], x[274], x[273], x[259], x[258], x[257], x[502], x[501], x[500], x[508], x[507], x[506], x[254], x[253], x[239], x[238], x[237], x[302], x[301], x[300], x[308], x[307], x[306], x[205], x[204], x[203], x[314], x[313], x[282], x[281], x[280], x[288], x[287], x[286], x[294], x[293], x[482], x[481], x[480], x[488], x[487], x[486], x[322], x[321], x[320], x[328], x[327], x[326], x[425], x[424], x[423], x[499], x[498], x[497], x[299], x[298], x[297], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[279], x[278], x[277], x[479], x[478], x[477], x[334], x[333], x[319], x[318], x[317], x[422], x[421], x[420], x[428], x[427], x[426], x[199], x[198], x[197], x[419], x[418], x[417], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[234], x[233], x[536], x[528], x[527], x[225], x[224], x[223]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[228], x[227], x[226], x[448], x[447], x[446], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[268], x[267], x[266], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[368], x[367], x[366], x[216], x[215], x[399], x[398], x[397], x[196], x[195], x[199], x[198], x[197], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[455], x[456], x[459], x[458], x[457], x[435], x[436], x[339], x[338], x[337], x[365], x[364], x[363], x[362], x[361], x[360], x[256], x[255], x[499], x[498], x[497], x[495], x[496], x[359], x[358], x[357], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[236], x[235], x[537], x[528], x[527], x[242], x[241], x[240]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[228], x[227], x[226], x[448], x[447], x[446], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[268], x[267], x[266], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[368], x[367], x[366], x[230], x[229], x[399], x[398], x[397], x[210], x[209], x[199], x[198], x[197], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[469], x[470], x[459], x[458], x[457], x[449], x[450], x[339], x[338], x[337], x[365], x[364], x[363], x[362], x[361], x[360], x[270], x[269], x[499], x[498], x[497], x[509], x[510], x[359], x[358], x[357], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[250], x[249], x[538], x[528], x[527], x[248], x[247], x[246]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[222], x[221], x[220], x[442], x[441], x[440], x[202], x[201], x[200], x[225], x[224], x[223], x[228], x[227], x[226], x[402], x[401], x[400], x[262], x[261], x[260], x[445], x[444], x[443], x[448], x[447], x[446], x[342], x[341], x[340], x[462], x[461], x[460], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[232], x[231], x[405], x[404], x[403], x[408], x[407], x[406], x[265], x[264], x[263], x[268], x[267], x[266], x[502], x[501], x[500], x[451], x[452], x[345], x[344], x[343], x[348], x[347], x[346], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[362], x[361], x[360], x[272], x[271], x[505], x[504], x[503], x[508], x[507], x[506], x[511], x[512], x[365], x[364], x[363], x[368], x[367], x[366], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[252], x[251], x[539], x[528], x[527], x[239], x[238], x[237]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[225], x[224], x[223], x[445], x[444], x[443], x[222], x[221], x[220], x[228], x[227], x[226], x[405], x[404], x[403], x[205], x[204], x[203], x[265], x[264], x[263], x[465], x[464], x[463], x[442], x[441], x[440], x[448], x[447], x[446], x[345], x[344], x[343], x[234], x[233], x[219], x[218], x[217], x[402], x[401], x[400], x[408], x[407], x[406], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[262], x[261], x[260], x[268], x[267], x[266], x[505], x[504], x[503], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[453], x[454], x[439], x[438], x[437], x[342], x[341], x[340], x[348], x[347], x[346], x[365], x[364], x[363], x[399], x[398], x[397], x[199], x[198], x[197], x[274], x[273], x[259], x[258], x[257], x[502], x[501], x[500], x[508], x[507], x[506], x[459], x[458], x[457], x[339], x[338], x[337], x[513], x[514], x[362], x[361], x[360], x[368], x[367], x[366], x[499], x[498], x[497], x[359], x[358], x[357], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[254], x[253], x[540], x[528], x[527], x[245], x[244], x[243]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[228], x[227], x[226], x[428], x[427], x[426], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[248], x[247], x[246], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[368], x[367], x[366], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[216], x[215], x[399], x[398], x[397], x[196], x[195], x[199], x[198], x[197], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[395], x[396], x[439], x[438], x[437], x[415], x[416], x[319], x[318], x[317], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[236], x[235], x[299], x[298], x[297], x[355], x[356], x[379], x[378], x[377], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[256], x[255], x[541], x[528], x[527], x[262], x[261], x[260]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[228], x[227], x[226], x[428], x[427], x[426], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[248], x[247], x[246], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[368], x[367], x[366], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[230], x[229], x[399], x[398], x[397], x[210], x[209], x[199], x[198], x[197], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[409], x[410], x[439], x[438], x[437], x[429], x[430], x[319], x[318], x[317], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[250], x[249], x[299], x[298], x[297], x[369], x[370], x[379], x[378], x[377], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[270], x[269], x[542], x[528], x[527], x[268], x[267], x[266]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[222], x[221], x[220], x[422], x[421], x[420], x[202], x[201], x[200], x[225], x[224], x[223], x[228], x[227], x[226], x[402], x[401], x[400], x[242], x[241], x[240], x[442], x[441], x[440], x[425], x[424], x[423], x[428], x[427], x[426], x[322], x[321], x[320], x[362], x[361], x[360], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[232], x[231], x[405], x[404], x[403], x[408], x[407], x[406], x[245], x[244], x[243], x[248], x[247], x[246], x[302], x[301], x[300], x[411], x[412], x[445], x[444], x[443], x[448], x[447], x[446], x[431], x[432], x[325], x[324], x[323], x[328], x[327], x[326], x[365], x[364], x[363], x[368], x[367], x[366], x[382], x[381], x[380], x[252], x[251], x[305], x[304], x[303], x[308], x[307], x[306], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[272], x[271], x[543], x[528], x[527], x[259], x[258], x[257]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[225], x[224], x[223], x[425], x[424], x[423], x[222], x[221], x[220], x[228], x[227], x[226], x[405], x[404], x[403], x[205], x[204], x[203], x[245], x[244], x[243], x[422], x[421], x[420], x[428], x[427], x[426], x[325], x[324], x[323], x[445], x[444], x[443], x[365], x[364], x[363], x[234], x[233], x[219], x[218], x[217], x[402], x[401], x[400], x[408], x[407], x[406], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[242], x[241], x[240], x[248], x[247], x[246], x[305], x[304], x[303], x[433], x[434], x[419], x[418], x[417], x[322], x[321], x[320], x[328], x[327], x[326], x[413], x[414], x[442], x[441], x[440], x[448], x[447], x[446], x[362], x[361], x[360], x[368], x[367], x[366], x[385], x[384], x[383], x[399], x[398], x[397], x[199], x[198], x[197], x[254], x[253], x[239], x[238], x[237], x[302], x[301], x[300], x[308], x[307], x[306], x[319], x[318], x[317], x[439], x[438], x[437], x[373], x[374], x[359], x[358], x[357], x[382], x[381], x[380], x[388], x[387], x[386], x[299], x[298], x[297], x[379], x[378], x[377], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[274], x[273], x[544], x[528], x[527], x[265], x[264], x[263]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[328], x[327], x[326], x[348], x[347], x[346], x[308], x[307], x[306], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[488], x[487], x[486], x[299], x[298], x[297], x[285], x[284], x[283], x[316], x[315], x[419], x[418], x[417], x[335], x[336], x[219], x[218], x[217], x[485], x[484], x[483], x[482], x[481], x[480], x[296], x[295], x[279], x[278], x[277], x[479], x[478], x[477], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[276], x[275], x[545], x[528], x[527], x[282], x[281], x[280]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[328], x[327], x[326], x[348], x[347], x[346], x[308], x[307], x[306], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[305], x[304], x[303], x[302], x[301], x[300], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[488], x[487], x[486], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[330], x[329], x[419], x[418], x[417], x[349], x[350], x[219], x[218], x[217], x[485], x[484], x[483], x[482], x[481], x[480], x[310], x[309], x[279], x[278], x[277], x[479], x[478], x[477], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[290], x[289], x[546], x[528], x[527], x[288], x[287], x[286]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[322], x[321], x[320], x[342], x[341], x[340], x[302], x[301], x[300], x[325], x[324], x[323], x[328], x[327], x[326], x[422], x[421], x[420], x[345], x[344], x[343], x[348], x[347], x[346], x[222], x[221], x[220], x[305], x[304], x[303], x[308], x[307], x[306], x[282], x[281], x[280], x[332], x[331], x[425], x[424], x[423], x[428], x[427], x[426], x[351], x[352], x[225], x[224], x[223], x[228], x[227], x[226], x[482], x[481], x[480], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[485], x[484], x[483], x[488], x[487], x[486], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[292], x[291], x[547], x[528], x[527], x[279], x[278], x[277]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[345], x[344], x[343], x[325], x[324], x[323], x[305], x[304], x[303], x[342], x[341], x[340], x[348], x[347], x[346], x[225], x[224], x[223], x[322], x[321], x[320], x[328], x[327], x[326], x[425], x[424], x[423], x[302], x[301], x[300], x[308], x[307], x[306], x[353], x[354], x[339], x[338], x[337], x[222], x[221], x[220], x[228], x[227], x[226], x[334], x[333], x[319], x[318], x[317], x[422], x[421], x[420], x[428], x[427], x[426], x[485], x[484], x[483], x[314], x[313], x[299], x[298], x[297], x[282], x[281], x[280], x[288], x[287], x[286], x[219], x[218], x[217], x[419], x[418], x[417], x[482], x[481], x[480], x[488], x[487], x[486], x[279], x[278], x[277], x[479], x[478], x[477], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[294], x[293], x[548], x[528], x[527], x[285], x[284], x[283]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[328], x[327], x[326], x[348], x[347], x[346], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[288], x[287], x[286], x[408], x[407], x[406], x[208], x[207], x[206], x[268], x[267], x[266], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[285], x[284], x[283], x[282], x[281], x[280], x[488], x[487], x[486], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[316], x[315], x[419], x[418], x[417], x[335], x[336], x[219], x[218], x[217], x[279], x[278], x[277], x[485], x[484], x[483], x[482], x[481], x[480], x[216], x[215], x[399], x[398], x[397], x[196], x[195], x[199], x[198], x[197], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[276], x[275], x[479], x[478], x[477], x[256], x[255], x[499], x[498], x[497], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[296], x[295], x[549], x[528], x[527], x[302], x[301], x[300]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[328], x[327], x[326], x[348], x[347], x[346], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[288], x[287], x[286], x[408], x[407], x[406], x[208], x[207], x[206], x[268], x[267], x[266], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[285], x[284], x[283], x[282], x[281], x[280], x[488], x[487], x[486], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[265], x[264], x[263], x[262], x[261], x[260], x[508], x[507], x[506], x[330], x[329], x[419], x[418], x[417], x[349], x[350], x[219], x[218], x[217], x[279], x[278], x[277], x[485], x[484], x[483], x[482], x[481], x[480], x[230], x[229], x[399], x[398], x[397], x[210], x[209], x[199], x[198], x[197], x[259], x[258], x[257], x[505], x[504], x[503], x[502], x[501], x[500], x[290], x[289], x[479], x[478], x[477], x[270], x[269], x[499], x[498], x[497], x[310], x[309], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[550], x[528], x[527], x[308], x[307], x[306]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[322], x[321], x[320], x[342], x[341], x[340], x[325], x[324], x[323], x[328], x[327], x[326], x[422], x[421], x[420], x[345], x[344], x[343], x[348], x[347], x[346], x[222], x[221], x[220], x[282], x[281], x[280], x[202], x[201], x[200], x[402], x[401], x[400], x[262], x[261], x[260], x[332], x[331], x[425], x[424], x[423], x[428], x[427], x[426], x[351], x[352], x[225], x[224], x[223], x[228], x[227], x[226], x[285], x[284], x[283], x[288], x[287], x[286], x[482], x[481], x[480], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[232], x[231], x[405], x[404], x[403], x[408], x[407], x[406], x[265], x[264], x[263], x[268], x[267], x[266], x[502], x[501], x[500], x[292], x[291], x[485], x[484], x[483], x[488], x[487], x[486], x[272], x[271], x[505], x[504], x[503], x[508], x[507], x[506], x[312], x[311], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[551], x[528], x[527], x[299], x[298], x[297]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[345], x[344], x[343], x[325], x[324], x[323], x[342], x[341], x[340], x[348], x[347], x[346], x[225], x[224], x[223], x[322], x[321], x[320], x[328], x[327], x[326], x[425], x[424], x[423], x[285], x[284], x[283], x[405], x[404], x[403], x[205], x[204], x[203], x[265], x[264], x[263], x[353], x[354], x[339], x[338], x[337], x[222], x[221], x[220], x[228], x[227], x[226], x[334], x[333], x[319], x[318], x[317], x[422], x[421], x[420], x[428], x[427], x[426], x[282], x[281], x[280], x[288], x[287], x[286], x[485], x[484], x[483], x[234], x[233], x[402], x[401], x[400], x[408], x[407], x[406], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[262], x[261], x[260], x[268], x[267], x[266], x[505], x[504], x[503], x[219], x[218], x[217], x[419], x[418], x[417], x[294], x[293], x[279], x[278], x[277], x[482], x[481], x[480], x[488], x[487], x[486], x[399], x[398], x[397], x[199], x[198], x[197], x[274], x[273], x[259], x[258], x[257], x[502], x[501], x[500], x[508], x[507], x[506], x[479], x[478], x[477], x[499], x[498], x[497], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[314], x[313], x[552], x[528], x[527], x[305], x[304], x[303]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[308], x[307], x[306], x[368], x[367], x[366], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[348], x[347], x[346], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[408], x[407], x[406], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[296], x[295], x[279], x[278], x[277], x[276], x[275], x[479], x[478], x[477], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[375], x[376], x[259], x[258], x[257], x[355], x[356], x[379], x[378], x[377], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[335], x[336], x[219], x[218], x[217], x[395], x[396], x[439], x[438], x[437], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[316], x[315], x[553], x[528], x[527], x[322], x[321], x[320]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[308], x[307], x[306], x[368], x[367], x[366], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[348], x[347], x[346], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[408], x[407], x[406], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[310], x[309], x[279], x[278], x[277], x[290], x[289], x[479], x[478], x[477], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[389], x[390], x[259], x[258], x[257], x[369], x[370], x[379], x[378], x[377], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[349], x[350], x[219], x[218], x[217], x[409], x[410], x[439], x[438], x[437], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[330], x[329], x[554], x[528], x[527], x[328], x[327], x[326]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[302], x[301], x[300], x[362], x[361], x[360], x[482], x[481], x[480], x[305], x[304], x[303], x[308], x[307], x[306], x[282], x[281], x[280], x[342], x[341], x[340], x[365], x[364], x[363], x[368], x[367], x[366], x[382], x[381], x[380], x[262], x[261], x[260], x[402], x[401], x[400], x[292], x[291], x[485], x[484], x[483], x[488], x[487], x[486], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[345], x[344], x[343], x[348], x[347], x[346], x[222], x[221], x[220], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[391], x[392], x[265], x[264], x[263], x[268], x[267], x[266], x[405], x[404], x[403], x[408], x[407], x[406], x[442], x[441], x[440], x[351], x[352], x[225], x[224], x[223], x[228], x[227], x[226], x[411], x[412], x[445], x[444], x[443], x[448], x[447], x[446], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[332], x[331], x[555], x[528], x[527], x[319], x[318], x[317]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[305], x[304], x[303], x[365], x[364], x[363], x[302], x[301], x[300], x[308], x[307], x[306], x[285], x[284], x[283], x[485], x[484], x[483], x[345], x[344], x[343], x[265], x[264], x[263], x[362], x[361], x[360], x[368], x[367], x[366], x[385], x[384], x[383], x[405], x[404], x[403], x[314], x[313], x[299], x[298], x[297], x[282], x[281], x[280], x[288], x[287], x[286], x[294], x[293], x[482], x[481], x[480], x[488], x[487], x[486], x[342], x[341], x[340], x[348], x[347], x[346], x[225], x[224], x[223], x[393], x[394], x[262], x[261], x[260], x[268], x[267], x[266], x[373], x[374], x[359], x[358], x[357], x[382], x[381], x[380], x[388], x[387], x[386], x[402], x[401], x[400], x[408], x[407], x[406], x[445], x[444], x[443], x[279], x[278], x[277], x[479], x[478], x[477], x[353], x[354], x[339], x[338], x[337], x[222], x[221], x[220], x[228], x[227], x[226], x[259], x[258], x[257], x[379], x[378], x[377], x[413], x[414], x[399], x[398], x[397], x[442], x[441], x[440], x[448], x[447], x[446], x[219], x[218], x[217], x[439], x[438], x[437], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[334], x[333], x[556], x[528], x[527], x[325], x[324], x[323]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[308], x[307], x[306], x[508], x[507], x[506], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[328], x[327], x[326], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[468], x[467], x[466], x[296], x[295], x[279], x[278], x[277], x[276], x[275], x[479], x[478], x[477], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[476], x[475], x[239], x[238], x[237], x[495], x[496], x[359], x[358], x[357], x[465], x[464], x[463], x[462], x[461], x[460], x[316], x[315], x[419], x[418], x[417], x[455], x[456], x[459], x[458], x[457], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[336], x[335], x[557], x[528], x[527], x[342], x[341], x[340]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[308], x[307], x[306], x[508], x[507], x[506], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[328], x[327], x[326], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[468], x[467], x[466], x[310], x[309], x[279], x[278], x[277], x[290], x[289], x[479], x[478], x[477], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[489], x[490], x[239], x[238], x[237], x[509], x[510], x[359], x[358], x[357], x[465], x[464], x[463], x[462], x[461], x[460], x[330], x[329], x[419], x[418], x[417], x[469], x[470], x[459], x[458], x[457], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[350], x[349], x[558], x[528], x[527], x[348], x[347], x[346]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[302], x[301], x[300], x[502], x[501], x[500], x[482], x[481], x[480], x[305], x[304], x[303], x[308], x[307], x[306], x[282], x[281], x[280], x[322], x[321], x[320], x[242], x[241], x[240], x[505], x[504], x[503], x[508], x[507], x[506], x[362], x[361], x[360], x[292], x[291], x[485], x[484], x[483], x[488], x[487], x[486], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[325], x[324], x[323], x[328], x[327], x[326], x[422], x[421], x[420], x[491], x[492], x[245], x[244], x[243], x[248], x[247], x[246], x[511], x[512], x[365], x[364], x[363], x[368], x[367], x[366], x[462], x[461], x[460], x[332], x[331], x[425], x[424], x[423], x[428], x[427], x[426], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[352], x[351], x[559], x[528], x[527], x[339], x[338], x[337]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[305], x[304], x[303], x[505], x[504], x[503], x[302], x[301], x[300], x[308], x[307], x[306], x[285], x[284], x[283], x[485], x[484], x[483], x[325], x[324], x[323], x[502], x[501], x[500], x[508], x[507], x[506], x[365], x[364], x[363], x[245], x[244], x[243], x[314], x[313], x[299], x[298], x[297], x[282], x[281], x[280], x[288], x[287], x[286], x[294], x[293], x[482], x[481], x[480], x[488], x[487], x[486], x[322], x[321], x[320], x[328], x[327], x[326], x[425], x[424], x[423], x[513], x[514], x[499], x[498], x[497], x[362], x[361], x[360], x[368], x[367], x[366], x[493], x[494], x[242], x[241], x[240], x[248], x[247], x[246], x[465], x[464], x[463], x[279], x[278], x[277], x[479], x[478], x[477], x[334], x[333], x[319], x[318], x[317], x[422], x[421], x[420], x[428], x[427], x[426], x[359], x[358], x[357], x[239], x[238], x[237], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[419], x[418], x[417], x[459], x[458], x[457], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[354], x[353], x[560], x[528], x[527], x[345], x[344], x[343]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[408], x[407], x[406], x[428], x[427], x[426], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[388], x[387], x[386], x[468], x[467], x[466], x[348], x[347], x[346], x[488], x[487], x[486], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[385], x[384], x[383], x[382], x[381], x[380], x[268], x[267], x[266], x[465], x[464], x[463], x[462], x[461], x[460], x[345], x[344], x[343], x[342], x[341], x[340], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[395], x[396], x[439], x[438], x[437], x[415], x[416], x[319], x[318], x[317], x[379], x[378], x[377], x[265], x[264], x[263], x[262], x[261], x[260], x[455], x[456], x[459], x[458], x[457], x[435], x[436], x[339], x[338], x[337], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[375], x[376], x[259], x[258], x[257], x[476], x[475], x[239], x[238], x[237], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[356], x[355], x[561], x[528], x[527], x[362], x[361], x[360]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[408], x[407], x[406], x[428], x[427], x[426], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[388], x[387], x[386], x[468], x[467], x[466], x[348], x[347], x[346], x[488], x[487], x[486], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[385], x[384], x[383], x[382], x[381], x[380], x[268], x[267], x[266], x[465], x[464], x[463], x[462], x[461], x[460], x[345], x[344], x[343], x[342], x[341], x[340], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[409], x[410], x[439], x[438], x[437], x[429], x[430], x[319], x[318], x[317], x[379], x[378], x[377], x[265], x[264], x[263], x[262], x[261], x[260], x[469], x[470], x[459], x[458], x[457], x[449], x[450], x[339], x[338], x[337], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[389], x[390], x[259], x[258], x[257], x[489], x[490], x[239], x[238], x[237], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[370], x[369], x[562], x[528], x[527], x[368], x[367], x[366]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[402], x[401], x[400], x[422], x[421], x[420], x[405], x[404], x[403], x[408], x[407], x[406], x[442], x[441], x[440], x[425], x[424], x[423], x[428], x[427], x[426], x[322], x[321], x[320], x[382], x[381], x[380], x[342], x[341], x[340], x[462], x[461], x[460], x[482], x[481], x[480], x[411], x[412], x[445], x[444], x[443], x[448], x[447], x[446], x[431], x[432], x[325], x[324], x[323], x[328], x[327], x[326], x[385], x[384], x[383], x[388], x[387], x[386], x[262], x[261], x[260], x[451], x[452], x[345], x[344], x[343], x[348], x[347], x[346], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[485], x[484], x[483], x[488], x[487], x[486], x[242], x[241], x[240], x[391], x[392], x[265], x[264], x[263], x[268], x[267], x[266], x[491], x[492], x[245], x[244], x[243], x[248], x[247], x[246], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[372], x[371], x[563], x[528], x[527], x[359], x[358], x[357]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[425], x[424], x[423], x[405], x[404], x[403], x[422], x[421], x[420], x[428], x[427], x[426], x[325], x[324], x[323], x[402], x[401], x[400], x[408], x[407], x[406], x[445], x[444], x[443], x[385], x[384], x[383], x[465], x[464], x[463], x[345], x[344], x[343], x[485], x[484], x[483], x[433], x[434], x[419], x[418], x[417], x[322], x[321], x[320], x[328], x[327], x[326], x[413], x[414], x[399], x[398], x[397], x[442], x[441], x[440], x[448], x[447], x[446], x[382], x[381], x[380], x[388], x[387], x[386], x[265], x[264], x[263], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[453], x[454], x[342], x[341], x[340], x[348], x[347], x[346], x[482], x[481], x[480], x[488], x[487], x[486], x[245], x[244], x[243], x[319], x[318], x[317], x[439], x[438], x[437], x[393], x[394], x[379], x[378], x[377], x[262], x[261], x[260], x[268], x[267], x[266], x[459], x[458], x[457], x[339], x[338], x[337], x[493], x[494], x[479], x[478], x[477], x[242], x[241], x[240], x[248], x[247], x[246], x[259], x[258], x[257], x[239], x[238], x[237], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[374], x[373], x[564], x[528], x[527], x[365], x[364], x[363]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[408], x[407], x[406], x[428], x[427], x[426], x[368], x[367], x[366], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[268], x[267], x[266], x[359], x[358], x[357], x[385], x[384], x[383], x[395], x[396], x[439], x[438], x[437], x[415], x[416], x[319], x[318], x[317], x[265], x[264], x[263], x[262], x[261], x[260], x[355], x[356], x[379], x[378], x[377], x[259], x[258], x[257], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[376], x[375], x[565], x[528], x[527], x[382], x[381], x[380]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[408], x[407], x[406], x[428], x[427], x[426], x[368], x[367], x[366], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[365], x[364], x[363], x[362], x[361], x[360], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[268], x[267], x[266], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[409], x[410], x[439], x[438], x[437], x[429], x[430], x[319], x[318], x[317], x[265], x[264], x[263], x[262], x[261], x[260], x[369], x[370], x[379], x[378], x[377], x[259], x[258], x[257], x[526], x[525], x[524], x[520], x[519], x[518], x[517], x[516], x[515], x[523], x[522], x[521], x[390], x[389], x[566], x[528], x[527], x[388], x[387], x[386]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[402], x[401], x[400], x[422], x[421], x[420], x[362], x[361], x[360], x[405], x[404], x[403], x[408], x[407], x[406], x[442], x[441], x[440], x[425], x[424], x[423], x[428], x[427], x[426], x[322], x[321], x[320], x[365], x[364], x[363], x[368], x[367], x[366], x[382], x[381], x[380], x[411], x[412], x[445], x[444], x[443], x[448], x[447], x[446], x[431], x[432], x[325], x[324], x[323], x[328], x[327], x[326], x[262], x[261], x[260], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[265], x[264], x[263], x[268], x[267], x[266], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[392], x[391], x[567], x[528], x[527], x[379], x[378], x[377]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[425], x[424], x[423], x[405], x[404], x[403], x[365], x[364], x[363], x[422], x[421], x[420], x[428], x[427], x[426], x[325], x[324], x[323], x[402], x[401], x[400], x[408], x[407], x[406], x[445], x[444], x[443], x[362], x[361], x[360], x[368], x[367], x[366], x[433], x[434], x[419], x[418], x[417], x[322], x[321], x[320], x[328], x[327], x[326], x[413], x[414], x[399], x[398], x[397], x[442], x[441], x[440], x[448], x[447], x[446], x[265], x[264], x[263], x[373], x[374], x[359], x[358], x[357], x[382], x[381], x[380], x[388], x[387], x[386], x[319], x[318], x[317], x[439], x[438], x[437], x[262], x[261], x[260], x[268], x[267], x[266], x[379], x[378], x[377], x[259], x[258], x[257], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[394], x[393], x[568], x[528], x[527], x[385], x[384], x[383]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[368], x[367], x[366], x[248], x[247], x[246], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[428], x[427], x[426], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[508], x[507], x[506], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[505], x[504], x[503], x[502], x[501], x[500], x[208], x[207], x[206], x[375], x[376], x[259], x[258], x[257], x[355], x[356], x[379], x[378], x[377], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[236], x[235], x[299], x[298], x[297], x[256], x[255], x[499], x[498], x[497], x[205], x[204], x[203], x[202], x[201], x[200], x[415], x[416], x[319], x[318], x[317], x[196], x[195], x[199], x[198], x[197], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[396], x[395], x[569], x[528], x[527], x[402], x[401], x[400]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[368], x[367], x[366], x[248], x[247], x[246], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[428], x[427], x[426], x[245], x[244], x[243], x[242], x[241], x[240], x[308], x[307], x[306], x[508], x[507], x[506], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[239], x[238], x[237], x[305], x[304], x[303], x[302], x[301], x[300], x[505], x[504], x[503], x[502], x[501], x[500], x[208], x[207], x[206], x[389], x[390], x[259], x[258], x[257], x[369], x[370], x[379], x[378], x[377], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[250], x[249], x[299], x[298], x[297], x[270], x[269], x[499], x[498], x[497], x[205], x[204], x[203], x[202], x[201], x[200], x[429], x[430], x[319], x[318], x[317], x[210], x[209], x[199], x[198], x[197], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[410], x[409], x[570], x[528], x[527], x[408], x[407], x[406]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[362], x[361], x[360], x[242], x[241], x[240], x[365], x[364], x[363], x[368], x[367], x[366], x[382], x[381], x[380], x[262], x[261], x[260], x[422], x[421], x[420], x[245], x[244], x[243], x[248], x[247], x[246], x[302], x[301], x[300], x[502], x[501], x[500], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[391], x[392], x[265], x[264], x[263], x[268], x[267], x[266], x[425], x[424], x[423], x[428], x[427], x[426], x[322], x[321], x[320], x[252], x[251], x[305], x[304], x[303], x[308], x[307], x[306], x[272], x[271], x[505], x[504], x[503], x[508], x[507], x[506], x[202], x[201], x[200], x[431], x[432], x[325], x[324], x[323], x[328], x[327], x[326], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[412], x[411], x[571], x[528], x[527], x[399], x[398], x[397]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[365], x[364], x[363], x[245], x[244], x[243], x[265], x[264], x[263], x[362], x[361], x[360], x[368], x[367], x[366], x[385], x[384], x[383], x[425], x[424], x[423], x[505], x[504], x[503], x[242], x[241], x[240], x[248], x[247], x[246], x[305], x[304], x[303], x[393], x[394], x[262], x[261], x[260], x[268], x[267], x[266], x[373], x[374], x[359], x[358], x[357], x[382], x[381], x[380], x[388], x[387], x[386], x[422], x[421], x[420], x[428], x[427], x[426], x[325], x[324], x[323], x[274], x[273], x[502], x[501], x[500], x[508], x[507], x[506], x[254], x[253], x[239], x[238], x[237], x[302], x[301], x[300], x[308], x[307], x[306], x[205], x[204], x[203], x[259], x[258], x[257], x[379], x[378], x[377], x[433], x[434], x[419], x[418], x[417], x[322], x[321], x[320], x[328], x[327], x[326], x[499], x[498], x[497], x[299], x[298], x[297], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[319], x[318], x[317], x[199], x[198], x[197], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[414], x[413], x[572], x[528], x[527], x[405], x[404], x[403]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[368], x[367], x[366], x[308], x[307], x[306], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[408], x[407], x[406], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[348], x[347], x[346], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[375], x[376], x[259], x[258], x[257], x[355], x[356], x[379], x[378], x[377], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[296], x[295], x[279], x[278], x[277], x[276], x[275], x[479], x[478], x[477], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[395], x[396], x[439], x[438], x[437], x[335], x[336], x[219], x[218], x[217], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[416], x[415], x[573], x[528], x[527], x[422], x[421], x[420]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[368], x[367], x[366], x[308], x[307], x[306], x[268], x[267], x[266], x[365], x[364], x[363], x[362], x[361], x[360], x[388], x[387], x[386], x[408], x[407], x[406], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[488], x[487], x[486], x[348], x[347], x[346], x[265], x[264], x[263], x[262], x[261], x[260], x[359], x[358], x[357], x[385], x[384], x[383], x[382], x[381], x[380], x[405], x[404], x[403], x[402], x[401], x[400], x[448], x[447], x[446], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[485], x[484], x[483], x[482], x[481], x[480], x[345], x[344], x[343], x[342], x[341], x[340], x[228], x[227], x[226], x[389], x[390], x[259], x[258], x[257], x[369], x[370], x[379], x[378], x[377], x[399], x[398], x[397], x[445], x[444], x[443], x[442], x[441], x[440], x[310], x[309], x[279], x[278], x[277], x[290], x[289], x[479], x[478], x[477], x[339], x[338], x[337], x[225], x[224], x[223], x[222], x[221], x[220], x[409], x[410], x[439], x[438], x[437], x[349], x[350], x[219], x[218], x[217], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[430], x[429], x[574], x[528], x[527], x[428], x[427], x[426]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[362], x[361], x[360], x[302], x[301], x[300], x[365], x[364], x[363], x[368], x[367], x[366], x[382], x[381], x[380], x[262], x[261], x[260], x[402], x[401], x[400], x[482], x[481], x[480], x[305], x[304], x[303], x[308], x[307], x[306], x[282], x[281], x[280], x[342], x[341], x[340], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[391], x[392], x[265], x[264], x[263], x[268], x[267], x[266], x[405], x[404], x[403], x[408], x[407], x[406], x[442], x[441], x[440], x[292], x[291], x[485], x[484], x[483], x[488], x[487], x[486], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[345], x[344], x[343], x[348], x[347], x[346], x[222], x[221], x[220], x[411], x[412], x[445], x[444], x[443], x[448], x[447], x[446], x[351], x[352], x[225], x[224], x[223], x[228], x[227], x[226], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[432], x[431], x[575], x[528], x[527], x[419], x[418], x[417]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[365], x[364], x[363], x[305], x[304], x[303], x[265], x[264], x[263], x[362], x[361], x[360], x[368], x[367], x[366], x[385], x[384], x[383], x[405], x[404], x[403], x[302], x[301], x[300], x[308], x[307], x[306], x[285], x[284], x[283], x[485], x[484], x[483], x[345], x[344], x[343], x[393], x[394], x[262], x[261], x[260], x[268], x[267], x[266], x[373], x[374], x[359], x[358], x[357], x[382], x[381], x[380], x[388], x[387], x[386], x[402], x[401], x[400], x[408], x[407], x[406], x[445], x[444], x[443], x[314], x[313], x[299], x[298], x[297], x[282], x[281], x[280], x[288], x[287], x[286], x[294], x[293], x[482], x[481], x[480], x[488], x[487], x[486], x[342], x[341], x[340], x[348], x[347], x[346], x[225], x[224], x[223], x[259], x[258], x[257], x[379], x[378], x[377], x[413], x[414], x[399], x[398], x[397], x[442], x[441], x[440], x[448], x[447], x[446], x[279], x[278], x[277], x[479], x[478], x[477], x[353], x[354], x[339], x[338], x[337], x[222], x[221], x[220], x[228], x[227], x[226], x[439], x[438], x[437], x[219], x[218], x[217], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[434], x[433], x[576], x[528], x[527], x[425], x[424], x[423]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[488], x[487], x[486], x[508], x[507], x[506], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[268], x[267], x[266], x[388], x[387], x[386], x[428], x[427], x[426], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[468], x[467], x[466], x[265], x[264], x[263], x[262], x[261], x[260], x[385], x[384], x[383], x[382], x[381], x[380], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[476], x[475], x[239], x[238], x[237], x[495], x[496], x[359], x[358], x[357], x[465], x[464], x[463], x[462], x[461], x[460], x[375], x[376], x[259], x[258], x[257], x[355], x[356], x[379], x[378], x[377], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[455], x[456], x[459], x[458], x[457], x[415], x[416], x[319], x[318], x[317], x[436], x[435], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[577], x[528], x[527], x[442], x[441], x[440]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[488], x[487], x[486], x[508], x[507], x[506], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[268], x[267], x[266], x[388], x[387], x[386], x[428], x[427], x[426], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[468], x[467], x[466], x[265], x[264], x[263], x[262], x[261], x[260], x[385], x[384], x[383], x[382], x[381], x[380], x[425], x[424], x[423], x[422], x[421], x[420], x[328], x[327], x[326], x[489], x[490], x[239], x[238], x[237], x[509], x[510], x[359], x[358], x[357], x[465], x[464], x[463], x[462], x[461], x[460], x[389], x[390], x[259], x[258], x[257], x[369], x[370], x[379], x[378], x[377], x[419], x[418], x[417], x[325], x[324], x[323], x[322], x[321], x[320], x[469], x[470], x[459], x[458], x[457], x[429], x[430], x[319], x[318], x[317], x[450], x[449], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[578], x[528], x[527], x[448], x[447], x[446]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[482], x[481], x[480], x[502], x[501], x[500], x[485], x[484], x[483], x[488], x[487], x[486], x[242], x[241], x[240], x[505], x[504], x[503], x[508], x[507], x[506], x[362], x[361], x[360], x[382], x[381], x[380], x[262], x[261], x[260], x[422], x[421], x[420], x[491], x[492], x[245], x[244], x[243], x[248], x[247], x[246], x[511], x[512], x[365], x[364], x[363], x[368], x[367], x[366], x[462], x[461], x[460], x[371], x[372], x[385], x[384], x[383], x[388], x[387], x[386], x[391], x[392], x[265], x[264], x[263], x[268], x[267], x[266], x[425], x[424], x[423], x[428], x[427], x[426], x[322], x[321], x[320], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[431], x[432], x[325], x[324], x[323], x[328], x[327], x[326], x[452], x[451], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[579], x[528], x[527], x[439], x[438], x[437]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[505], x[504], x[503], x[485], x[484], x[483], x[502], x[501], x[500], x[508], x[507], x[506], x[365], x[364], x[363], x[482], x[481], x[480], x[488], x[487], x[486], x[245], x[244], x[243], x[265], x[264], x[263], x[385], x[384], x[383], x[425], x[424], x[423], x[513], x[514], x[499], x[498], x[497], x[362], x[361], x[360], x[368], x[367], x[366], x[493], x[494], x[479], x[478], x[477], x[242], x[241], x[240], x[248], x[247], x[246], x[465], x[464], x[463], x[393], x[394], x[262], x[261], x[260], x[268], x[267], x[266], x[373], x[374], x[382], x[381], x[380], x[388], x[387], x[386], x[422], x[421], x[420], x[428], x[427], x[426], x[325], x[324], x[323], x[359], x[358], x[357], x[239], x[238], x[237], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[259], x[258], x[257], x[379], x[378], x[377], x[433], x[434], x[419], x[418], x[417], x[322], x[321], x[320], x[328], x[327], x[326], x[459], x[458], x[457], x[319], x[318], x[317], x[454], x[453], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[580], x[528], x[527], x[445], x[444], x[443]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[488], x[487], x[486], x[508], x[507], x[506], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[448], x[447], x[446], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[476], x[475], x[239], x[238], x[237], x[495], x[496], x[359], x[358], x[357], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[435], x[436], x[339], x[338], x[337], x[456], x[455], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[581], x[528], x[527], x[462], x[461], x[460]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[488], x[487], x[486], x[508], x[507], x[506], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[448], x[447], x[446], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[489], x[490], x[239], x[238], x[237], x[509], x[510], x[359], x[358], x[357], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[449], x[450], x[339], x[338], x[337], x[470], x[469], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[582], x[528], x[527], x[468], x[467], x[466]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[482], x[481], x[480], x[502], x[501], x[500], x[485], x[484], x[483], x[488], x[487], x[486], x[242], x[241], x[240], x[505], x[504], x[503], x[508], x[507], x[506], x[362], x[361], x[360], x[442], x[441], x[440], x[491], x[492], x[245], x[244], x[243], x[248], x[247], x[246], x[511], x[512], x[365], x[364], x[363], x[368], x[367], x[366], x[445], x[444], x[443], x[448], x[447], x[446], x[342], x[341], x[340], x[451], x[452], x[345], x[344], x[343], x[348], x[347], x[346], x[472], x[471], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[583], x[528], x[527], x[459], x[458], x[457]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[505], x[504], x[503], x[485], x[484], x[483], x[502], x[501], x[500], x[508], x[507], x[506], x[365], x[364], x[363], x[482], x[481], x[480], x[488], x[487], x[486], x[245], x[244], x[243], x[445], x[444], x[443], x[513], x[514], x[499], x[498], x[497], x[362], x[361], x[360], x[368], x[367], x[366], x[493], x[494], x[479], x[478], x[477], x[242], x[241], x[240], x[248], x[247], x[246], x[442], x[441], x[440], x[448], x[447], x[446], x[345], x[344], x[343], x[359], x[358], x[357], x[239], x[238], x[237], x[453], x[454], x[439], x[438], x[437], x[342], x[341], x[340], x[348], x[347], x[346], x[339], x[338], x[337], x[474], x[473], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[584], x[528], x[527], x[465], x[464], x[463]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[448], x[447], x[446], x[328], x[327], x[326], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[508], x[507], x[506], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[228], x[227], x[226], x[308], x[307], x[306], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[225], x[224], x[223], x[222], x[221], x[220], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[455], x[456], x[459], x[458], x[457], x[435], x[436], x[339], x[338], x[337], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[316], x[315], x[419], x[418], x[417], x[335], x[336], x[219], x[218], x[217], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[495], x[496], x[359], x[358], x[357], x[296], x[295], x[279], x[278], x[277], x[476], x[475], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[585], x[528], x[527], x[482], x[481], x[480]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[448], x[447], x[446], x[328], x[327], x[326], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[508], x[507], x[506], x[325], x[324], x[323], x[322], x[321], x[320], x[428], x[427], x[426], x[228], x[227], x[226], x[308], x[307], x[306], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[505], x[504], x[503], x[502], x[501], x[500], x[368], x[367], x[366], x[319], x[318], x[317], x[425], x[424], x[423], x[422], x[421], x[420], x[225], x[224], x[223], x[222], x[221], x[220], x[305], x[304], x[303], x[302], x[301], x[300], x[288], x[287], x[286], x[469], x[470], x[459], x[458], x[457], x[449], x[450], x[339], x[338], x[337], x[499], x[498], x[497], x[365], x[364], x[363], x[362], x[361], x[360], x[330], x[329], x[419], x[418], x[417], x[349], x[350], x[219], x[218], x[217], x[299], x[298], x[297], x[285], x[284], x[283], x[282], x[281], x[280], x[509], x[510], x[359], x[358], x[357], x[310], x[309], x[279], x[278], x[277], x[490], x[489], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[586], x[528], x[527], x[488], x[487], x[486]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[442], x[441], x[440], x[322], x[321], x[320], x[445], x[444], x[443], x[448], x[447], x[446], x[342], x[341], x[340], x[462], x[461], x[460], x[502], x[501], x[500], x[325], x[324], x[323], x[328], x[327], x[326], x[422], x[421], x[420], x[222], x[221], x[220], x[302], x[301], x[300], x[451], x[452], x[345], x[344], x[343], x[348], x[347], x[346], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[505], x[504], x[503], x[508], x[507], x[506], x[362], x[361], x[360], x[332], x[331], x[425], x[424], x[423], x[428], x[427], x[426], x[351], x[352], x[225], x[224], x[223], x[228], x[227], x[226], x[305], x[304], x[303], x[308], x[307], x[306], x[282], x[281], x[280], x[511], x[512], x[365], x[364], x[363], x[368], x[367], x[366], x[312], x[311], x[285], x[284], x[283], x[288], x[287], x[286], x[492], x[491], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[587], x[528], x[527], x[479], x[478], x[477]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[445], x[444], x[443], x[325], x[324], x[323], x[465], x[464], x[463], x[442], x[441], x[440], x[448], x[447], x[446], x[345], x[344], x[343], x[505], x[504], x[503], x[225], x[224], x[223], x[322], x[321], x[320], x[328], x[327], x[326], x[425], x[424], x[423], x[305], x[304], x[303], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[453], x[454], x[439], x[438], x[437], x[342], x[341], x[340], x[348], x[347], x[346], x[502], x[501], x[500], x[508], x[507], x[506], x[365], x[364], x[363], x[353], x[354], x[222], x[221], x[220], x[228], x[227], x[226], x[334], x[333], x[319], x[318], x[317], x[422], x[421], x[420], x[428], x[427], x[426], x[302], x[301], x[300], x[308], x[307], x[306], x[285], x[284], x[283], x[459], x[458], x[457], x[339], x[338], x[337], x[513], x[514], x[499], x[498], x[497], x[362], x[361], x[360], x[368], x[367], x[366], x[219], x[218], x[217], x[419], x[418], x[417], x[314], x[313], x[299], x[298], x[297], x[282], x[281], x[280], x[288], x[287], x[286], x[359], x[358], x[357], x[279], x[278], x[277], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[494], x[493], x[588], x[528], x[527], x[485], x[484], x[483]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[448], x[447], x[446], x[228], x[227], x[226], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[488], x[487], x[486], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[308], x[307], x[306], x[455], x[456], x[459], x[458], x[457], x[435], x[436], x[339], x[338], x[337], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[216], x[215], x[399], x[398], x[397], x[196], x[195], x[199], x[198], x[197], x[305], x[304], x[303], x[302], x[301], x[300], x[476], x[475], x[239], x[238], x[237], x[236], x[235], x[299], x[298], x[297], x[496], x[495], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[589], x[528], x[527], x[502], x[501], x[500]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[448], x[447], x[446], x[228], x[227], x[226], x[468], x[467], x[466], x[445], x[444], x[443], x[442], x[441], x[440], x[348], x[347], x[346], x[488], x[487], x[486], x[225], x[224], x[223], x[222], x[221], x[220], x[408], x[407], x[406], x[208], x[207], x[206], x[465], x[464], x[463], x[462], x[461], x[460], x[439], x[438], x[437], x[345], x[344], x[343], x[342], x[341], x[340], x[485], x[484], x[483], x[482], x[481], x[480], x[248], x[247], x[246], x[219], x[218], x[217], x[405], x[404], x[403], x[402], x[401], x[400], x[205], x[204], x[203], x[202], x[201], x[200], x[308], x[307], x[306], x[469], x[470], x[459], x[458], x[457], x[449], x[450], x[339], x[338], x[337], x[479], x[478], x[477], x[245], x[244], x[243], x[242], x[241], x[240], x[230], x[229], x[399], x[398], x[397], x[210], x[209], x[199], x[198], x[197], x[305], x[304], x[303], x[302], x[301], x[300], x[489], x[490], x[239], x[238], x[237], x[250], x[249], x[299], x[298], x[297], x[526], x[525], x[524], x[520], x[519], x[518], x[517], x[516], x[515], x[523], x[522], x[521], x[510], x[509], x[590], x[528], x[527], x[508], x[507], x[506]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[442], x[441], x[440], x[222], x[221], x[220], x[445], x[444], x[443], x[448], x[447], x[446], x[342], x[341], x[340], x[462], x[461], x[460], x[482], x[481], x[480], x[202], x[201], x[200], x[225], x[224], x[223], x[228], x[227], x[226], x[402], x[401], x[400], x[451], x[452], x[345], x[344], x[343], x[348], x[347], x[346], x[472], x[471], x[465], x[464], x[463], x[468], x[467], x[466], x[485], x[484], x[483], x[488], x[487], x[486], x[242], x[241], x[240], x[212], x[211], x[205], x[204], x[203], x[208], x[207], x[206], x[232], x[231], x[405], x[404], x[403], x[408], x[407], x[406], x[302], x[301], x[300], x[491], x[492], x[245], x[244], x[243], x[248], x[247], x[246], x[252], x[251], x[305], x[304], x[303], x[308], x[307], x[306], x[512], x[511], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[591], x[528], x[527], x[499], x[498], x[497]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[445], x[444], x[443], x[225], x[224], x[223], x[465], x[464], x[463], x[442], x[441], x[440], x[448], x[447], x[446], x[345], x[344], x[343], x[485], x[484], x[483], x[222], x[221], x[220], x[228], x[227], x[226], x[405], x[404], x[403], x[205], x[204], x[203], x[474], x[473], x[462], x[461], x[460], x[468], x[467], x[466], x[453], x[454], x[439], x[438], x[437], x[342], x[341], x[340], x[348], x[347], x[346], x[482], x[481], x[480], x[488], x[487], x[486], x[245], x[244], x[243], x[234], x[233], x[219], x[218], x[217], x[402], x[401], x[400], x[408], x[407], x[406], x[214], x[213], x[202], x[201], x[200], x[208], x[207], x[206], x[305], x[304], x[303], x[459], x[458], x[457], x[339], x[338], x[337], x[493], x[494], x[479], x[478], x[477], x[242], x[241], x[240], x[248], x[247], x[246], x[399], x[398], x[397], x[199], x[198], x[197], x[254], x[253], x[302], x[301], x[300], x[308], x[307], x[306], x[239], x[238], x[237], x[299], x[298], x[297], x[526], x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[513], x[592], x[528], x[527], x[505], x[504], x[503]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[523], x[522], x[521], x[526], x[525], x[524], x[517], x[516], x[515], x[520], x[519], x[518], x[527]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[520], x[519], x[518], x[523], x[522], x[521], x[526], x[525], x[524], x[517], x[516], x[515], x[527]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[520], x[519], x[518], x[517], x[516], x[515], x[523], x[522], x[521], x[526], x[525], x[524], x[527]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[526], x[525], x[524], x[520], x[519], x[518], x[517], x[516], x[515], x[523], x[522], x[521], x[527]}), .y(y[197]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (t[15] & ~t[16]);
  assign t[12] = (t[17] & ~t[18]);
  assign t[13] = (t[19] & ~t[20]);
  assign t[14] = (t[21] & ~t[22]);
  assign t[15] = t[23] ^ x[2];
  assign t[16] = t[24] ^ x[1];
  assign t[17] = t[25] ^ x[5];
  assign t[18] = t[26] ^ x[4];
  assign t[19] = t[27] ^ x[8];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[7];
  assign t[21] = t[29] ^ x[11];
  assign t[22] = t[30] ^ x[10];
  assign t[23] = (x[0]);
  assign t[24] = (x[0]);
  assign t[25] = (x[3]);
  assign t[26] = (x[3]);
  assign t[27] = (x[6]);
  assign t[28] = (x[6]);
  assign t[29] = (x[9]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (t[15] & ~t[16]);
  assign t[12] = (t[17] & ~t[18]);
  assign t[13] = (t[19] & ~t[20]);
  assign t[14] = (t[21] & ~t[22]);
  assign t[15] = t[23] ^ x[2];
  assign t[16] = t[24] ^ x[1];
  assign t[17] = t[25] ^ x[5];
  assign t[18] = t[26] ^ x[4];
  assign t[19] = t[27] ^ x[8];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[7];
  assign t[21] = t[29] ^ x[11];
  assign t[22] = t[30] ^ x[10];
  assign t[23] = (x[0]);
  assign t[24] = (x[0]);
  assign t[25] = (x[3]);
  assign t[26] = (x[3]);
  assign t[27] = (x[6]);
  assign t[28] = (x[6]);
  assign t[29] = (x[9]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[2];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[11];
  assign t[31] = (x[1]);
  assign t[32] = (x[1]);
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[2];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[11];
  assign t[31] = (x[1]);
  assign t[32] = (x[1]);
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1]);
  assign t[31] = (x[1]);
  assign t[32] = (x[4]);
  assign t[33] = (x[4]);
  assign t[34] = (x[7]);
  assign t[35] = (x[7]);
  assign t[36] = (x[10]);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1]);
  assign t[31] = (x[1]);
  assign t[32] = (x[4]);
  assign t[33] = (x[4]);
  assign t[34] = (x[7]);
  assign t[35] = (x[7]);
  assign t[36] = (x[10]);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (t[20] & ~t[21]);
  assign t[17] = (t[22] & ~t[23]);
  assign t[18] = (t[24] & ~t[25]);
  assign t[19] = (t[26] & ~t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = t[35] ^ x[11];
  assign t[28] = (x[1]);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4]);
  assign t[31] = (x[4]);
  assign t[32] = (x[7]);
  assign t[33] = (x[7]);
  assign t[34] = (x[10]);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (t[20] & ~t[21]);
  assign t[17] = (t[22] & ~t[23]);
  assign t[18] = (t[24] & ~t[25]);
  assign t[19] = (t[26] & ~t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = t[35] ^ x[11];
  assign t[28] = (x[1]);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4]);
  assign t[31] = (x[4]);
  assign t[32] = (x[7]);
  assign t[33] = (x[7]);
  assign t[34] = (x[10]);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = (t[23] & ~t[24]);
  assign t[18] = (t[25] & ~t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[6];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[9];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[12];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = (x[1]);
  assign t[28] = (x[1]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7]);
  assign t[32] = (x[7]);
  assign t[33] = (x[10]);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = (t[23] & ~t[24]);
  assign t[18] = (t[25] & ~t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[6];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[9];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[12];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = (x[1]);
  assign t[28] = (x[1]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7]);
  assign t[32] = (x[7]);
  assign t[33] = (x[10]);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [10:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[4];
  assign t[12] = t[15] ^ x[7];
  assign t[13] = t[16] ^ x[10];
  assign t[14] = (t[17] & ~t[18]);
  assign t[15] = (t[19] & ~t[20]);
  assign t[16] = (t[21] & ~t[22]);
  assign t[17] = t[23] ^ x[4];
  assign t[18] = t[24] ^ x[3];
  assign t[19] = t[25] ^ x[7];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[10];
  assign t[22] = t[28] ^ x[9];
  assign t[23] = (x[2]);
  assign t[24] = (x[2]);
  assign t[25] = (x[5]);
  assign t[26] = (x[5]);
  assign t[27] = (x[8]);
  assign t[28] = (x[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[4];
  assign t[15] = t[19] ^ x[7];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[4];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[2]);
  assign t[32] = (x[5]);
  assign t[33] = (x[5]);
  assign t[34] = (x[8]);
  assign t[35] = (x[8]);
  assign t[36] = (x[11]);
  assign t[37] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [13:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[4];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[10];
  assign t[16] = t[20] ^ x[13];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[4];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[7];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[5]);
  assign t[32] = (x[5]);
  assign t[33] = (x[8]);
  assign t[34] = (x[8]);
  assign t[35] = (x[11]);
  assign t[36] = (x[11]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[142] | t[143]);
  assign t[105] = ~(t[144] | t[145]);
  assign t[106] = ~(t[226]);
  assign t[107] = ~(t[227]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[148] | t[149]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[228] | t[150]);
  assign t[111] = t[151] ? x[98] : x[97];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = ~(t[229]);
  assign t[114] = ~(t[230]);
  assign t[115] = ~(t[154] | t[155]);
  assign t[116] = t[204] ? x[106] : x[105];
  assign t[117] = t[156] | t[157];
  assign t[118] = ~(t[204]);
  assign t[119] = ~(t[158] & t[205]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[159] & t[160]);
  assign t[121] = ~(t[77] | t[161]);
  assign t[122] = ~(t[77] | t[162]);
  assign t[123] = t[205] & t[163];
  assign t[124] = t[159] | t[158];
  assign t[125] = ~(t[164] & t[160]);
  assign t[126] = ~(x[4] & t[165]);
  assign t[127] = ~(t[159] & t[205]);
  assign t[128] = ~(t[158] & t[160]);
  assign t[129] = ~(t[204]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[140]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[218] | t[219]);
  assign t[133] = ~(t[166] | t[144]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[232]);
  assign t[136] = ~(t[220] | t[221]);
  assign t[137] = ~(t[233]);
  assign t[138] = ~(t[234]);
  assign t[139] = ~(t[169] | t[170]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[171] | t[144]);
  assign t[141] = ~(t[172] | t[173]);
  assign t[142] = ~(t[235]);
  assign t[143] = ~(t[224] | t[225]);
  assign t[144] = ~(t[118] | t[174]);
  assign t[145] = t[175] | t[176];
  assign t[146] = ~(t[236]);
  assign t[147] = ~(t[226] | t[227]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[177] | t[178]);
  assign t[151] = ~(t[129]);
  assign t[152] = ~(t[156] | t[179]);
  assign t[153] = ~(t[47]);
  assign t[154] = ~(t[239]);
  assign t[155] = ~(t[229] | t[230]);
  assign t[156] = ~(t[180] & t[181]);
  assign t[157] = ~(t[182] & t[86]);
  assign t[158] = x[4] & t[203];
  assign t[159] = ~(x[4] | t[203]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[205]);
  assign t[161] = t[202] ? t[119] : t[120];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[118] | t[202]);
  assign t[164] = ~(x[4] | t[185]);
  assign t[165] = ~(t[203] | t[160]);
  assign t[166] = ~(t[118] | t[186]);
  assign t[167] = ~(t[31]);
  assign t[168] = ~(t[77] | t[187]);
  assign t[169] = ~(t[240]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[233] | t[234]);
  assign t[171] = ~(t[118] | t[188]);
  assign t[172] = ~(t[189] & t[190]);
  assign t[173] = ~(t[80] & t[191]);
  assign t[174] = t[202] ? t[125] : t[184];
  assign t[175] = ~(t[77] | t[192]);
  assign t[176] = ~(t[180]);
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[237] | t[238]);
  assign t[179] = ~(t[193] & t[191]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[163] & t[194]);
  assign t[181] = ~(t[165] & t[195]);
  assign t[182] = ~(t[47] | t[175]);
  assign t[183] = ~(t[205] & t[164]);
  assign t[184] = ~(x[4] & t[196]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[120] : t[128];
  assign t[187] = t[202] ? t[183] : t[184];
  assign t[188] = t[202] ? t[128] : t[120];
  assign t[189] = ~(t[166] | t[197]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[118] & t[198]);
  assign t[191] = t[118] | t[199];
  assign t[192] = t[202] ? t[127] : t[128];
  assign t[193] = ~(t[144]);
  assign t[194] = ~(t[183] & t[126]);
  assign t[195] = t[77] & t[202];
  assign t[196] = ~(t[203] | t[205]);
  assign t[197] = ~(t[77] | t[200]);
  assign t[198] = ~(t[184] & t[183]);
  assign t[199] = t[202] ? t[184] : t[125];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[125] : t[126];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[204] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[34]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[10];
  assign t[244] = t[285] ^ x[13];
  assign t[245] = t[286] ^ x[16];
  assign t[246] = t[287] ^ x[19];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[36];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = x[4] ? t[38] : t[37];
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[70];
  assign t[262] = t[303] ^ x[73];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[81];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[96];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = ~(t[41] ^ t[42]);
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = x[4] ? t[46] : t[45];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[47] | t[48]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[10];
  assign t[327] = t[409] ^ x[9];
  assign t[328] = t[410] ^ x[13];
  assign t[329] = t[411] ^ x[12];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[16];
  assign t[331] = t[413] ^ x[15];
  assign t[332] = t[414] ^ x[19];
  assign t[333] = t[415] ^ x[18];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[206] | t[53]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[36];
  assign t[343] = t[425] ^ x[35];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[54] ^ t[55]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[70];
  assign t[363] = t[445] ^ x[69];
  assign t[364] = t[446] ^ x[73];
  assign t[365] = t[447] ^ x[72];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[81];
  assign t[369] = t[451] ^ x[80];
  assign t[36] = ~(t[35] ^ t[58]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[96];
  assign t[379] = t[461] ^ x[95];
  assign t[37] = ~(t[59] | t[60]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[8]);
  assign t[409] = (x[8]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[11]);
  assign t[411] = (x[11]);
  assign t[412] = (x[14]);
  assign t[413] = (x[14]);
  assign t[414] = (x[17]);
  assign t[415] = (x[17]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[34]);
  assign t[425] = (x[34]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[68]);
  assign t[445] = (x[68]);
  assign t[446] = (x[71]);
  assign t[447] = (x[71]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[79]);
  assign t[451] = (x[79]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[94]);
  assign t[461] = (x[94]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[79] & t[80]);
  assign t[49] = ~(t[77] | t[81]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[77] | t[82]);
  assign t[51] = ~(t[208]);
  assign t[52] = ~(t[209]);
  assign t[53] = ~(t[83] | t[84]);
  assign t[54] = t[85] ? x[33] : x[32];
  assign t[55] = ~(t[86] & t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[210] | t[90]);
  assign t[58] = ~(t[91] ^ t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[211] | t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[212]);
  assign t[64] = ~(t[213]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[214] | t[104]);
  assign t[68] = t[204] ? x[50] : x[49];
  assign t[69] = ~(t[30] & t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[215] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[216] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118]);
  assign t[78] = t[202] ? t[120] : t[119];
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] & t[124]);
  assign t[81] = t[202] ? t[126] : t[125];
  assign t[82] = t[202] ? t[128] : t[127];
  assign t[83] = ~(t[217]);
  assign t[84] = ~(t[208] | t[209]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[122] | t[50]);
  assign t[87] = ~(t[123] | t[130]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = t[85] ? x[67] : x[66];
  assign t[92] = ~(t[133] & t[134]);
  assign t[93] = ~(t[220]);
  assign t[94] = ~(t[221]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = ~(t[137] | t[138]);
  assign t[97] = ~(t[222] | t[139]);
  assign t[98] = t[85] ? x[78] : x[77];
  assign t[99] = ~(t[140] & t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[142] | t[143]);
  assign t[105] = ~(t[144] | t[145]);
  assign t[106] = ~(t[226]);
  assign t[107] = ~(t[227]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[148] | t[149]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[228] | t[150]);
  assign t[111] = t[151] ? x[98] : x[97];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = ~(t[229]);
  assign t[114] = ~(t[230]);
  assign t[115] = ~(t[154] | t[155]);
  assign t[116] = t[204] ? x[106] : x[105];
  assign t[117] = t[156] | t[157];
  assign t[118] = ~(t[204]);
  assign t[119] = ~(t[158] & t[205]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[159] & t[160]);
  assign t[121] = ~(t[77] | t[161]);
  assign t[122] = ~(t[77] | t[162]);
  assign t[123] = t[205] & t[163];
  assign t[124] = t[159] | t[158];
  assign t[125] = ~(t[164] & t[160]);
  assign t[126] = ~(x[4] & t[165]);
  assign t[127] = ~(t[159] & t[205]);
  assign t[128] = ~(t[158] & t[160]);
  assign t[129] = ~(t[204]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[140]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[218] | t[219]);
  assign t[133] = ~(t[166] | t[144]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[232]);
  assign t[136] = ~(t[220] | t[221]);
  assign t[137] = ~(t[233]);
  assign t[138] = ~(t[234]);
  assign t[139] = ~(t[169] | t[170]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[171] | t[144]);
  assign t[141] = ~(t[172] | t[173]);
  assign t[142] = ~(t[235]);
  assign t[143] = ~(t[224] | t[225]);
  assign t[144] = ~(t[118] | t[174]);
  assign t[145] = t[175] | t[176];
  assign t[146] = ~(t[236]);
  assign t[147] = ~(t[226] | t[227]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[177] | t[178]);
  assign t[151] = ~(t[129]);
  assign t[152] = ~(t[156] | t[179]);
  assign t[153] = ~(t[47]);
  assign t[154] = ~(t[239]);
  assign t[155] = ~(t[229] | t[230]);
  assign t[156] = ~(t[180] & t[181]);
  assign t[157] = ~(t[182] & t[86]);
  assign t[158] = x[4] & t[203];
  assign t[159] = ~(x[4] | t[203]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[205]);
  assign t[161] = t[202] ? t[119] : t[120];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[118] | t[202]);
  assign t[164] = ~(x[4] | t[185]);
  assign t[165] = ~(t[203] | t[160]);
  assign t[166] = ~(t[118] | t[186]);
  assign t[167] = ~(t[31]);
  assign t[168] = ~(t[77] | t[187]);
  assign t[169] = ~(t[240]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[233] | t[234]);
  assign t[171] = ~(t[118] | t[188]);
  assign t[172] = ~(t[189] & t[190]);
  assign t[173] = ~(t[80] & t[191]);
  assign t[174] = t[202] ? t[125] : t[184];
  assign t[175] = ~(t[77] | t[192]);
  assign t[176] = ~(t[180]);
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[237] | t[238]);
  assign t[179] = ~(t[193] & t[191]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[163] & t[194]);
  assign t[181] = ~(t[165] & t[195]);
  assign t[182] = ~(t[47] | t[175]);
  assign t[183] = ~(t[205] & t[164]);
  assign t[184] = ~(x[4] & t[196]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[120] : t[128];
  assign t[187] = t[202] ? t[183] : t[184];
  assign t[188] = t[202] ? t[128] : t[120];
  assign t[189] = ~(t[166] | t[197]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[118] & t[198]);
  assign t[191] = t[118] | t[199];
  assign t[192] = t[202] ? t[127] : t[128];
  assign t[193] = ~(t[144]);
  assign t[194] = ~(t[183] & t[126]);
  assign t[195] = t[77] & t[202];
  assign t[196] = ~(t[203] | t[205]);
  assign t[197] = ~(t[77] | t[200]);
  assign t[198] = ~(t[184] & t[183]);
  assign t[199] = t[202] ? t[184] : t[125];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[125] : t[126];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[204] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[34]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[10];
  assign t[244] = t[285] ^ x[13];
  assign t[245] = t[286] ^ x[16];
  assign t[246] = t[287] ^ x[19];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[36];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = x[4] ? t[38] : t[37];
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[70];
  assign t[262] = t[303] ^ x[73];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[81];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[96];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = ~(t[41] ^ t[42]);
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = x[4] ? t[46] : t[45];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[47] | t[48]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[10];
  assign t[327] = t[409] ^ x[9];
  assign t[328] = t[410] ^ x[13];
  assign t[329] = t[411] ^ x[12];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[16];
  assign t[331] = t[413] ^ x[15];
  assign t[332] = t[414] ^ x[19];
  assign t[333] = t[415] ^ x[18];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[206] | t[53]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[36];
  assign t[343] = t[425] ^ x[35];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[54] ^ t[55]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[70];
  assign t[363] = t[445] ^ x[69];
  assign t[364] = t[446] ^ x[73];
  assign t[365] = t[447] ^ x[72];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[81];
  assign t[369] = t[451] ^ x[80];
  assign t[36] = ~(t[35] ^ t[58]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[96];
  assign t[379] = t[461] ^ x[95];
  assign t[37] = ~(t[59] | t[60]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[8]);
  assign t[409] = (x[8]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[11]);
  assign t[411] = (x[11]);
  assign t[412] = (x[14]);
  assign t[413] = (x[14]);
  assign t[414] = (x[17]);
  assign t[415] = (x[17]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[34]);
  assign t[425] = (x[34]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[68]);
  assign t[445] = (x[68]);
  assign t[446] = (x[71]);
  assign t[447] = (x[71]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[79]);
  assign t[451] = (x[79]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[94]);
  assign t[461] = (x[94]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[79] & t[80]);
  assign t[49] = ~(t[77] | t[81]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[77] | t[82]);
  assign t[51] = ~(t[208]);
  assign t[52] = ~(t[209]);
  assign t[53] = ~(t[83] | t[84]);
  assign t[54] = t[85] ? x[33] : x[32];
  assign t[55] = ~(t[86] & t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[210] | t[90]);
  assign t[58] = ~(t[91] ^ t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[211] | t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[212]);
  assign t[64] = ~(t[213]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[214] | t[104]);
  assign t[68] = t[204] ? x[50] : x[49];
  assign t[69] = ~(t[30] & t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[215] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[216] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118]);
  assign t[78] = t[202] ? t[120] : t[119];
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] & t[124]);
  assign t[81] = t[202] ? t[126] : t[125];
  assign t[82] = t[202] ? t[128] : t[127];
  assign t[83] = ~(t[217]);
  assign t[84] = ~(t[208] | t[209]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[122] | t[50]);
  assign t[87] = ~(t[123] | t[130]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = t[85] ? x[67] : x[66];
  assign t[92] = ~(t[133] & t[134]);
  assign t[93] = ~(t[220]);
  assign t[94] = ~(t[221]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = ~(t[137] | t[138]);
  assign t[97] = ~(t[222] | t[139]);
  assign t[98] = t[85] ? x[78] : x[77];
  assign t[99] = ~(t[140] & t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [112:0] x;
 output y;

 wire [313:0] t;
  assign t[0] = t[1] ? t[2] : t[90];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = t[154] ^ x[2];
  assign t[123] = t[155] ^ x[8];
  assign t[124] = t[156] ^ x[11];
  assign t[125] = t[157] ^ x[14];
  assign t[126] = t[158] ^ x[17];
  assign t[127] = t[159] ^ x[22];
  assign t[128] = t[160] ^ x[25];
  assign t[129] = t[161] ^ x[30];
  assign t[12] = t[93] ? x[18] : x[19];
  assign t[130] = t[162] ^ x[33];
  assign t[131] = t[163] ^ x[38];
  assign t[132] = t[164] ^ x[41];
  assign t[133] = t[165] ^ x[44];
  assign t[134] = t[166] ^ x[49];
  assign t[135] = t[167] ^ x[52];
  assign t[136] = t[168] ^ x[57];
  assign t[137] = t[169] ^ x[60];
  assign t[138] = t[170] ^ x[63];
  assign t[139] = t[171] ^ x[66];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[69];
  assign t[141] = t[173] ^ x[74];
  assign t[142] = t[174] ^ x[77];
  assign t[143] = t[175] ^ x[82];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[88];
  assign t[146] = t[178] ^ x[91];
  assign t[147] = t[179] ^ x[94];
  assign t[148] = t[180] ^ x[97];
  assign t[149] = t[181] ^ x[100];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[103];
  assign t[151] = t[183] ^ x[106];
  assign t[152] = t[184] ^ x[109];
  assign t[153] = t[185] ^ x[112];
  assign t[154] = (t[186] & ~t[187]);
  assign t[155] = (t[188] & ~t[189]);
  assign t[156] = (t[190] & ~t[191]);
  assign t[157] = (t[192] & ~t[193]);
  assign t[158] = (t[194] & ~t[195]);
  assign t[159] = (t[196] & ~t[197]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (t[198] & ~t[199]);
  assign t[161] = (t[200] & ~t[201]);
  assign t[162] = (t[202] & ~t[203]);
  assign t[163] = (t[204] & ~t[205]);
  assign t[164] = (t[206] & ~t[207]);
  assign t[165] = (t[208] & ~t[209]);
  assign t[166] = (t[210] & ~t[211]);
  assign t[167] = (t[212] & ~t[213]);
  assign t[168] = (t[214] & ~t[215]);
  assign t[169] = (t[216] & ~t[217]);
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = (t[218] & ~t[219]);
  assign t[171] = (t[220] & ~t[221]);
  assign t[172] = (t[222] & ~t[223]);
  assign t[173] = (t[224] & ~t[225]);
  assign t[174] = (t[226] & ~t[227]);
  assign t[175] = (t[228] & ~t[229]);
  assign t[176] = (t[230] & ~t[231]);
  assign t[177] = (t[232] & ~t[233]);
  assign t[178] = (t[234] & ~t[235]);
  assign t[179] = (t[236] & ~t[237]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (t[238] & ~t[239]);
  assign t[181] = (t[240] & ~t[241]);
  assign t[182] = (t[242] & ~t[243]);
  assign t[183] = (t[244] & ~t[245]);
  assign t[184] = (t[246] & ~t[247]);
  assign t[185] = (t[248] & ~t[249]);
  assign t[186] = t[250] ^ x[2];
  assign t[187] = t[251] ^ x[1];
  assign t[188] = t[252] ^ x[8];
  assign t[189] = t[253] ^ x[7];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[254] ^ x[11];
  assign t[191] = t[255] ^ x[10];
  assign t[192] = t[256] ^ x[14];
  assign t[193] = t[257] ^ x[13];
  assign t[194] = t[258] ^ x[17];
  assign t[195] = t[259] ^ x[16];
  assign t[196] = t[260] ^ x[22];
  assign t[197] = t[261] ^ x[21];
  assign t[198] = t[262] ^ x[25];
  assign t[199] = t[263] ^ x[24];
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[264] ^ x[30];
  assign t[201] = t[265] ^ x[29];
  assign t[202] = t[266] ^ x[33];
  assign t[203] = t[267] ^ x[32];
  assign t[204] = t[268] ^ x[38];
  assign t[205] = t[269] ^ x[37];
  assign t[206] = t[270] ^ x[41];
  assign t[207] = t[271] ^ x[40];
  assign t[208] = t[272] ^ x[44];
  assign t[209] = t[273] ^ x[43];
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = t[274] ^ x[49];
  assign t[211] = t[275] ^ x[48];
  assign t[212] = t[276] ^ x[52];
  assign t[213] = t[277] ^ x[51];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[56];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[59];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[62];
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[65];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[68];
  assign t[224] = t[288] ^ x[74];
  assign t[225] = t[289] ^ x[73];
  assign t[226] = t[290] ^ x[77];
  assign t[227] = t[291] ^ x[76];
  assign t[228] = t[292] ^ x[82];
  assign t[229] = t[293] ^ x[81];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[294] ^ x[85];
  assign t[231] = t[295] ^ x[84];
  assign t[232] = t[296] ^ x[88];
  assign t[233] = t[297] ^ x[87];
  assign t[234] = t[298] ^ x[91];
  assign t[235] = t[299] ^ x[90];
  assign t[236] = t[300] ^ x[94];
  assign t[237] = t[301] ^ x[93];
  assign t[238] = t[302] ^ x[97];
  assign t[239] = t[303] ^ x[96];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[304] ^ x[100];
  assign t[241] = t[305] ^ x[99];
  assign t[242] = t[306] ^ x[103];
  assign t[243] = t[307] ^ x[102];
  assign t[244] = t[308] ^ x[106];
  assign t[245] = t[309] ^ x[105];
  assign t[246] = t[310] ^ x[109];
  assign t[247] = t[311] ^ x[108];
  assign t[248] = t[312] ^ x[112];
  assign t[249] = t[313] ^ x[111];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[0]);
  assign t[251] = (x[0]);
  assign t[252] = (x[6]);
  assign t[253] = (x[6]);
  assign t[254] = (x[9]);
  assign t[255] = (x[9]);
  assign t[256] = (x[12]);
  assign t[257] = (x[12]);
  assign t[258] = (x[15]);
  assign t[259] = (x[15]);
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = (x[20]);
  assign t[261] = (x[20]);
  assign t[262] = (x[23]);
  assign t[263] = (x[23]);
  assign t[264] = (x[28]);
  assign t[265] = (x[28]);
  assign t[266] = (x[31]);
  assign t[267] = (x[31]);
  assign t[268] = (x[36]);
  assign t[269] = (x[36]);
  assign t[26] = ~(t[95] & t[41]);
  assign t[270] = (x[39]);
  assign t[271] = (x[39]);
  assign t[272] = (x[42]);
  assign t[273] = (x[42]);
  assign t[274] = (x[47]);
  assign t[275] = (x[47]);
  assign t[276] = (x[50]);
  assign t[277] = (x[50]);
  assign t[278] = (x[55]);
  assign t[279] = (x[55]);
  assign t[27] = ~(t[96] & t[42]);
  assign t[280] = (x[58]);
  assign t[281] = (x[58]);
  assign t[282] = (x[61]);
  assign t[283] = (x[61]);
  assign t[284] = (x[64]);
  assign t[285] = (x[64]);
  assign t[286] = (x[67]);
  assign t[287] = (x[67]);
  assign t[288] = (x[72]);
  assign t[289] = (x[72]);
  assign t[28] = t[43] ? x[27] : x[26];
  assign t[290] = (x[75]);
  assign t[291] = (x[75]);
  assign t[292] = (x[80]);
  assign t[293] = (x[80]);
  assign t[294] = (x[83]);
  assign t[295] = (x[83]);
  assign t[296] = (x[86]);
  assign t[297] = (x[86]);
  assign t[298] = (x[89]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[92]);
  assign t[301] = (x[92]);
  assign t[302] = (x[95]);
  assign t[303] = (x[95]);
  assign t[304] = (x[98]);
  assign t[305] = (x[98]);
  assign t[306] = (x[101]);
  assign t[307] = (x[101]);
  assign t[308] = (x[104]);
  assign t[309] = (x[104]);
  assign t[30] = t[46] ^ t[47];
  assign t[310] = (x[107]);
  assign t[311] = (x[107]);
  assign t[312] = (x[110]);
  assign t[313] = (x[110]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[31];
  assign t[33] = ~(t[97] & t[51]);
  assign t[34] = ~(t[98] & t[52]);
  assign t[35] = t[43] ? x[35] : x[34];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] ^ t[37];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[99]);
  assign t[42] = ~(t[99] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[100] & t[64]);
  assign t[45] = ~(t[101] & t[65]);
  assign t[46] = t[43] ? x[46] : x[45];
  assign t[47] = ~(t[66] & t[67]);
  assign t[48] = ~(t[102] & t[68]);
  assign t[49] = ~(t[103] & t[69]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[43] ? x[54] : x[53];
  assign t[51] = ~(t[104]);
  assign t[52] = ~(t[104] & t[70]);
  assign t[53] = ~(t[105] & t[71]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = t[93] ? x[71] : x[70];
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[93] ? x[79] : x[78];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[95]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[111]);
  assign t[65] = ~(t[111] & t[79]);
  assign t[66] = ~(t[112] & t[80]);
  assign t[67] = ~(t[113] & t[81]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[97]);
  assign t[71] = ~(t[115]);
  assign t[72] = ~(t[115] & t[83]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117]);
  assign t[76] = ~(t[117] & t[85]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[100]);
  assign t[7] = ~(t[91] & t[92]);
  assign t[80] = ~(t[120]);
  assign t[81] = ~(t[120] & t[88]);
  assign t[82] = ~(t[102]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[107]);
  assign t[85] = ~(t[109]);
  assign t[86] = ~(t[121]);
  assign t[87] = ~(t[121] & t[89]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[118]);
  assign t[8] = ~(t[93] & t[94]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [112:0] x;
 output y;

 wire [313:0] t;
  assign t[0] = t[1] ? t[2] : t[90];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = t[154] ^ x[2];
  assign t[123] = t[155] ^ x[8];
  assign t[124] = t[156] ^ x[11];
  assign t[125] = t[157] ^ x[14];
  assign t[126] = t[158] ^ x[17];
  assign t[127] = t[159] ^ x[22];
  assign t[128] = t[160] ^ x[25];
  assign t[129] = t[161] ^ x[30];
  assign t[12] = t[93] ? x[18] : x[19];
  assign t[130] = t[162] ^ x[33];
  assign t[131] = t[163] ^ x[38];
  assign t[132] = t[164] ^ x[41];
  assign t[133] = t[165] ^ x[44];
  assign t[134] = t[166] ^ x[49];
  assign t[135] = t[167] ^ x[52];
  assign t[136] = t[168] ^ x[57];
  assign t[137] = t[169] ^ x[60];
  assign t[138] = t[170] ^ x[63];
  assign t[139] = t[171] ^ x[66];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[69];
  assign t[141] = t[173] ^ x[74];
  assign t[142] = t[174] ^ x[77];
  assign t[143] = t[175] ^ x[82];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[88];
  assign t[146] = t[178] ^ x[91];
  assign t[147] = t[179] ^ x[94];
  assign t[148] = t[180] ^ x[97];
  assign t[149] = t[181] ^ x[100];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[103];
  assign t[151] = t[183] ^ x[106];
  assign t[152] = t[184] ^ x[109];
  assign t[153] = t[185] ^ x[112];
  assign t[154] = (t[186] & ~t[187]);
  assign t[155] = (t[188] & ~t[189]);
  assign t[156] = (t[190] & ~t[191]);
  assign t[157] = (t[192] & ~t[193]);
  assign t[158] = (t[194] & ~t[195]);
  assign t[159] = (t[196] & ~t[197]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (t[198] & ~t[199]);
  assign t[161] = (t[200] & ~t[201]);
  assign t[162] = (t[202] & ~t[203]);
  assign t[163] = (t[204] & ~t[205]);
  assign t[164] = (t[206] & ~t[207]);
  assign t[165] = (t[208] & ~t[209]);
  assign t[166] = (t[210] & ~t[211]);
  assign t[167] = (t[212] & ~t[213]);
  assign t[168] = (t[214] & ~t[215]);
  assign t[169] = (t[216] & ~t[217]);
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = (t[218] & ~t[219]);
  assign t[171] = (t[220] & ~t[221]);
  assign t[172] = (t[222] & ~t[223]);
  assign t[173] = (t[224] & ~t[225]);
  assign t[174] = (t[226] & ~t[227]);
  assign t[175] = (t[228] & ~t[229]);
  assign t[176] = (t[230] & ~t[231]);
  assign t[177] = (t[232] & ~t[233]);
  assign t[178] = (t[234] & ~t[235]);
  assign t[179] = (t[236] & ~t[237]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (t[238] & ~t[239]);
  assign t[181] = (t[240] & ~t[241]);
  assign t[182] = (t[242] & ~t[243]);
  assign t[183] = (t[244] & ~t[245]);
  assign t[184] = (t[246] & ~t[247]);
  assign t[185] = (t[248] & ~t[249]);
  assign t[186] = t[250] ^ x[2];
  assign t[187] = t[251] ^ x[1];
  assign t[188] = t[252] ^ x[8];
  assign t[189] = t[253] ^ x[7];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[254] ^ x[11];
  assign t[191] = t[255] ^ x[10];
  assign t[192] = t[256] ^ x[14];
  assign t[193] = t[257] ^ x[13];
  assign t[194] = t[258] ^ x[17];
  assign t[195] = t[259] ^ x[16];
  assign t[196] = t[260] ^ x[22];
  assign t[197] = t[261] ^ x[21];
  assign t[198] = t[262] ^ x[25];
  assign t[199] = t[263] ^ x[24];
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[264] ^ x[30];
  assign t[201] = t[265] ^ x[29];
  assign t[202] = t[266] ^ x[33];
  assign t[203] = t[267] ^ x[32];
  assign t[204] = t[268] ^ x[38];
  assign t[205] = t[269] ^ x[37];
  assign t[206] = t[270] ^ x[41];
  assign t[207] = t[271] ^ x[40];
  assign t[208] = t[272] ^ x[44];
  assign t[209] = t[273] ^ x[43];
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = t[274] ^ x[49];
  assign t[211] = t[275] ^ x[48];
  assign t[212] = t[276] ^ x[52];
  assign t[213] = t[277] ^ x[51];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[56];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[59];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[62];
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[65];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[68];
  assign t[224] = t[288] ^ x[74];
  assign t[225] = t[289] ^ x[73];
  assign t[226] = t[290] ^ x[77];
  assign t[227] = t[291] ^ x[76];
  assign t[228] = t[292] ^ x[82];
  assign t[229] = t[293] ^ x[81];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[294] ^ x[85];
  assign t[231] = t[295] ^ x[84];
  assign t[232] = t[296] ^ x[88];
  assign t[233] = t[297] ^ x[87];
  assign t[234] = t[298] ^ x[91];
  assign t[235] = t[299] ^ x[90];
  assign t[236] = t[300] ^ x[94];
  assign t[237] = t[301] ^ x[93];
  assign t[238] = t[302] ^ x[97];
  assign t[239] = t[303] ^ x[96];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[304] ^ x[100];
  assign t[241] = t[305] ^ x[99];
  assign t[242] = t[306] ^ x[103];
  assign t[243] = t[307] ^ x[102];
  assign t[244] = t[308] ^ x[106];
  assign t[245] = t[309] ^ x[105];
  assign t[246] = t[310] ^ x[109];
  assign t[247] = t[311] ^ x[108];
  assign t[248] = t[312] ^ x[112];
  assign t[249] = t[313] ^ x[111];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[0]);
  assign t[251] = (x[0]);
  assign t[252] = (x[6]);
  assign t[253] = (x[6]);
  assign t[254] = (x[9]);
  assign t[255] = (x[9]);
  assign t[256] = (x[12]);
  assign t[257] = (x[12]);
  assign t[258] = (x[15]);
  assign t[259] = (x[15]);
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = (x[20]);
  assign t[261] = (x[20]);
  assign t[262] = (x[23]);
  assign t[263] = (x[23]);
  assign t[264] = (x[28]);
  assign t[265] = (x[28]);
  assign t[266] = (x[31]);
  assign t[267] = (x[31]);
  assign t[268] = (x[36]);
  assign t[269] = (x[36]);
  assign t[26] = ~(t[95] & t[41]);
  assign t[270] = (x[39]);
  assign t[271] = (x[39]);
  assign t[272] = (x[42]);
  assign t[273] = (x[42]);
  assign t[274] = (x[47]);
  assign t[275] = (x[47]);
  assign t[276] = (x[50]);
  assign t[277] = (x[50]);
  assign t[278] = (x[55]);
  assign t[279] = (x[55]);
  assign t[27] = ~(t[96] & t[42]);
  assign t[280] = (x[58]);
  assign t[281] = (x[58]);
  assign t[282] = (x[61]);
  assign t[283] = (x[61]);
  assign t[284] = (x[64]);
  assign t[285] = (x[64]);
  assign t[286] = (x[67]);
  assign t[287] = (x[67]);
  assign t[288] = (x[72]);
  assign t[289] = (x[72]);
  assign t[28] = t[43] ? x[27] : x[26];
  assign t[290] = (x[75]);
  assign t[291] = (x[75]);
  assign t[292] = (x[80]);
  assign t[293] = (x[80]);
  assign t[294] = (x[83]);
  assign t[295] = (x[83]);
  assign t[296] = (x[86]);
  assign t[297] = (x[86]);
  assign t[298] = (x[89]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[92]);
  assign t[301] = (x[92]);
  assign t[302] = (x[95]);
  assign t[303] = (x[95]);
  assign t[304] = (x[98]);
  assign t[305] = (x[98]);
  assign t[306] = (x[101]);
  assign t[307] = (x[101]);
  assign t[308] = (x[104]);
  assign t[309] = (x[104]);
  assign t[30] = t[46] ^ t[47];
  assign t[310] = (x[107]);
  assign t[311] = (x[107]);
  assign t[312] = (x[110]);
  assign t[313] = (x[110]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[31];
  assign t[33] = ~(t[97] & t[51]);
  assign t[34] = ~(t[98] & t[52]);
  assign t[35] = t[43] ? x[35] : x[34];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] ^ t[37];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[99]);
  assign t[42] = ~(t[99] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[100] & t[64]);
  assign t[45] = ~(t[101] & t[65]);
  assign t[46] = t[43] ? x[46] : x[45];
  assign t[47] = ~(t[66] & t[67]);
  assign t[48] = ~(t[102] & t[68]);
  assign t[49] = ~(t[103] & t[69]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[43] ? x[54] : x[53];
  assign t[51] = ~(t[104]);
  assign t[52] = ~(t[104] & t[70]);
  assign t[53] = ~(t[105] & t[71]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = t[93] ? x[71] : x[70];
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[93] ? x[79] : x[78];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[95]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[111]);
  assign t[65] = ~(t[111] & t[79]);
  assign t[66] = ~(t[112] & t[80]);
  assign t[67] = ~(t[113] & t[81]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[97]);
  assign t[71] = ~(t[115]);
  assign t[72] = ~(t[115] & t[83]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117]);
  assign t[76] = ~(t[117] & t[85]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[100]);
  assign t[7] = ~(t[91] & t[92]);
  assign t[80] = ~(t[120]);
  assign t[81] = ~(t[120] & t[88]);
  assign t[82] = ~(t[102]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[107]);
  assign t[85] = ~(t[109]);
  assign t[86] = ~(t[121]);
  assign t[87] = ~(t[121] & t[89]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[118]);
  assign t[8] = ~(t[93] & t[94]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[109] & t[110]);
  assign t[105] = ~(t[140] & t[139]);
  assign t[106] = ~(t[149]);
  assign t[107] = ~(t[144] & t[143]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[148] & t[147]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[112] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[112] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = t[30] ^ t[24];
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = ~(t[35] & t[36]);
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = t[37] ^ t[38];
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = x[4] ? t[40] : t[39];
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = ~(t[43] & t[44]);
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = ~(t[45] & t[116]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = t[46] ? x[24] : x[23];
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[49] ^ t[31];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[52] ^ t[53];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[54] & t[55]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[56] & t[117]);
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = t[57] ? x[29] : x[28];
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[118]);
  assign t[44] = ~(t[119]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[120]);
  assign t[49] = t[46] ? x[40] : x[39];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[121]);
  assign t[52] = t[46] ? x[45] : x[44];
  assign t[53] = ~(t[76] & t[77]);
  assign t[54] = ~(t[122]);
  assign t[55] = ~(t[123]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[69]);
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[124]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[125]);
  assign t[62] = t[112] ? x[59] : x[58];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[126]);
  assign t[66] = t[112] ? x[64] : x[63];
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[112]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[93] & t[94]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[97] & t[132]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[103]);
  assign t[87] = ~(t[104] & t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[107] & t[108]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[109] & t[110]);
  assign t[105] = ~(t[140] & t[139]);
  assign t[106] = ~(t[149]);
  assign t[107] = ~(t[144] & t[143]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[148] & t[147]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[112] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[112] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = t[30] ^ t[24];
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = ~(t[35] & t[36]);
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = t[37] ^ t[38];
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = x[4] ? t[40] : t[39];
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = ~(t[43] & t[44]);
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = ~(t[45] & t[116]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = t[46] ? x[24] : x[23];
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[49] ^ t[31];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[52] ^ t[53];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[54] & t[55]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[56] & t[117]);
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = t[57] ? x[29] : x[28];
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[118]);
  assign t[44] = ~(t[119]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[120]);
  assign t[49] = t[46] ? x[40] : x[39];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[121]);
  assign t[52] = t[46] ? x[45] : x[44];
  assign t[53] = ~(t[76] & t[77]);
  assign t[54] = ~(t[122]);
  assign t[55] = ~(t[123]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[69]);
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[124]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[125]);
  assign t[62] = t[112] ? x[59] : x[58];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[126]);
  assign t[66] = t[112] ? x[64] : x[63];
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[112]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[93] & t[94]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[97] & t[132]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[103]);
  assign t[87] = ~(t[104] & t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[107] & t[108]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [139:0] x;
 output y;

 wire [386:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[2];
  assign t[142] = t[183] ^ x[8];
  assign t[143] = t[184] ^ x[11];
  assign t[144] = t[185] ^ x[14];
  assign t[145] = t[186] ^ x[17];
  assign t[146] = t[187] ^ x[22];
  assign t[147] = t[188] ^ x[27];
  assign t[148] = t[189] ^ x[32];
  assign t[149] = t[190] ^ x[35];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[38];
  assign t[151] = t[192] ^ x[43];
  assign t[152] = t[193] ^ x[48];
  assign t[153] = t[194] ^ x[51];
  assign t[154] = t[195] ^ x[54];
  assign t[155] = t[196] ^ x[57];
  assign t[156] = t[197] ^ x[62];
  assign t[157] = t[198] ^ x[67];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[73];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[76];
  assign t[161] = t[202] ^ x[79];
  assign t[162] = t[203] ^ x[82];
  assign t[163] = t[204] ^ x[85];
  assign t[164] = t[205] ^ x[88];
  assign t[165] = t[206] ^ x[91];
  assign t[166] = t[207] ^ x[94];
  assign t[167] = t[208] ^ x[97];
  assign t[168] = t[209] ^ x[100];
  assign t[169] = t[210] ^ x[103];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[106];
  assign t[171] = t[212] ^ x[109];
  assign t[172] = t[213] ^ x[112];
  assign t[173] = t[214] ^ x[115];
  assign t[174] = t[215] ^ x[118];
  assign t[175] = t[216] ^ x[121];
  assign t[176] = t[217] ^ x[124];
  assign t[177] = t[218] ^ x[127];
  assign t[178] = t[219] ^ x[130];
  assign t[179] = t[220] ^ x[133];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[136];
  assign t[181] = t[222] ^ x[139];
  assign t[182] = (t[223] & ~t[224]);
  assign t[183] = (t[225] & ~t[226]);
  assign t[184] = (t[227] & ~t[228]);
  assign t[185] = (t[229] & ~t[230]);
  assign t[186] = (t[231] & ~t[232]);
  assign t[187] = (t[233] & ~t[234]);
  assign t[188] = (t[235] & ~t[236]);
  assign t[189] = (t[237] & ~t[238]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[239] & ~t[240]);
  assign t[191] = (t[241] & ~t[242]);
  assign t[192] = (t[243] & ~t[244]);
  assign t[193] = (t[245] & ~t[246]);
  assign t[194] = (t[247] & ~t[248]);
  assign t[195] = (t[249] & ~t[250]);
  assign t[196] = (t[251] & ~t[252]);
  assign t[197] = (t[253] & ~t[254]);
  assign t[198] = (t[255] & ~t[256]);
  assign t[199] = (t[257] & ~t[258]);
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[259] & ~t[260]);
  assign t[201] = (t[261] & ~t[262]);
  assign t[202] = (t[263] & ~t[264]);
  assign t[203] = (t[265] & ~t[266]);
  assign t[204] = (t[267] & ~t[268]);
  assign t[205] = (t[269] & ~t[270]);
  assign t[206] = (t[271] & ~t[272]);
  assign t[207] = (t[273] & ~t[274]);
  assign t[208] = (t[275] & ~t[276]);
  assign t[209] = (t[277] & ~t[278]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = (t[279] & ~t[280]);
  assign t[211] = (t[281] & ~t[282]);
  assign t[212] = (t[283] & ~t[284]);
  assign t[213] = (t[285] & ~t[286]);
  assign t[214] = (t[287] & ~t[288]);
  assign t[215] = (t[289] & ~t[290]);
  assign t[216] = (t[291] & ~t[292]);
  assign t[217] = (t[293] & ~t[294]);
  assign t[218] = (t[295] & ~t[296]);
  assign t[219] = (t[297] & ~t[298]);
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[220] = (t[299] & ~t[300]);
  assign t[221] = (t[301] & ~t[302]);
  assign t[222] = (t[303] & ~t[304]);
  assign t[223] = t[305] ^ x[2];
  assign t[224] = t[306] ^ x[1];
  assign t[225] = t[307] ^ x[8];
  assign t[226] = t[308] ^ x[7];
  assign t[227] = t[309] ^ x[11];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[14];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[17];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[22];
  assign t[234] = t[316] ^ x[21];
  assign t[235] = t[317] ^ x[27];
  assign t[236] = t[318] ^ x[26];
  assign t[237] = t[319] ^ x[32];
  assign t[238] = t[320] ^ x[31];
  assign t[239] = t[321] ^ x[35];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[322] ^ x[34];
  assign t[241] = t[323] ^ x[38];
  assign t[242] = t[324] ^ x[37];
  assign t[243] = t[325] ^ x[43];
  assign t[244] = t[326] ^ x[42];
  assign t[245] = t[327] ^ x[48];
  assign t[246] = t[328] ^ x[47];
  assign t[247] = t[329] ^ x[51];
  assign t[248] = t[330] ^ x[50];
  assign t[249] = t[331] ^ x[54];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[53];
  assign t[251] = t[333] ^ x[57];
  assign t[252] = t[334] ^ x[56];
  assign t[253] = t[335] ^ x[62];
  assign t[254] = t[336] ^ x[61];
  assign t[255] = t[337] ^ x[67];
  assign t[256] = t[338] ^ x[66];
  assign t[257] = t[339] ^ x[70];
  assign t[258] = t[340] ^ x[69];
  assign t[259] = t[341] ^ x[73];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[72];
  assign t[261] = t[343] ^ x[76];
  assign t[262] = t[344] ^ x[75];
  assign t[263] = t[345] ^ x[79];
  assign t[264] = t[346] ^ x[78];
  assign t[265] = t[347] ^ x[82];
  assign t[266] = t[348] ^ x[81];
  assign t[267] = t[349] ^ x[85];
  assign t[268] = t[350] ^ x[84];
  assign t[269] = t[351] ^ x[88];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[87];
  assign t[271] = t[353] ^ x[91];
  assign t[272] = t[354] ^ x[90];
  assign t[273] = t[355] ^ x[94];
  assign t[274] = t[356] ^ x[93];
  assign t[275] = t[357] ^ x[97];
  assign t[276] = t[358] ^ x[96];
  assign t[277] = t[359] ^ x[100];
  assign t[278] = t[360] ^ x[99];
  assign t[279] = t[361] ^ x[103];
  assign t[27] = t[43] | t[105];
  assign t[280] = t[362] ^ x[102];
  assign t[281] = t[363] ^ x[106];
  assign t[282] = t[364] ^ x[105];
  assign t[283] = t[365] ^ x[109];
  assign t[284] = t[366] ^ x[108];
  assign t[285] = t[367] ^ x[112];
  assign t[286] = t[368] ^ x[111];
  assign t[287] = t[369] ^ x[115];
  assign t[288] = t[370] ^ x[114];
  assign t[289] = t[371] ^ x[118];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[117];
  assign t[291] = t[373] ^ x[121];
  assign t[292] = t[374] ^ x[120];
  assign t[293] = t[375] ^ x[124];
  assign t[294] = t[376] ^ x[123];
  assign t[295] = t[377] ^ x[127];
  assign t[296] = t[378] ^ x[126];
  assign t[297] = t[379] ^ x[130];
  assign t[298] = t[380] ^ x[129];
  assign t[299] = t[381] ^ x[133];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[132];
  assign t[301] = t[383] ^ x[136];
  assign t[302] = t[384] ^ x[135];
  assign t[303] = t[385] ^ x[139];
  assign t[304] = t[386] ^ x[138];
  assign t[305] = (x[0]);
  assign t[306] = (x[0]);
  assign t[307] = (x[6]);
  assign t[308] = (x[6]);
  assign t[309] = (x[9]);
  assign t[30] = t[47] ^ t[29];
  assign t[310] = (x[9]);
  assign t[311] = (x[12]);
  assign t[312] = (x[12]);
  assign t[313] = (x[15]);
  assign t[314] = (x[15]);
  assign t[315] = (x[20]);
  assign t[316] = (x[20]);
  assign t[317] = (x[25]);
  assign t[318] = (x[25]);
  assign t[319] = (x[30]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = (x[30]);
  assign t[321] = (x[33]);
  assign t[322] = (x[33]);
  assign t[323] = (x[36]);
  assign t[324] = (x[36]);
  assign t[325] = (x[41]);
  assign t[326] = (x[41]);
  assign t[327] = (x[46]);
  assign t[328] = (x[46]);
  assign t[329] = (x[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[330] = (x[49]);
  assign t[331] = (x[52]);
  assign t[332] = (x[52]);
  assign t[333] = (x[55]);
  assign t[334] = (x[55]);
  assign t[335] = (x[60]);
  assign t[336] = (x[60]);
  assign t[337] = (x[65]);
  assign t[338] = (x[65]);
  assign t[339] = (x[68]);
  assign t[33] = ~(t[52] & t[53]);
  assign t[340] = (x[68]);
  assign t[341] = (x[71]);
  assign t[342] = (x[71]);
  assign t[343] = (x[74]);
  assign t[344] = (x[74]);
  assign t[345] = (x[77]);
  assign t[346] = (x[77]);
  assign t[347] = (x[80]);
  assign t[348] = (x[80]);
  assign t[349] = (x[83]);
  assign t[34] = t[54] | t[106];
  assign t[350] = (x[83]);
  assign t[351] = (x[86]);
  assign t[352] = (x[86]);
  assign t[353] = (x[89]);
  assign t[354] = (x[89]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[98]);
  assign t[35] = t[55] ? x[29] : x[28];
  assign t[360] = (x[98]);
  assign t[361] = (x[101]);
  assign t[362] = (x[101]);
  assign t[363] = (x[104]);
  assign t[364] = (x[104]);
  assign t[365] = (x[107]);
  assign t[366] = (x[107]);
  assign t[367] = (x[110]);
  assign t[368] = (x[110]);
  assign t[369] = (x[113]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[113]);
  assign t[371] = (x[116]);
  assign t[372] = (x[116]);
  assign t[373] = (x[119]);
  assign t[374] = (x[119]);
  assign t[375] = (x[122]);
  assign t[376] = (x[122]);
  assign t[377] = (x[125]);
  assign t[378] = (x[125]);
  assign t[379] = (x[128]);
  assign t[37] = ~(t[58] & t[59]);
  assign t[380] = (x[128]);
  assign t[381] = (x[131]);
  assign t[382] = (x[131]);
  assign t[383] = (x[134]);
  assign t[384] = (x[134]);
  assign t[385] = (x[137]);
  assign t[386] = (x[137]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[62] & t[63]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[64] ^ t[39];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[65] | t[41]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = t[69] | t[109];
  assign t[47] = t[44] ? x[40] : x[39];
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = t[72] | t[110];
  assign t[4] = ~(x[3]);
  assign t[50] = t[44] ? x[45] : x[44];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[75] | t[52]);
  assign t[55] = ~(t[66]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[113];
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = t[81] | t[114];
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[103] ? x[59] : x[58];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[115];
  assign t[64] = t[103] ? x[64] : x[63];
  assign t[65] = ~(t[116]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[87] | t[67]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[119]);
  assign t[71] = ~(t[120]);
  assign t[72] = ~(t[88] | t[70]);
  assign t[73] = ~(t[89] & t[90]);
  assign t[74] = t[91] | t[121];
  assign t[75] = ~(t[122]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[125]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[93] | t[79]);
  assign t[82] = ~(t[94] & t[95]);
  assign t[83] = t[96] | t[127];
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[97] | t[84]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[98] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[99] | t[94]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [139:0] x;
 output y;

 wire [386:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[2];
  assign t[142] = t[183] ^ x[8];
  assign t[143] = t[184] ^ x[11];
  assign t[144] = t[185] ^ x[14];
  assign t[145] = t[186] ^ x[17];
  assign t[146] = t[187] ^ x[22];
  assign t[147] = t[188] ^ x[27];
  assign t[148] = t[189] ^ x[32];
  assign t[149] = t[190] ^ x[35];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[38];
  assign t[151] = t[192] ^ x[43];
  assign t[152] = t[193] ^ x[48];
  assign t[153] = t[194] ^ x[51];
  assign t[154] = t[195] ^ x[54];
  assign t[155] = t[196] ^ x[57];
  assign t[156] = t[197] ^ x[62];
  assign t[157] = t[198] ^ x[67];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[73];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[76];
  assign t[161] = t[202] ^ x[79];
  assign t[162] = t[203] ^ x[82];
  assign t[163] = t[204] ^ x[85];
  assign t[164] = t[205] ^ x[88];
  assign t[165] = t[206] ^ x[91];
  assign t[166] = t[207] ^ x[94];
  assign t[167] = t[208] ^ x[97];
  assign t[168] = t[209] ^ x[100];
  assign t[169] = t[210] ^ x[103];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[106];
  assign t[171] = t[212] ^ x[109];
  assign t[172] = t[213] ^ x[112];
  assign t[173] = t[214] ^ x[115];
  assign t[174] = t[215] ^ x[118];
  assign t[175] = t[216] ^ x[121];
  assign t[176] = t[217] ^ x[124];
  assign t[177] = t[218] ^ x[127];
  assign t[178] = t[219] ^ x[130];
  assign t[179] = t[220] ^ x[133];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[136];
  assign t[181] = t[222] ^ x[139];
  assign t[182] = (t[223] & ~t[224]);
  assign t[183] = (t[225] & ~t[226]);
  assign t[184] = (t[227] & ~t[228]);
  assign t[185] = (t[229] & ~t[230]);
  assign t[186] = (t[231] & ~t[232]);
  assign t[187] = (t[233] & ~t[234]);
  assign t[188] = (t[235] & ~t[236]);
  assign t[189] = (t[237] & ~t[238]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[239] & ~t[240]);
  assign t[191] = (t[241] & ~t[242]);
  assign t[192] = (t[243] & ~t[244]);
  assign t[193] = (t[245] & ~t[246]);
  assign t[194] = (t[247] & ~t[248]);
  assign t[195] = (t[249] & ~t[250]);
  assign t[196] = (t[251] & ~t[252]);
  assign t[197] = (t[253] & ~t[254]);
  assign t[198] = (t[255] & ~t[256]);
  assign t[199] = (t[257] & ~t[258]);
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[259] & ~t[260]);
  assign t[201] = (t[261] & ~t[262]);
  assign t[202] = (t[263] & ~t[264]);
  assign t[203] = (t[265] & ~t[266]);
  assign t[204] = (t[267] & ~t[268]);
  assign t[205] = (t[269] & ~t[270]);
  assign t[206] = (t[271] & ~t[272]);
  assign t[207] = (t[273] & ~t[274]);
  assign t[208] = (t[275] & ~t[276]);
  assign t[209] = (t[277] & ~t[278]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = (t[279] & ~t[280]);
  assign t[211] = (t[281] & ~t[282]);
  assign t[212] = (t[283] & ~t[284]);
  assign t[213] = (t[285] & ~t[286]);
  assign t[214] = (t[287] & ~t[288]);
  assign t[215] = (t[289] & ~t[290]);
  assign t[216] = (t[291] & ~t[292]);
  assign t[217] = (t[293] & ~t[294]);
  assign t[218] = (t[295] & ~t[296]);
  assign t[219] = (t[297] & ~t[298]);
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[220] = (t[299] & ~t[300]);
  assign t[221] = (t[301] & ~t[302]);
  assign t[222] = (t[303] & ~t[304]);
  assign t[223] = t[305] ^ x[2];
  assign t[224] = t[306] ^ x[1];
  assign t[225] = t[307] ^ x[8];
  assign t[226] = t[308] ^ x[7];
  assign t[227] = t[309] ^ x[11];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[14];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[17];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[22];
  assign t[234] = t[316] ^ x[21];
  assign t[235] = t[317] ^ x[27];
  assign t[236] = t[318] ^ x[26];
  assign t[237] = t[319] ^ x[32];
  assign t[238] = t[320] ^ x[31];
  assign t[239] = t[321] ^ x[35];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[322] ^ x[34];
  assign t[241] = t[323] ^ x[38];
  assign t[242] = t[324] ^ x[37];
  assign t[243] = t[325] ^ x[43];
  assign t[244] = t[326] ^ x[42];
  assign t[245] = t[327] ^ x[48];
  assign t[246] = t[328] ^ x[47];
  assign t[247] = t[329] ^ x[51];
  assign t[248] = t[330] ^ x[50];
  assign t[249] = t[331] ^ x[54];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[53];
  assign t[251] = t[333] ^ x[57];
  assign t[252] = t[334] ^ x[56];
  assign t[253] = t[335] ^ x[62];
  assign t[254] = t[336] ^ x[61];
  assign t[255] = t[337] ^ x[67];
  assign t[256] = t[338] ^ x[66];
  assign t[257] = t[339] ^ x[70];
  assign t[258] = t[340] ^ x[69];
  assign t[259] = t[341] ^ x[73];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[72];
  assign t[261] = t[343] ^ x[76];
  assign t[262] = t[344] ^ x[75];
  assign t[263] = t[345] ^ x[79];
  assign t[264] = t[346] ^ x[78];
  assign t[265] = t[347] ^ x[82];
  assign t[266] = t[348] ^ x[81];
  assign t[267] = t[349] ^ x[85];
  assign t[268] = t[350] ^ x[84];
  assign t[269] = t[351] ^ x[88];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[87];
  assign t[271] = t[353] ^ x[91];
  assign t[272] = t[354] ^ x[90];
  assign t[273] = t[355] ^ x[94];
  assign t[274] = t[356] ^ x[93];
  assign t[275] = t[357] ^ x[97];
  assign t[276] = t[358] ^ x[96];
  assign t[277] = t[359] ^ x[100];
  assign t[278] = t[360] ^ x[99];
  assign t[279] = t[361] ^ x[103];
  assign t[27] = t[43] | t[105];
  assign t[280] = t[362] ^ x[102];
  assign t[281] = t[363] ^ x[106];
  assign t[282] = t[364] ^ x[105];
  assign t[283] = t[365] ^ x[109];
  assign t[284] = t[366] ^ x[108];
  assign t[285] = t[367] ^ x[112];
  assign t[286] = t[368] ^ x[111];
  assign t[287] = t[369] ^ x[115];
  assign t[288] = t[370] ^ x[114];
  assign t[289] = t[371] ^ x[118];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[117];
  assign t[291] = t[373] ^ x[121];
  assign t[292] = t[374] ^ x[120];
  assign t[293] = t[375] ^ x[124];
  assign t[294] = t[376] ^ x[123];
  assign t[295] = t[377] ^ x[127];
  assign t[296] = t[378] ^ x[126];
  assign t[297] = t[379] ^ x[130];
  assign t[298] = t[380] ^ x[129];
  assign t[299] = t[381] ^ x[133];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[132];
  assign t[301] = t[383] ^ x[136];
  assign t[302] = t[384] ^ x[135];
  assign t[303] = t[385] ^ x[139];
  assign t[304] = t[386] ^ x[138];
  assign t[305] = (x[0]);
  assign t[306] = (x[0]);
  assign t[307] = (x[6]);
  assign t[308] = (x[6]);
  assign t[309] = (x[9]);
  assign t[30] = t[47] ^ t[29];
  assign t[310] = (x[9]);
  assign t[311] = (x[12]);
  assign t[312] = (x[12]);
  assign t[313] = (x[15]);
  assign t[314] = (x[15]);
  assign t[315] = (x[20]);
  assign t[316] = (x[20]);
  assign t[317] = (x[25]);
  assign t[318] = (x[25]);
  assign t[319] = (x[30]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = (x[30]);
  assign t[321] = (x[33]);
  assign t[322] = (x[33]);
  assign t[323] = (x[36]);
  assign t[324] = (x[36]);
  assign t[325] = (x[41]);
  assign t[326] = (x[41]);
  assign t[327] = (x[46]);
  assign t[328] = (x[46]);
  assign t[329] = (x[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[330] = (x[49]);
  assign t[331] = (x[52]);
  assign t[332] = (x[52]);
  assign t[333] = (x[55]);
  assign t[334] = (x[55]);
  assign t[335] = (x[60]);
  assign t[336] = (x[60]);
  assign t[337] = (x[65]);
  assign t[338] = (x[65]);
  assign t[339] = (x[68]);
  assign t[33] = ~(t[52] & t[53]);
  assign t[340] = (x[68]);
  assign t[341] = (x[71]);
  assign t[342] = (x[71]);
  assign t[343] = (x[74]);
  assign t[344] = (x[74]);
  assign t[345] = (x[77]);
  assign t[346] = (x[77]);
  assign t[347] = (x[80]);
  assign t[348] = (x[80]);
  assign t[349] = (x[83]);
  assign t[34] = t[54] | t[106];
  assign t[350] = (x[83]);
  assign t[351] = (x[86]);
  assign t[352] = (x[86]);
  assign t[353] = (x[89]);
  assign t[354] = (x[89]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[98]);
  assign t[35] = t[55] ? x[29] : x[28];
  assign t[360] = (x[98]);
  assign t[361] = (x[101]);
  assign t[362] = (x[101]);
  assign t[363] = (x[104]);
  assign t[364] = (x[104]);
  assign t[365] = (x[107]);
  assign t[366] = (x[107]);
  assign t[367] = (x[110]);
  assign t[368] = (x[110]);
  assign t[369] = (x[113]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[113]);
  assign t[371] = (x[116]);
  assign t[372] = (x[116]);
  assign t[373] = (x[119]);
  assign t[374] = (x[119]);
  assign t[375] = (x[122]);
  assign t[376] = (x[122]);
  assign t[377] = (x[125]);
  assign t[378] = (x[125]);
  assign t[379] = (x[128]);
  assign t[37] = ~(t[58] & t[59]);
  assign t[380] = (x[128]);
  assign t[381] = (x[131]);
  assign t[382] = (x[131]);
  assign t[383] = (x[134]);
  assign t[384] = (x[134]);
  assign t[385] = (x[137]);
  assign t[386] = (x[137]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[62] & t[63]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[64] ^ t[39];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[65] | t[41]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = t[69] | t[109];
  assign t[47] = t[44] ? x[40] : x[39];
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = t[72] | t[110];
  assign t[4] = ~(x[3]);
  assign t[50] = t[44] ? x[45] : x[44];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[75] | t[52]);
  assign t[55] = ~(t[66]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[113];
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = t[81] | t[114];
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[103] ? x[59] : x[58];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[115];
  assign t[64] = t[103] ? x[64] : x[63];
  assign t[65] = ~(t[116]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[87] | t[67]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[119]);
  assign t[71] = ~(t[120]);
  assign t[72] = ~(t[88] | t[70]);
  assign t[73] = ~(t[89] & t[90]);
  assign t[74] = t[91] | t[121];
  assign t[75] = ~(t[122]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[125]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[93] | t[79]);
  assign t[82] = ~(t[94] & t[95]);
  assign t[83] = t[96] | t[127];
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[97] | t[84]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[98] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[99] | t[94]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [151:0] x;
 output y;

 wire [519:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[227] | t[145]);
  assign t[101] = t[146] ? x[79] : x[78];
  assign t[102] = ~(t[147] & t[83]);
  assign t[103] = ~(t[228]);
  assign t[104] = ~(t[229]);
  assign t[105] = ~(t[148] | t[149]);
  assign t[106] = t[146] ? x[87] : x[86];
  assign t[107] = ~(t[150] & t[151]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[152] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = ~(t[158] | t[159]);
  assign t[118] = ~(t[235] | t[160]);
  assign t[119] = t[93] ? x[107] : x[106];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[161] & t[162]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[163] | t[164]);
  assign t[124] = t[208] ? x[115] : x[114];
  assign t[125] = t[165] | t[166];
  assign t[126] = ~(t[167] & t[209]);
  assign t[127] = ~(t[168] & t[169]);
  assign t[128] = ~(t[80] | t[170]);
  assign t[129] = ~(t[80] | t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[168] | t[167];
  assign t[132] = ~(x[4] & t[173]);
  assign t[133] = ~(t[174] & t[169]);
  assign t[134] = t[206] ? t[176] : t[175];
  assign t[135] = ~(t[172] & t[177]);
  assign t[136] = ~(t[238]);
  assign t[137] = ~(t[223] | t[224]);
  assign t[138] = ~(t[208]);
  assign t[139] = ~(t[113]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[80] | t[178]);
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[240]);
  assign t[144] = ~(t[241]);
  assign t[145] = ~(t[179] | t[180]);
  assign t[146] = ~(t[138]);
  assign t[147] = ~(t[165] | t[181]);
  assign t[148] = ~(t[242]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[182]);
  assign t[151] = ~(t[183] & t[184]);
  assign t[152] = ~(t[243]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[80] | t[185]);
  assign t[155] = ~(t[80] | t[186]);
  assign t[156] = ~(t[244]);
  assign t[157] = ~(t[233] | t[234]);
  assign t[158] = ~(t[245]);
  assign t[159] = ~(t[246]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[187] | t[188]);
  assign t[161] = ~(t[165] | t[189]);
  assign t[162] = ~(t[48]);
  assign t[163] = ~(t[247]);
  assign t[164] = ~(t[236] | t[237]);
  assign t[165] = ~(t[135] & t[151]);
  assign t[166] = ~(t[190] & t[191]);
  assign t[167] = x[4] & t[207];
  assign t[168] = ~(x[4] | t[207]);
  assign t[169] = ~(t[209]);
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = t[206] ? t[126] : t[127];
  assign t[171] = t[206] ? t[132] : t[192];
  assign t[172] = ~(t[84] | t[206]);
  assign t[173] = ~(t[207] | t[209]);
  assign t[174] = ~(x[4] | t[193]);
  assign t[175] = ~(t[167] & t[169]);
  assign t[176] = ~(t[168] & t[209]);
  assign t[177] = ~(t[192] & t[194]);
  assign t[178] = t[206] ? t[192] : t[132];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[240] | t[241]);
  assign t[181] = t[140] | t[86];
  assign t[182] = ~(t[195] & t[196]);
  assign t[183] = ~(t[207] | t[169]);
  assign t[184] = t[80] & t[206];
  assign t[185] = t[206] ? t[194] : t[133];
  assign t[186] = t[206] ? t[175] : t[176];
  assign t[187] = ~(t[249]);
  assign t[188] = ~(t[245] | t[246]);
  assign t[189] = ~(t[197] & t[198]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[48] | t[86]);
  assign t[191] = ~(t[129] | t[155]);
  assign t[192] = ~(t[209] & t[174]);
  assign t[193] = ~(t[207]);
  assign t[194] = ~(x[4] & t[183]);
  assign t[195] = ~(t[199] | t[200]);
  assign t[196] = ~(t[84] & t[201]);
  assign t[197] = ~(t[50]);
  assign t[198] = t[84] | t[202];
  assign t[199] = ~(t[84] | t[203]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[80] | t[204]);
  assign t[201] = ~(t[132] & t[192]);
  assign t[202] = t[206] ? t[132] : t[133];
  assign t[203] = t[206] ? t[127] : t[175];
  assign t[204] = t[206] ? t[133] : t[194];
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[208] ? x[6] : x[7];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[295] ^ x[2];
  assign t[251] = t[296] ^ x[10];
  assign t[252] = t[297] ^ x[13];
  assign t[253] = t[298] ^ x[16];
  assign t[254] = t[299] ^ x[19];
  assign t[255] = t[300] ^ x[22];
  assign t[256] = t[301] ^ x[25];
  assign t[257] = t[302] ^ x[28];
  assign t[258] = t[303] ^ x[31];
  assign t[259] = t[304] ^ x[34];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[305] ^ x[39];
  assign t[261] = t[306] ^ x[42];
  assign t[262] = t[307] ^ x[45];
  assign t[263] = t[308] ^ x[48];
  assign t[264] = t[309] ^ x[51];
  assign t[265] = t[310] ^ x[56];
  assign t[266] = t[311] ^ x[59];
  assign t[267] = t[312] ^ x[62];
  assign t[268] = t[313] ^ x[65];
  assign t[269] = t[314] ^ x[68];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[315] ^ x[71];
  assign t[271] = t[316] ^ x[74];
  assign t[272] = t[317] ^ x[77];
  assign t[273] = t[318] ^ x[82];
  assign t[274] = t[319] ^ x[85];
  assign t[275] = t[320] ^ x[90];
  assign t[276] = t[321] ^ x[93];
  assign t[277] = t[322] ^ x[96];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[102];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[325] ^ x[105];
  assign t[281] = t[326] ^ x[110];
  assign t[282] = t[327] ^ x[113];
  assign t[283] = t[328] ^ x[118];
  assign t[284] = t[329] ^ x[121];
  assign t[285] = t[330] ^ x[124];
  assign t[286] = t[331] ^ x[127];
  assign t[287] = t[332] ^ x[130];
  assign t[288] = t[333] ^ x[133];
  assign t[289] = t[334] ^ x[136];
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = t[335] ^ x[139];
  assign t[291] = t[336] ^ x[142];
  assign t[292] = t[337] ^ x[145];
  assign t[293] = t[338] ^ x[148];
  assign t[294] = t[339] ^ x[151];
  assign t[295] = (t[340] & ~t[341]);
  assign t[296] = (t[342] & ~t[343]);
  assign t[297] = (t[344] & ~t[345]);
  assign t[298] = (t[346] & ~t[347]);
  assign t[299] = (t[348] & ~t[349]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[350] & ~t[351]);
  assign t[301] = (t[352] & ~t[353]);
  assign t[302] = (t[354] & ~t[355]);
  assign t[303] = (t[356] & ~t[357]);
  assign t[304] = (t[358] & ~t[359]);
  assign t[305] = (t[360] & ~t[361]);
  assign t[306] = (t[362] & ~t[363]);
  assign t[307] = (t[364] & ~t[365]);
  assign t[308] = (t[366] & ~t[367]);
  assign t[309] = (t[368] & ~t[369]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[310] = (t[370] & ~t[371]);
  assign t[311] = (t[372] & ~t[373]);
  assign t[312] = (t[374] & ~t[375]);
  assign t[313] = (t[376] & ~t[377]);
  assign t[314] = (t[378] & ~t[379]);
  assign t[315] = (t[380] & ~t[381]);
  assign t[316] = (t[382] & ~t[383]);
  assign t[317] = (t[384] & ~t[385]);
  assign t[318] = (t[386] & ~t[387]);
  assign t[319] = (t[388] & ~t[389]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[390] & ~t[391]);
  assign t[321] = (t[392] & ~t[393]);
  assign t[322] = (t[394] & ~t[395]);
  assign t[323] = (t[396] & ~t[397]);
  assign t[324] = (t[398] & ~t[399]);
  assign t[325] = (t[400] & ~t[401]);
  assign t[326] = (t[402] & ~t[403]);
  assign t[327] = (t[404] & ~t[405]);
  assign t[328] = (t[406] & ~t[407]);
  assign t[329] = (t[408] & ~t[409]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[410] & ~t[411]);
  assign t[331] = (t[412] & ~t[413]);
  assign t[332] = (t[414] & ~t[415]);
  assign t[333] = (t[416] & ~t[417]);
  assign t[334] = (t[418] & ~t[419]);
  assign t[335] = (t[420] & ~t[421]);
  assign t[336] = (t[422] & ~t[423]);
  assign t[337] = (t[424] & ~t[425]);
  assign t[338] = (t[426] & ~t[427]);
  assign t[339] = (t[428] & ~t[429]);
  assign t[33] = ~(t[210] | t[54]);
  assign t[340] = t[430] ^ x[2];
  assign t[341] = t[431] ^ x[1];
  assign t[342] = t[432] ^ x[10];
  assign t[343] = t[433] ^ x[9];
  assign t[344] = t[434] ^ x[13];
  assign t[345] = t[435] ^ x[12];
  assign t[346] = t[436] ^ x[16];
  assign t[347] = t[437] ^ x[15];
  assign t[348] = t[438] ^ x[19];
  assign t[349] = t[439] ^ x[18];
  assign t[34] = ~(t[55] | t[56]);
  assign t[350] = t[440] ^ x[22];
  assign t[351] = t[441] ^ x[21];
  assign t[352] = t[442] ^ x[25];
  assign t[353] = t[443] ^ x[24];
  assign t[354] = t[444] ^ x[28];
  assign t[355] = t[445] ^ x[27];
  assign t[356] = t[446] ^ x[31];
  assign t[357] = t[447] ^ x[30];
  assign t[358] = t[448] ^ x[34];
  assign t[359] = t[449] ^ x[33];
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[360] = t[450] ^ x[39];
  assign t[361] = t[451] ^ x[38];
  assign t[362] = t[452] ^ x[42];
  assign t[363] = t[453] ^ x[41];
  assign t[364] = t[454] ^ x[45];
  assign t[365] = t[455] ^ x[44];
  assign t[366] = t[456] ^ x[48];
  assign t[367] = t[457] ^ x[47];
  assign t[368] = t[458] ^ x[51];
  assign t[369] = t[459] ^ x[50];
  assign t[36] = ~(t[59] | t[60]);
  assign t[370] = t[460] ^ x[56];
  assign t[371] = t[461] ^ x[55];
  assign t[372] = t[462] ^ x[59];
  assign t[373] = t[463] ^ x[58];
  assign t[374] = t[464] ^ x[62];
  assign t[375] = t[465] ^ x[61];
  assign t[376] = t[466] ^ x[65];
  assign t[377] = t[467] ^ x[64];
  assign t[378] = t[468] ^ x[68];
  assign t[379] = t[469] ^ x[67];
  assign t[37] = ~(t[61] ^ t[62]);
  assign t[380] = t[470] ^ x[71];
  assign t[381] = t[471] ^ x[70];
  assign t[382] = t[472] ^ x[74];
  assign t[383] = t[473] ^ x[73];
  assign t[384] = t[474] ^ x[77];
  assign t[385] = t[475] ^ x[76];
  assign t[386] = t[476] ^ x[82];
  assign t[387] = t[477] ^ x[81];
  assign t[388] = t[478] ^ x[85];
  assign t[389] = t[479] ^ x[84];
  assign t[38] = ~(t[63] | t[64]);
  assign t[390] = t[480] ^ x[90];
  assign t[391] = t[481] ^ x[89];
  assign t[392] = t[482] ^ x[93];
  assign t[393] = t[483] ^ x[92];
  assign t[394] = t[484] ^ x[96];
  assign t[395] = t[485] ^ x[95];
  assign t[396] = t[486] ^ x[99];
  assign t[397] = t[487] ^ x[98];
  assign t[398] = t[488] ^ x[102];
  assign t[399] = t[489] ^ x[101];
  assign t[39] = ~(t[44] ^ t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[105];
  assign t[401] = t[491] ^ x[104];
  assign t[402] = t[492] ^ x[110];
  assign t[403] = t[493] ^ x[109];
  assign t[404] = t[494] ^ x[113];
  assign t[405] = t[495] ^ x[112];
  assign t[406] = t[496] ^ x[118];
  assign t[407] = t[497] ^ x[117];
  assign t[408] = t[498] ^ x[121];
  assign t[409] = t[499] ^ x[120];
  assign t[40] = ~(t[66] | t[67]);
  assign t[410] = t[500] ^ x[124];
  assign t[411] = t[501] ^ x[123];
  assign t[412] = t[502] ^ x[127];
  assign t[413] = t[503] ^ x[126];
  assign t[414] = t[504] ^ x[130];
  assign t[415] = t[505] ^ x[129];
  assign t[416] = t[506] ^ x[133];
  assign t[417] = t[507] ^ x[132];
  assign t[418] = t[508] ^ x[136];
  assign t[419] = t[509] ^ x[135];
  assign t[41] = ~(t[211] | t[68]);
  assign t[420] = t[510] ^ x[139];
  assign t[421] = t[511] ^ x[138];
  assign t[422] = t[512] ^ x[142];
  assign t[423] = t[513] ^ x[141];
  assign t[424] = t[514] ^ x[145];
  assign t[425] = t[515] ^ x[144];
  assign t[426] = t[516] ^ x[148];
  assign t[427] = t[517] ^ x[147];
  assign t[428] = t[518] ^ x[151];
  assign t[429] = t[519] ^ x[150];
  assign t[42] = ~(t[69] | t[70]);
  assign t[430] = (x[0]);
  assign t[431] = (x[0]);
  assign t[432] = (x[8]);
  assign t[433] = (x[8]);
  assign t[434] = (x[11]);
  assign t[435] = (x[11]);
  assign t[436] = (x[14]);
  assign t[437] = (x[14]);
  assign t[438] = (x[17]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[440] = (x[20]);
  assign t[441] = (x[20]);
  assign t[442] = (x[23]);
  assign t[443] = (x[23]);
  assign t[444] = (x[26]);
  assign t[445] = (x[26]);
  assign t[446] = (x[29]);
  assign t[447] = (x[29]);
  assign t[448] = (x[32]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[450] = (x[37]);
  assign t[451] = (x[37]);
  assign t[452] = (x[40]);
  assign t[453] = (x[40]);
  assign t[454] = (x[43]);
  assign t[455] = (x[43]);
  assign t[456] = (x[46]);
  assign t[457] = (x[46]);
  assign t[458] = (x[49]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[460] = (x[54]);
  assign t[461] = (x[54]);
  assign t[462] = (x[57]);
  assign t[463] = (x[57]);
  assign t[464] = (x[60]);
  assign t[465] = (x[60]);
  assign t[466] = (x[63]);
  assign t[467] = (x[63]);
  assign t[468] = (x[66]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[470] = (x[69]);
  assign t[471] = (x[69]);
  assign t[472] = (x[72]);
  assign t[473] = (x[72]);
  assign t[474] = (x[75]);
  assign t[475] = (x[75]);
  assign t[476] = (x[80]);
  assign t[477] = (x[80]);
  assign t[478] = (x[83]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[46] ^ t[79]);
  assign t[480] = (x[88]);
  assign t[481] = (x[88]);
  assign t[482] = (x[91]);
  assign t[483] = (x[91]);
  assign t[484] = (x[94]);
  assign t[485] = (x[94]);
  assign t[486] = (x[97]);
  assign t[487] = (x[97]);
  assign t[488] = (x[100]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[80] | t[81]);
  assign t[490] = (x[103]);
  assign t[491] = (x[103]);
  assign t[492] = (x[108]);
  assign t[493] = (x[108]);
  assign t[494] = (x[111]);
  assign t[495] = (x[111]);
  assign t[496] = (x[116]);
  assign t[497] = (x[116]);
  assign t[498] = (x[119]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[82] & t[83]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[122]);
  assign t[501] = (x[122]);
  assign t[502] = (x[125]);
  assign t[503] = (x[125]);
  assign t[504] = (x[128]);
  assign t[505] = (x[128]);
  assign t[506] = (x[131]);
  assign t[507] = (x[131]);
  assign t[508] = (x[134]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[84] | t[85]);
  assign t[510] = (x[137]);
  assign t[511] = (x[137]);
  assign t[512] = (x[140]);
  assign t[513] = (x[140]);
  assign t[514] = (x[143]);
  assign t[515] = (x[143]);
  assign t[516] = (x[146]);
  assign t[517] = (x[146]);
  assign t[518] = (x[149]);
  assign t[519] = (x[149]);
  assign t[51] = t[86] | t[87];
  assign t[52] = ~(t[212]);
  assign t[53] = ~(t[213]);
  assign t[54] = ~(t[88] | t[89]);
  assign t[55] = ~(t[90] | t[91]);
  assign t[56] = ~(t[214] | t[92]);
  assign t[57] = t[93] ? x[36] : x[35];
  assign t[58] = ~(t[94] & t[95]);
  assign t[59] = ~(t[96] | t[97]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[215] | t[98]);
  assign t[61] = ~(t[99] | t[100]);
  assign t[62] = ~(t[101] ^ t[102]);
  assign t[63] = ~(t[103] | t[104]);
  assign t[64] = ~(t[216] | t[105]);
  assign t[65] = ~(t[106] ^ t[107]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[218]);
  assign t[68] = ~(t[108] | t[109]);
  assign t[69] = ~(t[110] | t[111]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[219] | t[112]);
  assign t[71] = t[208] ? x[53] : x[52];
  assign t[72] = ~(t[30] & t[113]);
  assign t[73] = ~(t[114] | t[115]);
  assign t[74] = ~(t[220] | t[116]);
  assign t[75] = ~(t[117] | t[118]);
  assign t[76] = ~(t[119] ^ t[120]);
  assign t[77] = ~(t[121] | t[122]);
  assign t[78] = ~(t[221] | t[123]);
  assign t[79] = ~(t[124] ^ t[125]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[84]);
  assign t[81] = t[206] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] & t[131]);
  assign t[84] = ~(t[208]);
  assign t[85] = t[206] ? t[133] : t[132];
  assign t[86] = ~(t[80] | t[134]);
  assign t[87] = ~(t[135]);
  assign t[88] = ~(t[222]);
  assign t[89] = ~(t[212] | t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[138]);
  assign t[94] = ~(t[128]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = ~(t[143] | t[144]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [151:0] x;
 output y;

 wire [519:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[227] | t[145]);
  assign t[101] = t[146] ? x[79] : x[78];
  assign t[102] = ~(t[147] & t[83]);
  assign t[103] = ~(t[228]);
  assign t[104] = ~(t[229]);
  assign t[105] = ~(t[148] | t[149]);
  assign t[106] = t[146] ? x[87] : x[86];
  assign t[107] = ~(t[150] & t[151]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[152] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = ~(t[158] | t[159]);
  assign t[118] = ~(t[235] | t[160]);
  assign t[119] = t[93] ? x[107] : x[106];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[161] & t[162]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[163] | t[164]);
  assign t[124] = t[208] ? x[115] : x[114];
  assign t[125] = t[165] | t[166];
  assign t[126] = ~(t[167] & t[209]);
  assign t[127] = ~(t[168] & t[169]);
  assign t[128] = ~(t[80] | t[170]);
  assign t[129] = ~(t[80] | t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[168] | t[167];
  assign t[132] = ~(x[4] & t[173]);
  assign t[133] = ~(t[174] & t[169]);
  assign t[134] = t[206] ? t[176] : t[175];
  assign t[135] = ~(t[172] & t[177]);
  assign t[136] = ~(t[238]);
  assign t[137] = ~(t[223] | t[224]);
  assign t[138] = ~(t[208]);
  assign t[139] = ~(t[113]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[80] | t[178]);
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[240]);
  assign t[144] = ~(t[241]);
  assign t[145] = ~(t[179] | t[180]);
  assign t[146] = ~(t[138]);
  assign t[147] = ~(t[165] | t[181]);
  assign t[148] = ~(t[242]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[182]);
  assign t[151] = ~(t[183] & t[184]);
  assign t[152] = ~(t[243]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[80] | t[185]);
  assign t[155] = ~(t[80] | t[186]);
  assign t[156] = ~(t[244]);
  assign t[157] = ~(t[233] | t[234]);
  assign t[158] = ~(t[245]);
  assign t[159] = ~(t[246]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[187] | t[188]);
  assign t[161] = ~(t[165] | t[189]);
  assign t[162] = ~(t[48]);
  assign t[163] = ~(t[247]);
  assign t[164] = ~(t[236] | t[237]);
  assign t[165] = ~(t[135] & t[151]);
  assign t[166] = ~(t[190] & t[191]);
  assign t[167] = x[4] & t[207];
  assign t[168] = ~(x[4] | t[207]);
  assign t[169] = ~(t[209]);
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = t[206] ? t[126] : t[127];
  assign t[171] = t[206] ? t[132] : t[192];
  assign t[172] = ~(t[84] | t[206]);
  assign t[173] = ~(t[207] | t[209]);
  assign t[174] = ~(x[4] | t[193]);
  assign t[175] = ~(t[167] & t[169]);
  assign t[176] = ~(t[168] & t[209]);
  assign t[177] = ~(t[192] & t[194]);
  assign t[178] = t[206] ? t[192] : t[132];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[240] | t[241]);
  assign t[181] = t[140] | t[86];
  assign t[182] = ~(t[195] & t[196]);
  assign t[183] = ~(t[207] | t[169]);
  assign t[184] = t[80] & t[206];
  assign t[185] = t[206] ? t[194] : t[133];
  assign t[186] = t[206] ? t[175] : t[176];
  assign t[187] = ~(t[249]);
  assign t[188] = ~(t[245] | t[246]);
  assign t[189] = ~(t[197] & t[198]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[48] | t[86]);
  assign t[191] = ~(t[129] | t[155]);
  assign t[192] = ~(t[209] & t[174]);
  assign t[193] = ~(t[207]);
  assign t[194] = ~(x[4] & t[183]);
  assign t[195] = ~(t[199] | t[200]);
  assign t[196] = ~(t[84] & t[201]);
  assign t[197] = ~(t[50]);
  assign t[198] = t[84] | t[202];
  assign t[199] = ~(t[84] | t[203]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[80] | t[204]);
  assign t[201] = ~(t[132] & t[192]);
  assign t[202] = t[206] ? t[132] : t[133];
  assign t[203] = t[206] ? t[127] : t[175];
  assign t[204] = t[206] ? t[133] : t[194];
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[208] ? x[6] : x[7];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[295] ^ x[2];
  assign t[251] = t[296] ^ x[10];
  assign t[252] = t[297] ^ x[13];
  assign t[253] = t[298] ^ x[16];
  assign t[254] = t[299] ^ x[19];
  assign t[255] = t[300] ^ x[22];
  assign t[256] = t[301] ^ x[25];
  assign t[257] = t[302] ^ x[28];
  assign t[258] = t[303] ^ x[31];
  assign t[259] = t[304] ^ x[34];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[305] ^ x[39];
  assign t[261] = t[306] ^ x[42];
  assign t[262] = t[307] ^ x[45];
  assign t[263] = t[308] ^ x[48];
  assign t[264] = t[309] ^ x[51];
  assign t[265] = t[310] ^ x[56];
  assign t[266] = t[311] ^ x[59];
  assign t[267] = t[312] ^ x[62];
  assign t[268] = t[313] ^ x[65];
  assign t[269] = t[314] ^ x[68];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[315] ^ x[71];
  assign t[271] = t[316] ^ x[74];
  assign t[272] = t[317] ^ x[77];
  assign t[273] = t[318] ^ x[82];
  assign t[274] = t[319] ^ x[85];
  assign t[275] = t[320] ^ x[90];
  assign t[276] = t[321] ^ x[93];
  assign t[277] = t[322] ^ x[96];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[102];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[325] ^ x[105];
  assign t[281] = t[326] ^ x[110];
  assign t[282] = t[327] ^ x[113];
  assign t[283] = t[328] ^ x[118];
  assign t[284] = t[329] ^ x[121];
  assign t[285] = t[330] ^ x[124];
  assign t[286] = t[331] ^ x[127];
  assign t[287] = t[332] ^ x[130];
  assign t[288] = t[333] ^ x[133];
  assign t[289] = t[334] ^ x[136];
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = t[335] ^ x[139];
  assign t[291] = t[336] ^ x[142];
  assign t[292] = t[337] ^ x[145];
  assign t[293] = t[338] ^ x[148];
  assign t[294] = t[339] ^ x[151];
  assign t[295] = (t[340] & ~t[341]);
  assign t[296] = (t[342] & ~t[343]);
  assign t[297] = (t[344] & ~t[345]);
  assign t[298] = (t[346] & ~t[347]);
  assign t[299] = (t[348] & ~t[349]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[350] & ~t[351]);
  assign t[301] = (t[352] & ~t[353]);
  assign t[302] = (t[354] & ~t[355]);
  assign t[303] = (t[356] & ~t[357]);
  assign t[304] = (t[358] & ~t[359]);
  assign t[305] = (t[360] & ~t[361]);
  assign t[306] = (t[362] & ~t[363]);
  assign t[307] = (t[364] & ~t[365]);
  assign t[308] = (t[366] & ~t[367]);
  assign t[309] = (t[368] & ~t[369]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[310] = (t[370] & ~t[371]);
  assign t[311] = (t[372] & ~t[373]);
  assign t[312] = (t[374] & ~t[375]);
  assign t[313] = (t[376] & ~t[377]);
  assign t[314] = (t[378] & ~t[379]);
  assign t[315] = (t[380] & ~t[381]);
  assign t[316] = (t[382] & ~t[383]);
  assign t[317] = (t[384] & ~t[385]);
  assign t[318] = (t[386] & ~t[387]);
  assign t[319] = (t[388] & ~t[389]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[390] & ~t[391]);
  assign t[321] = (t[392] & ~t[393]);
  assign t[322] = (t[394] & ~t[395]);
  assign t[323] = (t[396] & ~t[397]);
  assign t[324] = (t[398] & ~t[399]);
  assign t[325] = (t[400] & ~t[401]);
  assign t[326] = (t[402] & ~t[403]);
  assign t[327] = (t[404] & ~t[405]);
  assign t[328] = (t[406] & ~t[407]);
  assign t[329] = (t[408] & ~t[409]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[410] & ~t[411]);
  assign t[331] = (t[412] & ~t[413]);
  assign t[332] = (t[414] & ~t[415]);
  assign t[333] = (t[416] & ~t[417]);
  assign t[334] = (t[418] & ~t[419]);
  assign t[335] = (t[420] & ~t[421]);
  assign t[336] = (t[422] & ~t[423]);
  assign t[337] = (t[424] & ~t[425]);
  assign t[338] = (t[426] & ~t[427]);
  assign t[339] = (t[428] & ~t[429]);
  assign t[33] = ~(t[210] | t[54]);
  assign t[340] = t[430] ^ x[2];
  assign t[341] = t[431] ^ x[1];
  assign t[342] = t[432] ^ x[10];
  assign t[343] = t[433] ^ x[9];
  assign t[344] = t[434] ^ x[13];
  assign t[345] = t[435] ^ x[12];
  assign t[346] = t[436] ^ x[16];
  assign t[347] = t[437] ^ x[15];
  assign t[348] = t[438] ^ x[19];
  assign t[349] = t[439] ^ x[18];
  assign t[34] = ~(t[55] | t[56]);
  assign t[350] = t[440] ^ x[22];
  assign t[351] = t[441] ^ x[21];
  assign t[352] = t[442] ^ x[25];
  assign t[353] = t[443] ^ x[24];
  assign t[354] = t[444] ^ x[28];
  assign t[355] = t[445] ^ x[27];
  assign t[356] = t[446] ^ x[31];
  assign t[357] = t[447] ^ x[30];
  assign t[358] = t[448] ^ x[34];
  assign t[359] = t[449] ^ x[33];
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[360] = t[450] ^ x[39];
  assign t[361] = t[451] ^ x[38];
  assign t[362] = t[452] ^ x[42];
  assign t[363] = t[453] ^ x[41];
  assign t[364] = t[454] ^ x[45];
  assign t[365] = t[455] ^ x[44];
  assign t[366] = t[456] ^ x[48];
  assign t[367] = t[457] ^ x[47];
  assign t[368] = t[458] ^ x[51];
  assign t[369] = t[459] ^ x[50];
  assign t[36] = ~(t[59] | t[60]);
  assign t[370] = t[460] ^ x[56];
  assign t[371] = t[461] ^ x[55];
  assign t[372] = t[462] ^ x[59];
  assign t[373] = t[463] ^ x[58];
  assign t[374] = t[464] ^ x[62];
  assign t[375] = t[465] ^ x[61];
  assign t[376] = t[466] ^ x[65];
  assign t[377] = t[467] ^ x[64];
  assign t[378] = t[468] ^ x[68];
  assign t[379] = t[469] ^ x[67];
  assign t[37] = ~(t[61] ^ t[62]);
  assign t[380] = t[470] ^ x[71];
  assign t[381] = t[471] ^ x[70];
  assign t[382] = t[472] ^ x[74];
  assign t[383] = t[473] ^ x[73];
  assign t[384] = t[474] ^ x[77];
  assign t[385] = t[475] ^ x[76];
  assign t[386] = t[476] ^ x[82];
  assign t[387] = t[477] ^ x[81];
  assign t[388] = t[478] ^ x[85];
  assign t[389] = t[479] ^ x[84];
  assign t[38] = ~(t[63] | t[64]);
  assign t[390] = t[480] ^ x[90];
  assign t[391] = t[481] ^ x[89];
  assign t[392] = t[482] ^ x[93];
  assign t[393] = t[483] ^ x[92];
  assign t[394] = t[484] ^ x[96];
  assign t[395] = t[485] ^ x[95];
  assign t[396] = t[486] ^ x[99];
  assign t[397] = t[487] ^ x[98];
  assign t[398] = t[488] ^ x[102];
  assign t[399] = t[489] ^ x[101];
  assign t[39] = ~(t[44] ^ t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[105];
  assign t[401] = t[491] ^ x[104];
  assign t[402] = t[492] ^ x[110];
  assign t[403] = t[493] ^ x[109];
  assign t[404] = t[494] ^ x[113];
  assign t[405] = t[495] ^ x[112];
  assign t[406] = t[496] ^ x[118];
  assign t[407] = t[497] ^ x[117];
  assign t[408] = t[498] ^ x[121];
  assign t[409] = t[499] ^ x[120];
  assign t[40] = ~(t[66] | t[67]);
  assign t[410] = t[500] ^ x[124];
  assign t[411] = t[501] ^ x[123];
  assign t[412] = t[502] ^ x[127];
  assign t[413] = t[503] ^ x[126];
  assign t[414] = t[504] ^ x[130];
  assign t[415] = t[505] ^ x[129];
  assign t[416] = t[506] ^ x[133];
  assign t[417] = t[507] ^ x[132];
  assign t[418] = t[508] ^ x[136];
  assign t[419] = t[509] ^ x[135];
  assign t[41] = ~(t[211] | t[68]);
  assign t[420] = t[510] ^ x[139];
  assign t[421] = t[511] ^ x[138];
  assign t[422] = t[512] ^ x[142];
  assign t[423] = t[513] ^ x[141];
  assign t[424] = t[514] ^ x[145];
  assign t[425] = t[515] ^ x[144];
  assign t[426] = t[516] ^ x[148];
  assign t[427] = t[517] ^ x[147];
  assign t[428] = t[518] ^ x[151];
  assign t[429] = t[519] ^ x[150];
  assign t[42] = ~(t[69] | t[70]);
  assign t[430] = (x[0]);
  assign t[431] = (x[0]);
  assign t[432] = (x[8]);
  assign t[433] = (x[8]);
  assign t[434] = (x[11]);
  assign t[435] = (x[11]);
  assign t[436] = (x[14]);
  assign t[437] = (x[14]);
  assign t[438] = (x[17]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[440] = (x[20]);
  assign t[441] = (x[20]);
  assign t[442] = (x[23]);
  assign t[443] = (x[23]);
  assign t[444] = (x[26]);
  assign t[445] = (x[26]);
  assign t[446] = (x[29]);
  assign t[447] = (x[29]);
  assign t[448] = (x[32]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[450] = (x[37]);
  assign t[451] = (x[37]);
  assign t[452] = (x[40]);
  assign t[453] = (x[40]);
  assign t[454] = (x[43]);
  assign t[455] = (x[43]);
  assign t[456] = (x[46]);
  assign t[457] = (x[46]);
  assign t[458] = (x[49]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[460] = (x[54]);
  assign t[461] = (x[54]);
  assign t[462] = (x[57]);
  assign t[463] = (x[57]);
  assign t[464] = (x[60]);
  assign t[465] = (x[60]);
  assign t[466] = (x[63]);
  assign t[467] = (x[63]);
  assign t[468] = (x[66]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[470] = (x[69]);
  assign t[471] = (x[69]);
  assign t[472] = (x[72]);
  assign t[473] = (x[72]);
  assign t[474] = (x[75]);
  assign t[475] = (x[75]);
  assign t[476] = (x[80]);
  assign t[477] = (x[80]);
  assign t[478] = (x[83]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[46] ^ t[79]);
  assign t[480] = (x[88]);
  assign t[481] = (x[88]);
  assign t[482] = (x[91]);
  assign t[483] = (x[91]);
  assign t[484] = (x[94]);
  assign t[485] = (x[94]);
  assign t[486] = (x[97]);
  assign t[487] = (x[97]);
  assign t[488] = (x[100]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[80] | t[81]);
  assign t[490] = (x[103]);
  assign t[491] = (x[103]);
  assign t[492] = (x[108]);
  assign t[493] = (x[108]);
  assign t[494] = (x[111]);
  assign t[495] = (x[111]);
  assign t[496] = (x[116]);
  assign t[497] = (x[116]);
  assign t[498] = (x[119]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[82] & t[83]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[122]);
  assign t[501] = (x[122]);
  assign t[502] = (x[125]);
  assign t[503] = (x[125]);
  assign t[504] = (x[128]);
  assign t[505] = (x[128]);
  assign t[506] = (x[131]);
  assign t[507] = (x[131]);
  assign t[508] = (x[134]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[84] | t[85]);
  assign t[510] = (x[137]);
  assign t[511] = (x[137]);
  assign t[512] = (x[140]);
  assign t[513] = (x[140]);
  assign t[514] = (x[143]);
  assign t[515] = (x[143]);
  assign t[516] = (x[146]);
  assign t[517] = (x[146]);
  assign t[518] = (x[149]);
  assign t[519] = (x[149]);
  assign t[51] = t[86] | t[87];
  assign t[52] = ~(t[212]);
  assign t[53] = ~(t[213]);
  assign t[54] = ~(t[88] | t[89]);
  assign t[55] = ~(t[90] | t[91]);
  assign t[56] = ~(t[214] | t[92]);
  assign t[57] = t[93] ? x[36] : x[35];
  assign t[58] = ~(t[94] & t[95]);
  assign t[59] = ~(t[96] | t[97]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[215] | t[98]);
  assign t[61] = ~(t[99] | t[100]);
  assign t[62] = ~(t[101] ^ t[102]);
  assign t[63] = ~(t[103] | t[104]);
  assign t[64] = ~(t[216] | t[105]);
  assign t[65] = ~(t[106] ^ t[107]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[218]);
  assign t[68] = ~(t[108] | t[109]);
  assign t[69] = ~(t[110] | t[111]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[219] | t[112]);
  assign t[71] = t[208] ? x[53] : x[52];
  assign t[72] = ~(t[30] & t[113]);
  assign t[73] = ~(t[114] | t[115]);
  assign t[74] = ~(t[220] | t[116]);
  assign t[75] = ~(t[117] | t[118]);
  assign t[76] = ~(t[119] ^ t[120]);
  assign t[77] = ~(t[121] | t[122]);
  assign t[78] = ~(t[221] | t[123]);
  assign t[79] = ~(t[124] ^ t[125]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[84]);
  assign t[81] = t[206] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] & t[131]);
  assign t[84] = ~(t[208]);
  assign t[85] = t[206] ? t[133] : t[132];
  assign t[86] = ~(t[80] | t[134]);
  assign t[87] = ~(t[135]);
  assign t[88] = ~(t[222]);
  assign t[89] = ~(t[212] | t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[138]);
  assign t[94] = ~(t[128]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = ~(t[143] | t[144]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [121:0] x;
 output y;

 wire [342:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[18] : x[19];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[2];
  assign t[134] = t[169] ^ x[8];
  assign t[135] = t[170] ^ x[11];
  assign t[136] = t[171] ^ x[14];
  assign t[137] = t[172] ^ x[17];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[25];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[30];
  assign t[141] = t[176] ^ x[33];
  assign t[142] = t[177] ^ x[38];
  assign t[143] = t[178] ^ x[41];
  assign t[144] = t[179] ^ x[44];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[50];
  assign t[147] = t[182] ^ x[55];
  assign t[148] = t[183] ^ x[58];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[66];
  assign t[151] = t[186] ^ x[69];
  assign t[152] = t[187] ^ x[72];
  assign t[153] = t[188] ^ x[75];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[83];
  assign t[156] = t[191] ^ x[88];
  assign t[157] = t[192] ^ x[91];
  assign t[158] = t[193] ^ x[94];
  assign t[159] = t[194] ^ x[97];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[106];
  assign t[163] = t[198] ^ x[109];
  assign t[164] = t[199] ^ x[112];
  assign t[165] = t[200] ^ x[115];
  assign t[166] = t[201] ^ x[118];
  assign t[167] = t[202] ^ x[121];
  assign t[168] = (t[203] & ~t[204]);
  assign t[169] = (t[205] & ~t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (t[207] & ~t[208]);
  assign t[171] = (t[209] & ~t[210]);
  assign t[172] = (t[211] & ~t[212]);
  assign t[173] = (t[213] & ~t[214]);
  assign t[174] = (t[215] & ~t[216]);
  assign t[175] = (t[217] & ~t[218]);
  assign t[176] = (t[219] & ~t[220]);
  assign t[177] = (t[221] & ~t[222]);
  assign t[178] = (t[223] & ~t[224]);
  assign t[179] = (t[225] & ~t[226]);
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = (t[227] & ~t[228]);
  assign t[181] = (t[229] & ~t[230]);
  assign t[182] = (t[231] & ~t[232]);
  assign t[183] = (t[233] & ~t[234]);
  assign t[184] = (t[235] & ~t[236]);
  assign t[185] = (t[237] & ~t[238]);
  assign t[186] = (t[239] & ~t[240]);
  assign t[187] = (t[241] & ~t[242]);
  assign t[188] = (t[243] & ~t[244]);
  assign t[189] = (t[245] & ~t[246]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (t[247] & ~t[248]);
  assign t[191] = (t[249] & ~t[250]);
  assign t[192] = (t[251] & ~t[252]);
  assign t[193] = (t[253] & ~t[254]);
  assign t[194] = (t[255] & ~t[256]);
  assign t[195] = (t[257] & ~t[258]);
  assign t[196] = (t[259] & ~t[260]);
  assign t[197] = (t[261] & ~t[262]);
  assign t[198] = (t[263] & ~t[264]);
  assign t[199] = (t[265] & ~t[266]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[267] & ~t[268]);
  assign t[201] = (t[269] & ~t[270]);
  assign t[202] = (t[271] & ~t[272]);
  assign t[203] = t[273] ^ x[2];
  assign t[204] = t[274] ^ x[1];
  assign t[205] = t[275] ^ x[8];
  assign t[206] = t[276] ^ x[7];
  assign t[207] = t[277] ^ x[11];
  assign t[208] = t[278] ^ x[10];
  assign t[209] = t[279] ^ x[14];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[280] ^ x[13];
  assign t[211] = t[281] ^ x[17];
  assign t[212] = t[282] ^ x[16];
  assign t[213] = t[283] ^ x[22];
  assign t[214] = t[284] ^ x[21];
  assign t[215] = t[285] ^ x[25];
  assign t[216] = t[286] ^ x[24];
  assign t[217] = t[287] ^ x[30];
  assign t[218] = t[288] ^ x[29];
  assign t[219] = t[289] ^ x[33];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[290] ^ x[32];
  assign t[221] = t[291] ^ x[38];
  assign t[222] = t[292] ^ x[37];
  assign t[223] = t[293] ^ x[41];
  assign t[224] = t[294] ^ x[40];
  assign t[225] = t[295] ^ x[44];
  assign t[226] = t[296] ^ x[43];
  assign t[227] = t[297] ^ x[47];
  assign t[228] = t[298] ^ x[46];
  assign t[229] = t[299] ^ x[50];
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = t[300] ^ x[49];
  assign t[231] = t[301] ^ x[55];
  assign t[232] = t[302] ^ x[54];
  assign t[233] = t[303] ^ x[58];
  assign t[234] = t[304] ^ x[57];
  assign t[235] = t[305] ^ x[63];
  assign t[236] = t[306] ^ x[62];
  assign t[237] = t[307] ^ x[66];
  assign t[238] = t[308] ^ x[65];
  assign t[239] = t[309] ^ x[69];
  assign t[23] = ~(t[101]);
  assign t[240] = t[310] ^ x[68];
  assign t[241] = t[311] ^ x[72];
  assign t[242] = t[312] ^ x[71];
  assign t[243] = t[313] ^ x[75];
  assign t[244] = t[314] ^ x[74];
  assign t[245] = t[315] ^ x[80];
  assign t[246] = t[316] ^ x[79];
  assign t[247] = t[317] ^ x[83];
  assign t[248] = t[318] ^ x[82];
  assign t[249] = t[319] ^ x[88];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[320] ^ x[87];
  assign t[251] = t[321] ^ x[91];
  assign t[252] = t[322] ^ x[90];
  assign t[253] = t[323] ^ x[94];
  assign t[254] = t[324] ^ x[93];
  assign t[255] = t[325] ^ x[97];
  assign t[256] = t[326] ^ x[96];
  assign t[257] = t[327] ^ x[100];
  assign t[258] = t[328] ^ x[99];
  assign t[259] = t[329] ^ x[103];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[330] ^ x[102];
  assign t[261] = t[331] ^ x[106];
  assign t[262] = t[332] ^ x[105];
  assign t[263] = t[333] ^ x[109];
  assign t[264] = t[334] ^ x[108];
  assign t[265] = t[335] ^ x[112];
  assign t[266] = t[336] ^ x[111];
  assign t[267] = t[337] ^ x[115];
  assign t[268] = t[338] ^ x[114];
  assign t[269] = t[339] ^ x[118];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[340] ^ x[117];
  assign t[271] = t[341] ^ x[121];
  assign t[272] = t[342] ^ x[120];
  assign t[273] = (x[0]);
  assign t[274] = (x[0]);
  assign t[275] = (x[6]);
  assign t[276] = (x[6]);
  assign t[277] = (x[9]);
  assign t[278] = (x[9]);
  assign t[279] = (x[12]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[12]);
  assign t[281] = (x[15]);
  assign t[282] = (x[15]);
  assign t[283] = (x[20]);
  assign t[284] = (x[20]);
  assign t[285] = (x[23]);
  assign t[286] = (x[23]);
  assign t[287] = (x[28]);
  assign t[288] = (x[28]);
  assign t[289] = (x[31]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[31]);
  assign t[291] = (x[36]);
  assign t[292] = (x[36]);
  assign t[293] = (x[39]);
  assign t[294] = (x[39]);
  assign t[295] = (x[42]);
  assign t[296] = (x[42]);
  assign t[297] = (x[45]);
  assign t[298] = (x[45]);
  assign t[299] = (x[48]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[48]);
  assign t[301] = (x[53]);
  assign t[302] = (x[53]);
  assign t[303] = (x[56]);
  assign t[304] = (x[56]);
  assign t[305] = (x[61]);
  assign t[306] = (x[61]);
  assign t[307] = (x[64]);
  assign t[308] = (x[64]);
  assign t[309] = (x[67]);
  assign t[30] = t[46] ? x[27] : x[26];
  assign t[310] = (x[67]);
  assign t[311] = (x[70]);
  assign t[312] = (x[70]);
  assign t[313] = (x[73]);
  assign t[314] = (x[73]);
  assign t[315] = (x[78]);
  assign t[316] = (x[78]);
  assign t[317] = (x[81]);
  assign t[318] = (x[81]);
  assign t[319] = (x[86]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[86]);
  assign t[321] = (x[89]);
  assign t[322] = (x[89]);
  assign t[323] = (x[92]);
  assign t[324] = (x[92]);
  assign t[325] = (x[95]);
  assign t[326] = (x[95]);
  assign t[327] = (x[98]);
  assign t[328] = (x[98]);
  assign t[329] = (x[101]);
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = (x[101]);
  assign t[331] = (x[104]);
  assign t[332] = (x[104]);
  assign t[333] = (x[107]);
  assign t[334] = (x[107]);
  assign t[335] = (x[110]);
  assign t[336] = (x[110]);
  assign t[337] = (x[113]);
  assign t[338] = (x[113]);
  assign t[339] = (x[116]);
  assign t[33] = t[51] ^ t[42];
  assign t[340] = (x[116]);
  assign t[341] = (x[119]);
  assign t[342] = (x[119]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[35] = t[54] ^ t[55];
  assign t[36] = ~(t[105] & t[56]);
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = t[101] ? x[35] : x[34];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[67]);
  assign t[46] = ~(t[23]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = t[72] ? x[52] : x[51];
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = t[72] ? x[60] : x[59];
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = t[101] ? x[77] : x[76];
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[101] ? x[85] : x[84];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[103]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[23]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[131]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[131] & t[96]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[124]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind151(x, y);
 input [121:0] x;
 output y;

 wire [342:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[18] : x[19];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[2];
  assign t[134] = t[169] ^ x[8];
  assign t[135] = t[170] ^ x[11];
  assign t[136] = t[171] ^ x[14];
  assign t[137] = t[172] ^ x[17];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[25];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[30];
  assign t[141] = t[176] ^ x[33];
  assign t[142] = t[177] ^ x[38];
  assign t[143] = t[178] ^ x[41];
  assign t[144] = t[179] ^ x[44];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[50];
  assign t[147] = t[182] ^ x[55];
  assign t[148] = t[183] ^ x[58];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[66];
  assign t[151] = t[186] ^ x[69];
  assign t[152] = t[187] ^ x[72];
  assign t[153] = t[188] ^ x[75];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[83];
  assign t[156] = t[191] ^ x[88];
  assign t[157] = t[192] ^ x[91];
  assign t[158] = t[193] ^ x[94];
  assign t[159] = t[194] ^ x[97];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[106];
  assign t[163] = t[198] ^ x[109];
  assign t[164] = t[199] ^ x[112];
  assign t[165] = t[200] ^ x[115];
  assign t[166] = t[201] ^ x[118];
  assign t[167] = t[202] ^ x[121];
  assign t[168] = (t[203] & ~t[204]);
  assign t[169] = (t[205] & ~t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (t[207] & ~t[208]);
  assign t[171] = (t[209] & ~t[210]);
  assign t[172] = (t[211] & ~t[212]);
  assign t[173] = (t[213] & ~t[214]);
  assign t[174] = (t[215] & ~t[216]);
  assign t[175] = (t[217] & ~t[218]);
  assign t[176] = (t[219] & ~t[220]);
  assign t[177] = (t[221] & ~t[222]);
  assign t[178] = (t[223] & ~t[224]);
  assign t[179] = (t[225] & ~t[226]);
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = (t[227] & ~t[228]);
  assign t[181] = (t[229] & ~t[230]);
  assign t[182] = (t[231] & ~t[232]);
  assign t[183] = (t[233] & ~t[234]);
  assign t[184] = (t[235] & ~t[236]);
  assign t[185] = (t[237] & ~t[238]);
  assign t[186] = (t[239] & ~t[240]);
  assign t[187] = (t[241] & ~t[242]);
  assign t[188] = (t[243] & ~t[244]);
  assign t[189] = (t[245] & ~t[246]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (t[247] & ~t[248]);
  assign t[191] = (t[249] & ~t[250]);
  assign t[192] = (t[251] & ~t[252]);
  assign t[193] = (t[253] & ~t[254]);
  assign t[194] = (t[255] & ~t[256]);
  assign t[195] = (t[257] & ~t[258]);
  assign t[196] = (t[259] & ~t[260]);
  assign t[197] = (t[261] & ~t[262]);
  assign t[198] = (t[263] & ~t[264]);
  assign t[199] = (t[265] & ~t[266]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[267] & ~t[268]);
  assign t[201] = (t[269] & ~t[270]);
  assign t[202] = (t[271] & ~t[272]);
  assign t[203] = t[273] ^ x[2];
  assign t[204] = t[274] ^ x[1];
  assign t[205] = t[275] ^ x[8];
  assign t[206] = t[276] ^ x[7];
  assign t[207] = t[277] ^ x[11];
  assign t[208] = t[278] ^ x[10];
  assign t[209] = t[279] ^ x[14];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[280] ^ x[13];
  assign t[211] = t[281] ^ x[17];
  assign t[212] = t[282] ^ x[16];
  assign t[213] = t[283] ^ x[22];
  assign t[214] = t[284] ^ x[21];
  assign t[215] = t[285] ^ x[25];
  assign t[216] = t[286] ^ x[24];
  assign t[217] = t[287] ^ x[30];
  assign t[218] = t[288] ^ x[29];
  assign t[219] = t[289] ^ x[33];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[290] ^ x[32];
  assign t[221] = t[291] ^ x[38];
  assign t[222] = t[292] ^ x[37];
  assign t[223] = t[293] ^ x[41];
  assign t[224] = t[294] ^ x[40];
  assign t[225] = t[295] ^ x[44];
  assign t[226] = t[296] ^ x[43];
  assign t[227] = t[297] ^ x[47];
  assign t[228] = t[298] ^ x[46];
  assign t[229] = t[299] ^ x[50];
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = t[300] ^ x[49];
  assign t[231] = t[301] ^ x[55];
  assign t[232] = t[302] ^ x[54];
  assign t[233] = t[303] ^ x[58];
  assign t[234] = t[304] ^ x[57];
  assign t[235] = t[305] ^ x[63];
  assign t[236] = t[306] ^ x[62];
  assign t[237] = t[307] ^ x[66];
  assign t[238] = t[308] ^ x[65];
  assign t[239] = t[309] ^ x[69];
  assign t[23] = ~(t[101]);
  assign t[240] = t[310] ^ x[68];
  assign t[241] = t[311] ^ x[72];
  assign t[242] = t[312] ^ x[71];
  assign t[243] = t[313] ^ x[75];
  assign t[244] = t[314] ^ x[74];
  assign t[245] = t[315] ^ x[80];
  assign t[246] = t[316] ^ x[79];
  assign t[247] = t[317] ^ x[83];
  assign t[248] = t[318] ^ x[82];
  assign t[249] = t[319] ^ x[88];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[320] ^ x[87];
  assign t[251] = t[321] ^ x[91];
  assign t[252] = t[322] ^ x[90];
  assign t[253] = t[323] ^ x[94];
  assign t[254] = t[324] ^ x[93];
  assign t[255] = t[325] ^ x[97];
  assign t[256] = t[326] ^ x[96];
  assign t[257] = t[327] ^ x[100];
  assign t[258] = t[328] ^ x[99];
  assign t[259] = t[329] ^ x[103];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[330] ^ x[102];
  assign t[261] = t[331] ^ x[106];
  assign t[262] = t[332] ^ x[105];
  assign t[263] = t[333] ^ x[109];
  assign t[264] = t[334] ^ x[108];
  assign t[265] = t[335] ^ x[112];
  assign t[266] = t[336] ^ x[111];
  assign t[267] = t[337] ^ x[115];
  assign t[268] = t[338] ^ x[114];
  assign t[269] = t[339] ^ x[118];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[340] ^ x[117];
  assign t[271] = t[341] ^ x[121];
  assign t[272] = t[342] ^ x[120];
  assign t[273] = (x[0]);
  assign t[274] = (x[0]);
  assign t[275] = (x[6]);
  assign t[276] = (x[6]);
  assign t[277] = (x[9]);
  assign t[278] = (x[9]);
  assign t[279] = (x[12]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[12]);
  assign t[281] = (x[15]);
  assign t[282] = (x[15]);
  assign t[283] = (x[20]);
  assign t[284] = (x[20]);
  assign t[285] = (x[23]);
  assign t[286] = (x[23]);
  assign t[287] = (x[28]);
  assign t[288] = (x[28]);
  assign t[289] = (x[31]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[31]);
  assign t[291] = (x[36]);
  assign t[292] = (x[36]);
  assign t[293] = (x[39]);
  assign t[294] = (x[39]);
  assign t[295] = (x[42]);
  assign t[296] = (x[42]);
  assign t[297] = (x[45]);
  assign t[298] = (x[45]);
  assign t[299] = (x[48]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[48]);
  assign t[301] = (x[53]);
  assign t[302] = (x[53]);
  assign t[303] = (x[56]);
  assign t[304] = (x[56]);
  assign t[305] = (x[61]);
  assign t[306] = (x[61]);
  assign t[307] = (x[64]);
  assign t[308] = (x[64]);
  assign t[309] = (x[67]);
  assign t[30] = t[46] ? x[27] : x[26];
  assign t[310] = (x[67]);
  assign t[311] = (x[70]);
  assign t[312] = (x[70]);
  assign t[313] = (x[73]);
  assign t[314] = (x[73]);
  assign t[315] = (x[78]);
  assign t[316] = (x[78]);
  assign t[317] = (x[81]);
  assign t[318] = (x[81]);
  assign t[319] = (x[86]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[86]);
  assign t[321] = (x[89]);
  assign t[322] = (x[89]);
  assign t[323] = (x[92]);
  assign t[324] = (x[92]);
  assign t[325] = (x[95]);
  assign t[326] = (x[95]);
  assign t[327] = (x[98]);
  assign t[328] = (x[98]);
  assign t[329] = (x[101]);
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = (x[101]);
  assign t[331] = (x[104]);
  assign t[332] = (x[104]);
  assign t[333] = (x[107]);
  assign t[334] = (x[107]);
  assign t[335] = (x[110]);
  assign t[336] = (x[110]);
  assign t[337] = (x[113]);
  assign t[338] = (x[113]);
  assign t[339] = (x[116]);
  assign t[33] = t[51] ^ t[42];
  assign t[340] = (x[116]);
  assign t[341] = (x[119]);
  assign t[342] = (x[119]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[35] = t[54] ^ t[55];
  assign t[36] = ~(t[105] & t[56]);
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = t[101] ? x[35] : x[34];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[67]);
  assign t[46] = ~(t[23]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = t[72] ? x[52] : x[51];
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = t[72] ? x[60] : x[59];
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = t[101] ? x[77] : x[76];
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[101] ? x[85] : x[84];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[103]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[23]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[131]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[131] & t[96]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[124]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [151:0] x;
 output y;

 wire [431:0] t;
  assign t[0] = t[1] ? t[2] : t[117];
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[113] & t[114]);
  assign t[104] = ~(t[144] & t[143]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[156]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[115] & t[116]);
  assign t[111] = ~(t[149] & t[148]);
  assign t[112] = ~(t[159]);
  assign t[113] = ~(t[154] & t[153]);
  assign t[114] = ~(t[160]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[18] : x[19];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = t[207] ^ x[2];
  assign t[163] = t[208] ^ x[8];
  assign t[164] = t[209] ^ x[11];
  assign t[165] = t[210] ^ x[14];
  assign t[166] = t[211] ^ x[17];
  assign t[167] = t[212] ^ x[22];
  assign t[168] = t[213] ^ x[27];
  assign t[169] = t[214] ^ x[32];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[35];
  assign t[171] = t[216] ^ x[38];
  assign t[172] = t[217] ^ x[41];
  assign t[173] = t[218] ^ x[46];
  assign t[174] = t[219] ^ x[51];
  assign t[175] = t[220] ^ x[54];
  assign t[176] = t[221] ^ x[57];
  assign t[177] = t[222] ^ x[60];
  assign t[178] = t[223] ^ x[65];
  assign t[179] = t[224] ^ x[70];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[73];
  assign t[181] = t[226] ^ x[76];
  assign t[182] = t[227] ^ x[79];
  assign t[183] = t[228] ^ x[82];
  assign t[184] = t[229] ^ x[85];
  assign t[185] = t[230] ^ x[88];
  assign t[186] = t[231] ^ x[91];
  assign t[187] = t[232] ^ x[94];
  assign t[188] = t[233] ^ x[97];
  assign t[189] = t[234] ^ x[100];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[103];
  assign t[191] = t[236] ^ x[106];
  assign t[192] = t[237] ^ x[109];
  assign t[193] = t[238] ^ x[112];
  assign t[194] = t[239] ^ x[115];
  assign t[195] = t[240] ^ x[118];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[124];
  assign t[198] = t[243] ^ x[127];
  assign t[199] = t[244] ^ x[130];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[133];
  assign t[201] = t[246] ^ x[136];
  assign t[202] = t[247] ^ x[139];
  assign t[203] = t[248] ^ x[142];
  assign t[204] = t[249] ^ x[145];
  assign t[205] = t[250] ^ x[148];
  assign t[206] = t[251] ^ x[151];
  assign t[207] = (t[252] & ~t[253]);
  assign t[208] = (t[254] & ~t[255]);
  assign t[209] = (t[256] & ~t[257]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[258] & ~t[259]);
  assign t[211] = (t[260] & ~t[261]);
  assign t[212] = (t[262] & ~t[263]);
  assign t[213] = (t[264] & ~t[265]);
  assign t[214] = (t[266] & ~t[267]);
  assign t[215] = (t[268] & ~t[269]);
  assign t[216] = (t[270] & ~t[271]);
  assign t[217] = (t[272] & ~t[273]);
  assign t[218] = (t[274] & ~t[275]);
  assign t[219] = (t[276] & ~t[277]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[278] & ~t[279]);
  assign t[221] = (t[280] & ~t[281]);
  assign t[222] = (t[282] & ~t[283]);
  assign t[223] = (t[284] & ~t[285]);
  assign t[224] = (t[286] & ~t[287]);
  assign t[225] = (t[288] & ~t[289]);
  assign t[226] = (t[290] & ~t[291]);
  assign t[227] = (t[292] & ~t[293]);
  assign t[228] = (t[294] & ~t[295]);
  assign t[229] = (t[296] & ~t[297]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[298] & ~t[299]);
  assign t[231] = (t[300] & ~t[301]);
  assign t[232] = (t[302] & ~t[303]);
  assign t[233] = (t[304] & ~t[305]);
  assign t[234] = (t[306] & ~t[307]);
  assign t[235] = (t[308] & ~t[309]);
  assign t[236] = (t[310] & ~t[311]);
  assign t[237] = (t[312] & ~t[313]);
  assign t[238] = (t[314] & ~t[315]);
  assign t[239] = (t[316] & ~t[317]);
  assign t[23] = ~(t[120]);
  assign t[240] = (t[318] & ~t[319]);
  assign t[241] = (t[320] & ~t[321]);
  assign t[242] = (t[322] & ~t[323]);
  assign t[243] = (t[324] & ~t[325]);
  assign t[244] = (t[326] & ~t[327]);
  assign t[245] = (t[328] & ~t[329]);
  assign t[246] = (t[330] & ~t[331]);
  assign t[247] = (t[332] & ~t[333]);
  assign t[248] = (t[334] & ~t[335]);
  assign t[249] = (t[336] & ~t[337]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (t[338] & ~t[339]);
  assign t[251] = (t[340] & ~t[341]);
  assign t[252] = t[342] ^ x[2];
  assign t[253] = t[343] ^ x[1];
  assign t[254] = t[344] ^ x[8];
  assign t[255] = t[345] ^ x[7];
  assign t[256] = t[346] ^ x[11];
  assign t[257] = t[347] ^ x[10];
  assign t[258] = t[348] ^ x[14];
  assign t[259] = t[349] ^ x[13];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[17];
  assign t[261] = t[351] ^ x[16];
  assign t[262] = t[352] ^ x[22];
  assign t[263] = t[353] ^ x[21];
  assign t[264] = t[354] ^ x[27];
  assign t[265] = t[355] ^ x[26];
  assign t[266] = t[356] ^ x[32];
  assign t[267] = t[357] ^ x[31];
  assign t[268] = t[358] ^ x[35];
  assign t[269] = t[359] ^ x[34];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[38];
  assign t[271] = t[361] ^ x[37];
  assign t[272] = t[362] ^ x[41];
  assign t[273] = t[363] ^ x[40];
  assign t[274] = t[364] ^ x[46];
  assign t[275] = t[365] ^ x[45];
  assign t[276] = t[366] ^ x[51];
  assign t[277] = t[367] ^ x[50];
  assign t[278] = t[368] ^ x[54];
  assign t[279] = t[369] ^ x[53];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[57];
  assign t[281] = t[371] ^ x[56];
  assign t[282] = t[372] ^ x[60];
  assign t[283] = t[373] ^ x[59];
  assign t[284] = t[374] ^ x[65];
  assign t[285] = t[375] ^ x[64];
  assign t[286] = t[376] ^ x[70];
  assign t[287] = t[377] ^ x[69];
  assign t[288] = t[378] ^ x[73];
  assign t[289] = t[379] ^ x[72];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[76];
  assign t[291] = t[381] ^ x[75];
  assign t[292] = t[382] ^ x[79];
  assign t[293] = t[383] ^ x[78];
  assign t[294] = t[384] ^ x[82];
  assign t[295] = t[385] ^ x[81];
  assign t[296] = t[386] ^ x[85];
  assign t[297] = t[387] ^ x[84];
  assign t[298] = t[388] ^ x[88];
  assign t[299] = t[389] ^ x[87];
  assign t[29] = ~(t[46] & t[122]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[91];
  assign t[301] = t[391] ^ x[90];
  assign t[302] = t[392] ^ x[94];
  assign t[303] = t[393] ^ x[93];
  assign t[304] = t[394] ^ x[97];
  assign t[305] = t[395] ^ x[96];
  assign t[306] = t[396] ^ x[100];
  assign t[307] = t[397] ^ x[99];
  assign t[308] = t[398] ^ x[103];
  assign t[309] = t[399] ^ x[102];
  assign t[30] = t[47] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[106];
  assign t[311] = t[401] ^ x[105];
  assign t[312] = t[402] ^ x[109];
  assign t[313] = t[403] ^ x[108];
  assign t[314] = t[404] ^ x[112];
  assign t[315] = t[405] ^ x[111];
  assign t[316] = t[406] ^ x[115];
  assign t[317] = t[407] ^ x[114];
  assign t[318] = t[408] ^ x[118];
  assign t[319] = t[409] ^ x[117];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[410] ^ x[121];
  assign t[321] = t[411] ^ x[120];
  assign t[322] = t[412] ^ x[124];
  assign t[323] = t[413] ^ x[123];
  assign t[324] = t[414] ^ x[127];
  assign t[325] = t[415] ^ x[126];
  assign t[326] = t[416] ^ x[130];
  assign t[327] = t[417] ^ x[129];
  assign t[328] = t[418] ^ x[133];
  assign t[329] = t[419] ^ x[132];
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = t[420] ^ x[136];
  assign t[331] = t[421] ^ x[135];
  assign t[332] = t[422] ^ x[139];
  assign t[333] = t[423] ^ x[138];
  assign t[334] = t[424] ^ x[142];
  assign t[335] = t[425] ^ x[141];
  assign t[336] = t[426] ^ x[145];
  assign t[337] = t[427] ^ x[144];
  assign t[338] = t[428] ^ x[148];
  assign t[339] = t[429] ^ x[147];
  assign t[33] = t[52] ^ t[40];
  assign t[340] = t[430] ^ x[151];
  assign t[341] = t[431] ^ x[150];
  assign t[342] = (x[0]);
  assign t[343] = (x[0]);
  assign t[344] = (x[6]);
  assign t[345] = (x[6]);
  assign t[346] = (x[9]);
  assign t[347] = (x[9]);
  assign t[348] = (x[12]);
  assign t[349] = (x[12]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[15]);
  assign t[351] = (x[15]);
  assign t[352] = (x[20]);
  assign t[353] = (x[20]);
  assign t[354] = (x[25]);
  assign t[355] = (x[25]);
  assign t[356] = (x[30]);
  assign t[357] = (x[30]);
  assign t[358] = (x[33]);
  assign t[359] = (x[33]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[36]);
  assign t[361] = (x[36]);
  assign t[362] = (x[39]);
  assign t[363] = (x[39]);
  assign t[364] = (x[44]);
  assign t[365] = (x[44]);
  assign t[366] = (x[49]);
  assign t[367] = (x[49]);
  assign t[368] = (x[52]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[57] & t[58]);
  assign t[370] = (x[55]);
  assign t[371] = (x[55]);
  assign t[372] = (x[58]);
  assign t[373] = (x[58]);
  assign t[374] = (x[63]);
  assign t[375] = (x[63]);
  assign t[376] = (x[68]);
  assign t[377] = (x[68]);
  assign t[378] = (x[71]);
  assign t[379] = (x[71]);
  assign t[37] = ~(t[59] & t[123]);
  assign t[380] = (x[74]);
  assign t[381] = (x[74]);
  assign t[382] = (x[77]);
  assign t[383] = (x[77]);
  assign t[384] = (x[80]);
  assign t[385] = (x[80]);
  assign t[386] = (x[83]);
  assign t[387] = (x[83]);
  assign t[388] = (x[86]);
  assign t[389] = (x[86]);
  assign t[38] = t[120] ? x[29] : x[28];
  assign t[390] = (x[89]);
  assign t[391] = (x[89]);
  assign t[392] = (x[92]);
  assign t[393] = (x[92]);
  assign t[394] = (x[95]);
  assign t[395] = (x[95]);
  assign t[396] = (x[98]);
  assign t[397] = (x[98]);
  assign t[398] = (x[101]);
  assign t[399] = (x[101]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[104]);
  assign t[401] = (x[104]);
  assign t[402] = (x[107]);
  assign t[403] = (x[107]);
  assign t[404] = (x[110]);
  assign t[405] = (x[110]);
  assign t[406] = (x[113]);
  assign t[407] = (x[113]);
  assign t[408] = (x[116]);
  assign t[409] = (x[116]);
  assign t[40] = ~(t[62] & t[63]);
  assign t[410] = (x[119]);
  assign t[411] = (x[119]);
  assign t[412] = (x[122]);
  assign t[413] = (x[122]);
  assign t[414] = (x[125]);
  assign t[415] = (x[125]);
  assign t[416] = (x[128]);
  assign t[417] = (x[128]);
  assign t[418] = (x[131]);
  assign t[419] = (x[131]);
  assign t[41] = t[64] ^ t[65];
  assign t[420] = (x[134]);
  assign t[421] = (x[134]);
  assign t[422] = (x[137]);
  assign t[423] = (x[137]);
  assign t[424] = (x[140]);
  assign t[425] = (x[140]);
  assign t[426] = (x[143]);
  assign t[427] = (x[143]);
  assign t[428] = (x[146]);
  assign t[429] = (x[146]);
  assign t[42] = ~(t[66] & t[67]);
  assign t[430] = (x[149]);
  assign t[431] = (x[149]);
  assign t[43] = t[68] ^ t[42];
  assign t[44] = ~(t[124]);
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[23]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[126]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[127]);
  assign t[52] = t[16] ? x[43] : x[42];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = ~(t[79] & t[128]);
  assign t[55] = t[16] ? x[48] : x[47];
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = ~(t[129]);
  assign t[58] = ~(t[130]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[86] & t[131]);
  assign t[62] = ~(t[87] & t[88]);
  assign t[63] = ~(t[89] & t[132]);
  assign t[64] = t[120] ? x[62] : x[61];
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[93]);
  assign t[67] = ~(t[94] & t[133]);
  assign t[68] = t[120] ? x[67] : x[66];
  assign t[69] = ~(t[125] & t[124]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[134]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[95] & t[96]);
  assign t[74] = ~(t[137]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[97] & t[98]);
  assign t[77] = ~(t[139]);
  assign t[78] = ~(t[140]);
  assign t[79] = ~(t[99] & t[100]);
  assign t[7] = ~(t[118] & t[119]);
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[103] & t[141]);
  assign t[82] = ~(t[130] & t[129]);
  assign t[83] = ~(t[142]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[104] & t[105]);
  assign t[87] = ~(t[145]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[120] & t[121]);
  assign t[90] = ~(t[108] & t[109]);
  assign t[91] = ~(t[110] & t[147]);
  assign t[92] = ~(t[148]);
  assign t[93] = ~(t[149]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[136] & t[135]);
  assign t[96] = ~(t[150]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[151]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [151:0] x;
 output y;

 wire [431:0] t;
  assign t[0] = t[1] ? t[2] : t[117];
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[113] & t[114]);
  assign t[104] = ~(t[144] & t[143]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[156]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[115] & t[116]);
  assign t[111] = ~(t[149] & t[148]);
  assign t[112] = ~(t[159]);
  assign t[113] = ~(t[154] & t[153]);
  assign t[114] = ~(t[160]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[18] : x[19];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = t[207] ^ x[2];
  assign t[163] = t[208] ^ x[8];
  assign t[164] = t[209] ^ x[11];
  assign t[165] = t[210] ^ x[14];
  assign t[166] = t[211] ^ x[17];
  assign t[167] = t[212] ^ x[22];
  assign t[168] = t[213] ^ x[27];
  assign t[169] = t[214] ^ x[32];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[35];
  assign t[171] = t[216] ^ x[38];
  assign t[172] = t[217] ^ x[41];
  assign t[173] = t[218] ^ x[46];
  assign t[174] = t[219] ^ x[51];
  assign t[175] = t[220] ^ x[54];
  assign t[176] = t[221] ^ x[57];
  assign t[177] = t[222] ^ x[60];
  assign t[178] = t[223] ^ x[65];
  assign t[179] = t[224] ^ x[70];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[73];
  assign t[181] = t[226] ^ x[76];
  assign t[182] = t[227] ^ x[79];
  assign t[183] = t[228] ^ x[82];
  assign t[184] = t[229] ^ x[85];
  assign t[185] = t[230] ^ x[88];
  assign t[186] = t[231] ^ x[91];
  assign t[187] = t[232] ^ x[94];
  assign t[188] = t[233] ^ x[97];
  assign t[189] = t[234] ^ x[100];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[103];
  assign t[191] = t[236] ^ x[106];
  assign t[192] = t[237] ^ x[109];
  assign t[193] = t[238] ^ x[112];
  assign t[194] = t[239] ^ x[115];
  assign t[195] = t[240] ^ x[118];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[124];
  assign t[198] = t[243] ^ x[127];
  assign t[199] = t[244] ^ x[130];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[133];
  assign t[201] = t[246] ^ x[136];
  assign t[202] = t[247] ^ x[139];
  assign t[203] = t[248] ^ x[142];
  assign t[204] = t[249] ^ x[145];
  assign t[205] = t[250] ^ x[148];
  assign t[206] = t[251] ^ x[151];
  assign t[207] = (t[252] & ~t[253]);
  assign t[208] = (t[254] & ~t[255]);
  assign t[209] = (t[256] & ~t[257]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[258] & ~t[259]);
  assign t[211] = (t[260] & ~t[261]);
  assign t[212] = (t[262] & ~t[263]);
  assign t[213] = (t[264] & ~t[265]);
  assign t[214] = (t[266] & ~t[267]);
  assign t[215] = (t[268] & ~t[269]);
  assign t[216] = (t[270] & ~t[271]);
  assign t[217] = (t[272] & ~t[273]);
  assign t[218] = (t[274] & ~t[275]);
  assign t[219] = (t[276] & ~t[277]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[278] & ~t[279]);
  assign t[221] = (t[280] & ~t[281]);
  assign t[222] = (t[282] & ~t[283]);
  assign t[223] = (t[284] & ~t[285]);
  assign t[224] = (t[286] & ~t[287]);
  assign t[225] = (t[288] & ~t[289]);
  assign t[226] = (t[290] & ~t[291]);
  assign t[227] = (t[292] & ~t[293]);
  assign t[228] = (t[294] & ~t[295]);
  assign t[229] = (t[296] & ~t[297]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[298] & ~t[299]);
  assign t[231] = (t[300] & ~t[301]);
  assign t[232] = (t[302] & ~t[303]);
  assign t[233] = (t[304] & ~t[305]);
  assign t[234] = (t[306] & ~t[307]);
  assign t[235] = (t[308] & ~t[309]);
  assign t[236] = (t[310] & ~t[311]);
  assign t[237] = (t[312] & ~t[313]);
  assign t[238] = (t[314] & ~t[315]);
  assign t[239] = (t[316] & ~t[317]);
  assign t[23] = ~(t[120]);
  assign t[240] = (t[318] & ~t[319]);
  assign t[241] = (t[320] & ~t[321]);
  assign t[242] = (t[322] & ~t[323]);
  assign t[243] = (t[324] & ~t[325]);
  assign t[244] = (t[326] & ~t[327]);
  assign t[245] = (t[328] & ~t[329]);
  assign t[246] = (t[330] & ~t[331]);
  assign t[247] = (t[332] & ~t[333]);
  assign t[248] = (t[334] & ~t[335]);
  assign t[249] = (t[336] & ~t[337]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (t[338] & ~t[339]);
  assign t[251] = (t[340] & ~t[341]);
  assign t[252] = t[342] ^ x[2];
  assign t[253] = t[343] ^ x[1];
  assign t[254] = t[344] ^ x[8];
  assign t[255] = t[345] ^ x[7];
  assign t[256] = t[346] ^ x[11];
  assign t[257] = t[347] ^ x[10];
  assign t[258] = t[348] ^ x[14];
  assign t[259] = t[349] ^ x[13];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[17];
  assign t[261] = t[351] ^ x[16];
  assign t[262] = t[352] ^ x[22];
  assign t[263] = t[353] ^ x[21];
  assign t[264] = t[354] ^ x[27];
  assign t[265] = t[355] ^ x[26];
  assign t[266] = t[356] ^ x[32];
  assign t[267] = t[357] ^ x[31];
  assign t[268] = t[358] ^ x[35];
  assign t[269] = t[359] ^ x[34];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[38];
  assign t[271] = t[361] ^ x[37];
  assign t[272] = t[362] ^ x[41];
  assign t[273] = t[363] ^ x[40];
  assign t[274] = t[364] ^ x[46];
  assign t[275] = t[365] ^ x[45];
  assign t[276] = t[366] ^ x[51];
  assign t[277] = t[367] ^ x[50];
  assign t[278] = t[368] ^ x[54];
  assign t[279] = t[369] ^ x[53];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[57];
  assign t[281] = t[371] ^ x[56];
  assign t[282] = t[372] ^ x[60];
  assign t[283] = t[373] ^ x[59];
  assign t[284] = t[374] ^ x[65];
  assign t[285] = t[375] ^ x[64];
  assign t[286] = t[376] ^ x[70];
  assign t[287] = t[377] ^ x[69];
  assign t[288] = t[378] ^ x[73];
  assign t[289] = t[379] ^ x[72];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[76];
  assign t[291] = t[381] ^ x[75];
  assign t[292] = t[382] ^ x[79];
  assign t[293] = t[383] ^ x[78];
  assign t[294] = t[384] ^ x[82];
  assign t[295] = t[385] ^ x[81];
  assign t[296] = t[386] ^ x[85];
  assign t[297] = t[387] ^ x[84];
  assign t[298] = t[388] ^ x[88];
  assign t[299] = t[389] ^ x[87];
  assign t[29] = ~(t[46] & t[122]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[91];
  assign t[301] = t[391] ^ x[90];
  assign t[302] = t[392] ^ x[94];
  assign t[303] = t[393] ^ x[93];
  assign t[304] = t[394] ^ x[97];
  assign t[305] = t[395] ^ x[96];
  assign t[306] = t[396] ^ x[100];
  assign t[307] = t[397] ^ x[99];
  assign t[308] = t[398] ^ x[103];
  assign t[309] = t[399] ^ x[102];
  assign t[30] = t[47] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[106];
  assign t[311] = t[401] ^ x[105];
  assign t[312] = t[402] ^ x[109];
  assign t[313] = t[403] ^ x[108];
  assign t[314] = t[404] ^ x[112];
  assign t[315] = t[405] ^ x[111];
  assign t[316] = t[406] ^ x[115];
  assign t[317] = t[407] ^ x[114];
  assign t[318] = t[408] ^ x[118];
  assign t[319] = t[409] ^ x[117];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[410] ^ x[121];
  assign t[321] = t[411] ^ x[120];
  assign t[322] = t[412] ^ x[124];
  assign t[323] = t[413] ^ x[123];
  assign t[324] = t[414] ^ x[127];
  assign t[325] = t[415] ^ x[126];
  assign t[326] = t[416] ^ x[130];
  assign t[327] = t[417] ^ x[129];
  assign t[328] = t[418] ^ x[133];
  assign t[329] = t[419] ^ x[132];
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = t[420] ^ x[136];
  assign t[331] = t[421] ^ x[135];
  assign t[332] = t[422] ^ x[139];
  assign t[333] = t[423] ^ x[138];
  assign t[334] = t[424] ^ x[142];
  assign t[335] = t[425] ^ x[141];
  assign t[336] = t[426] ^ x[145];
  assign t[337] = t[427] ^ x[144];
  assign t[338] = t[428] ^ x[148];
  assign t[339] = t[429] ^ x[147];
  assign t[33] = t[52] ^ t[40];
  assign t[340] = t[430] ^ x[151];
  assign t[341] = t[431] ^ x[150];
  assign t[342] = (x[0]);
  assign t[343] = (x[0]);
  assign t[344] = (x[6]);
  assign t[345] = (x[6]);
  assign t[346] = (x[9]);
  assign t[347] = (x[9]);
  assign t[348] = (x[12]);
  assign t[349] = (x[12]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[15]);
  assign t[351] = (x[15]);
  assign t[352] = (x[20]);
  assign t[353] = (x[20]);
  assign t[354] = (x[25]);
  assign t[355] = (x[25]);
  assign t[356] = (x[30]);
  assign t[357] = (x[30]);
  assign t[358] = (x[33]);
  assign t[359] = (x[33]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[36]);
  assign t[361] = (x[36]);
  assign t[362] = (x[39]);
  assign t[363] = (x[39]);
  assign t[364] = (x[44]);
  assign t[365] = (x[44]);
  assign t[366] = (x[49]);
  assign t[367] = (x[49]);
  assign t[368] = (x[52]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[57] & t[58]);
  assign t[370] = (x[55]);
  assign t[371] = (x[55]);
  assign t[372] = (x[58]);
  assign t[373] = (x[58]);
  assign t[374] = (x[63]);
  assign t[375] = (x[63]);
  assign t[376] = (x[68]);
  assign t[377] = (x[68]);
  assign t[378] = (x[71]);
  assign t[379] = (x[71]);
  assign t[37] = ~(t[59] & t[123]);
  assign t[380] = (x[74]);
  assign t[381] = (x[74]);
  assign t[382] = (x[77]);
  assign t[383] = (x[77]);
  assign t[384] = (x[80]);
  assign t[385] = (x[80]);
  assign t[386] = (x[83]);
  assign t[387] = (x[83]);
  assign t[388] = (x[86]);
  assign t[389] = (x[86]);
  assign t[38] = t[120] ? x[29] : x[28];
  assign t[390] = (x[89]);
  assign t[391] = (x[89]);
  assign t[392] = (x[92]);
  assign t[393] = (x[92]);
  assign t[394] = (x[95]);
  assign t[395] = (x[95]);
  assign t[396] = (x[98]);
  assign t[397] = (x[98]);
  assign t[398] = (x[101]);
  assign t[399] = (x[101]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[104]);
  assign t[401] = (x[104]);
  assign t[402] = (x[107]);
  assign t[403] = (x[107]);
  assign t[404] = (x[110]);
  assign t[405] = (x[110]);
  assign t[406] = (x[113]);
  assign t[407] = (x[113]);
  assign t[408] = (x[116]);
  assign t[409] = (x[116]);
  assign t[40] = ~(t[62] & t[63]);
  assign t[410] = (x[119]);
  assign t[411] = (x[119]);
  assign t[412] = (x[122]);
  assign t[413] = (x[122]);
  assign t[414] = (x[125]);
  assign t[415] = (x[125]);
  assign t[416] = (x[128]);
  assign t[417] = (x[128]);
  assign t[418] = (x[131]);
  assign t[419] = (x[131]);
  assign t[41] = t[64] ^ t[65];
  assign t[420] = (x[134]);
  assign t[421] = (x[134]);
  assign t[422] = (x[137]);
  assign t[423] = (x[137]);
  assign t[424] = (x[140]);
  assign t[425] = (x[140]);
  assign t[426] = (x[143]);
  assign t[427] = (x[143]);
  assign t[428] = (x[146]);
  assign t[429] = (x[146]);
  assign t[42] = ~(t[66] & t[67]);
  assign t[430] = (x[149]);
  assign t[431] = (x[149]);
  assign t[43] = t[68] ^ t[42];
  assign t[44] = ~(t[124]);
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[23]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[126]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[127]);
  assign t[52] = t[16] ? x[43] : x[42];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = ~(t[79] & t[128]);
  assign t[55] = t[16] ? x[48] : x[47];
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = ~(t[129]);
  assign t[58] = ~(t[130]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[86] & t[131]);
  assign t[62] = ~(t[87] & t[88]);
  assign t[63] = ~(t[89] & t[132]);
  assign t[64] = t[120] ? x[62] : x[61];
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[93]);
  assign t[67] = ~(t[94] & t[133]);
  assign t[68] = t[120] ? x[67] : x[66];
  assign t[69] = ~(t[125] & t[124]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[134]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[95] & t[96]);
  assign t[74] = ~(t[137]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[97] & t[98]);
  assign t[77] = ~(t[139]);
  assign t[78] = ~(t[140]);
  assign t[79] = ~(t[99] & t[100]);
  assign t[7] = ~(t[118] & t[119]);
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[103] & t[141]);
  assign t[82] = ~(t[130] & t[129]);
  assign t[83] = ~(t[142]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[104] & t[105]);
  assign t[87] = ~(t[145]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[120] & t[121]);
  assign t[90] = ~(t[108] & t[109]);
  assign t[91] = ~(t[110] & t[147]);
  assign t[92] = ~(t[148]);
  assign t[93] = ~(t[149]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[136] & t[135]);
  assign t[96] = ~(t[150]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[151]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [151:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[107];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[106] | t[101]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[150]);
  assign t[106] = ~(t[151]);
  assign t[107] = (t[152]);
  assign t[108] = (t[153]);
  assign t[109] = (t[154]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = t[197] ^ x[2];
  assign t[153] = t[198] ^ x[8];
  assign t[154] = t[199] ^ x[11];
  assign t[155] = t[200] ^ x[14];
  assign t[156] = t[201] ^ x[17];
  assign t[157] = t[202] ^ x[22];
  assign t[158] = t[203] ^ x[27];
  assign t[159] = t[204] ^ x[32];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[205] ^ x[35];
  assign t[161] = t[206] ^ x[38];
  assign t[162] = t[207] ^ x[41];
  assign t[163] = t[208] ^ x[46];
  assign t[164] = t[209] ^ x[51];
  assign t[165] = t[210] ^ x[54];
  assign t[166] = t[211] ^ x[57];
  assign t[167] = t[212] ^ x[60];
  assign t[168] = t[213] ^ x[65];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[73];
  assign t[171] = t[216] ^ x[76];
  assign t[172] = t[217] ^ x[79];
  assign t[173] = t[218] ^ x[82];
  assign t[174] = t[219] ^ x[85];
  assign t[175] = t[220] ^ x[88];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[94];
  assign t[178] = t[223] ^ x[97];
  assign t[179] = t[224] ^ x[100];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[103];
  assign t[181] = t[226] ^ x[106];
  assign t[182] = t[227] ^ x[109];
  assign t[183] = t[228] ^ x[112];
  assign t[184] = t[229] ^ x[115];
  assign t[185] = t[230] ^ x[118];
  assign t[186] = t[231] ^ x[121];
  assign t[187] = t[232] ^ x[124];
  assign t[188] = t[233] ^ x[127];
  assign t[189] = t[234] ^ x[130];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[133];
  assign t[191] = t[236] ^ x[136];
  assign t[192] = t[237] ^ x[139];
  assign t[193] = t[238] ^ x[142];
  assign t[194] = t[239] ^ x[145];
  assign t[195] = t[240] ^ x[148];
  assign t[196] = t[241] ^ x[151];
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = (t[316] & ~t[317]);
  assign t[235] = (t[318] & ~t[319]);
  assign t[236] = (t[320] & ~t[321]);
  assign t[237] = (t[322] & ~t[323]);
  assign t[238] = (t[324] & ~t[325]);
  assign t[239] = (t[326] & ~t[327]);
  assign t[23] = ~(t[110]);
  assign t[240] = (t[328] & ~t[329]);
  assign t[241] = (t[330] & ~t[331]);
  assign t[242] = t[332] ^ x[2];
  assign t[243] = t[333] ^ x[1];
  assign t[244] = t[334] ^ x[8];
  assign t[245] = t[335] ^ x[7];
  assign t[246] = t[336] ^ x[11];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[14];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[340] ^ x[17];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[22];
  assign t[253] = t[343] ^ x[21];
  assign t[254] = t[344] ^ x[27];
  assign t[255] = t[345] ^ x[26];
  assign t[256] = t[346] ^ x[32];
  assign t[257] = t[347] ^ x[31];
  assign t[258] = t[348] ^ x[35];
  assign t[259] = t[349] ^ x[34];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[38];
  assign t[261] = t[351] ^ x[37];
  assign t[262] = t[352] ^ x[41];
  assign t[263] = t[353] ^ x[40];
  assign t[264] = t[354] ^ x[46];
  assign t[265] = t[355] ^ x[45];
  assign t[266] = t[356] ^ x[51];
  assign t[267] = t[357] ^ x[50];
  assign t[268] = t[358] ^ x[54];
  assign t[269] = t[359] ^ x[53];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[57];
  assign t[271] = t[361] ^ x[56];
  assign t[272] = t[362] ^ x[60];
  assign t[273] = t[363] ^ x[59];
  assign t[274] = t[364] ^ x[65];
  assign t[275] = t[365] ^ x[64];
  assign t[276] = t[366] ^ x[70];
  assign t[277] = t[367] ^ x[69];
  assign t[278] = t[368] ^ x[73];
  assign t[279] = t[369] ^ x[72];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[76];
  assign t[281] = t[371] ^ x[75];
  assign t[282] = t[372] ^ x[79];
  assign t[283] = t[373] ^ x[78];
  assign t[284] = t[374] ^ x[82];
  assign t[285] = t[375] ^ x[81];
  assign t[286] = t[376] ^ x[85];
  assign t[287] = t[377] ^ x[84];
  assign t[288] = t[378] ^ x[88];
  assign t[289] = t[379] ^ x[87];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[91];
  assign t[291] = t[381] ^ x[90];
  assign t[292] = t[382] ^ x[94];
  assign t[293] = t[383] ^ x[93];
  assign t[294] = t[384] ^ x[97];
  assign t[295] = t[385] ^ x[96];
  assign t[296] = t[386] ^ x[100];
  assign t[297] = t[387] ^ x[99];
  assign t[298] = t[388] ^ x[103];
  assign t[299] = t[389] ^ x[102];
  assign t[29] = t[46] | t[112];
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[106];
  assign t[301] = t[391] ^ x[105];
  assign t[302] = t[392] ^ x[109];
  assign t[303] = t[393] ^ x[108];
  assign t[304] = t[394] ^ x[112];
  assign t[305] = t[395] ^ x[111];
  assign t[306] = t[396] ^ x[115];
  assign t[307] = t[397] ^ x[114];
  assign t[308] = t[398] ^ x[118];
  assign t[309] = t[399] ^ x[117];
  assign t[30] = t[16] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[121];
  assign t[311] = t[401] ^ x[120];
  assign t[312] = t[402] ^ x[124];
  assign t[313] = t[403] ^ x[123];
  assign t[314] = t[404] ^ x[127];
  assign t[315] = t[405] ^ x[126];
  assign t[316] = t[406] ^ x[130];
  assign t[317] = t[407] ^ x[129];
  assign t[318] = t[408] ^ x[133];
  assign t[319] = t[409] ^ x[132];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[410] ^ x[136];
  assign t[321] = t[411] ^ x[135];
  assign t[322] = t[412] ^ x[139];
  assign t[323] = t[413] ^ x[138];
  assign t[324] = t[414] ^ x[142];
  assign t[325] = t[415] ^ x[141];
  assign t[326] = t[416] ^ x[145];
  assign t[327] = t[417] ^ x[144];
  assign t[328] = t[418] ^ x[148];
  assign t[329] = t[419] ^ x[147];
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = t[420] ^ x[151];
  assign t[331] = t[421] ^ x[150];
  assign t[332] = (x[0]);
  assign t[333] = (x[0]);
  assign t[334] = (x[6]);
  assign t[335] = (x[6]);
  assign t[336] = (x[9]);
  assign t[337] = (x[9]);
  assign t[338] = (x[12]);
  assign t[339] = (x[12]);
  assign t[33] = t[51] ^ t[40];
  assign t[340] = (x[15]);
  assign t[341] = (x[15]);
  assign t[342] = (x[20]);
  assign t[343] = (x[20]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[30]);
  assign t[347] = (x[30]);
  assign t[348] = (x[33]);
  assign t[349] = (x[33]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[36]);
  assign t[351] = (x[36]);
  assign t[352] = (x[39]);
  assign t[353] = (x[39]);
  assign t[354] = (x[44]);
  assign t[355] = (x[44]);
  assign t[356] = (x[49]);
  assign t[357] = (x[49]);
  assign t[358] = (x[52]);
  assign t[359] = (x[52]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[55]);
  assign t[361] = (x[55]);
  assign t[362] = (x[58]);
  assign t[363] = (x[58]);
  assign t[364] = (x[63]);
  assign t[365] = (x[63]);
  assign t[366] = (x[68]);
  assign t[367] = (x[68]);
  assign t[368] = (x[71]);
  assign t[369] = (x[71]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[74]);
  assign t[371] = (x[74]);
  assign t[372] = (x[77]);
  assign t[373] = (x[77]);
  assign t[374] = (x[80]);
  assign t[375] = (x[80]);
  assign t[376] = (x[83]);
  assign t[377] = (x[83]);
  assign t[378] = (x[86]);
  assign t[379] = (x[86]);
  assign t[37] = t[58] | t[113];
  assign t[380] = (x[89]);
  assign t[381] = (x[89]);
  assign t[382] = (x[92]);
  assign t[383] = (x[92]);
  assign t[384] = (x[95]);
  assign t[385] = (x[95]);
  assign t[386] = (x[98]);
  assign t[387] = (x[98]);
  assign t[388] = (x[101]);
  assign t[389] = (x[101]);
  assign t[38] = t[110] ? x[29] : x[28];
  assign t[390] = (x[104]);
  assign t[391] = (x[104]);
  assign t[392] = (x[107]);
  assign t[393] = (x[107]);
  assign t[394] = (x[110]);
  assign t[395] = (x[110]);
  assign t[396] = (x[113]);
  assign t[397] = (x[113]);
  assign t[398] = (x[116]);
  assign t[399] = (x[116]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[119]);
  assign t[401] = (x[119]);
  assign t[402] = (x[122]);
  assign t[403] = (x[122]);
  assign t[404] = (x[125]);
  assign t[405] = (x[125]);
  assign t[406] = (x[128]);
  assign t[407] = (x[128]);
  assign t[408] = (x[131]);
  assign t[409] = (x[131]);
  assign t[40] = ~(t[61] & t[62]);
  assign t[410] = (x[134]);
  assign t[411] = (x[134]);
  assign t[412] = (x[137]);
  assign t[413] = (x[137]);
  assign t[414] = (x[140]);
  assign t[415] = (x[140]);
  assign t[416] = (x[143]);
  assign t[417] = (x[143]);
  assign t[418] = (x[146]);
  assign t[419] = (x[146]);
  assign t[41] = t[63] ^ t[64];
  assign t[420] = (x[149]);
  assign t[421] = (x[149]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[114]);
  assign t[45] = ~(t[115]);
  assign t[46] = ~(t[68] | t[44]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[116];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[74] | t[117];
  assign t[51] = t[75] ? x[43] : x[42];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[118];
  assign t[54] = t[75] ? x[48] : x[47];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[119]);
  assign t[57] = ~(t[120]);
  assign t[58] = ~(t[81] | t[56]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[84] | t[121];
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = t[87] | t[122];
  assign t[63] = t[110] ? x[62] : x[61];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = t[92] | t[123];
  assign t[67] = t[110] ? x[67] : x[66];
  assign t[68] = ~(t[124]);
  assign t[69] = ~(t[125]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[93] | t[69]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[94] | t[72]);
  assign t[75] = ~(t[23]);
  assign t[76] = ~(t[129]);
  assign t[77] = ~(t[130]);
  assign t[78] = ~(t[95] | t[76]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = ~(t[108] & t[109]);
  assign t[80] = t[98] | t[131];
  assign t[81] = ~(t[132]);
  assign t[82] = ~(t[133]);
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[135]);
  assign t[86] = ~(t[136]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[137];
  assign t[8] = ~(t[110] & t[111]);
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[141]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[105] | t[96]);
  assign t[99] = ~(t[145]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [151:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[107];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[106] | t[101]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[150]);
  assign t[106] = ~(t[151]);
  assign t[107] = (t[152]);
  assign t[108] = (t[153]);
  assign t[109] = (t[154]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = t[197] ^ x[2];
  assign t[153] = t[198] ^ x[8];
  assign t[154] = t[199] ^ x[11];
  assign t[155] = t[200] ^ x[14];
  assign t[156] = t[201] ^ x[17];
  assign t[157] = t[202] ^ x[22];
  assign t[158] = t[203] ^ x[27];
  assign t[159] = t[204] ^ x[32];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[205] ^ x[35];
  assign t[161] = t[206] ^ x[38];
  assign t[162] = t[207] ^ x[41];
  assign t[163] = t[208] ^ x[46];
  assign t[164] = t[209] ^ x[51];
  assign t[165] = t[210] ^ x[54];
  assign t[166] = t[211] ^ x[57];
  assign t[167] = t[212] ^ x[60];
  assign t[168] = t[213] ^ x[65];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[73];
  assign t[171] = t[216] ^ x[76];
  assign t[172] = t[217] ^ x[79];
  assign t[173] = t[218] ^ x[82];
  assign t[174] = t[219] ^ x[85];
  assign t[175] = t[220] ^ x[88];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[94];
  assign t[178] = t[223] ^ x[97];
  assign t[179] = t[224] ^ x[100];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[103];
  assign t[181] = t[226] ^ x[106];
  assign t[182] = t[227] ^ x[109];
  assign t[183] = t[228] ^ x[112];
  assign t[184] = t[229] ^ x[115];
  assign t[185] = t[230] ^ x[118];
  assign t[186] = t[231] ^ x[121];
  assign t[187] = t[232] ^ x[124];
  assign t[188] = t[233] ^ x[127];
  assign t[189] = t[234] ^ x[130];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[133];
  assign t[191] = t[236] ^ x[136];
  assign t[192] = t[237] ^ x[139];
  assign t[193] = t[238] ^ x[142];
  assign t[194] = t[239] ^ x[145];
  assign t[195] = t[240] ^ x[148];
  assign t[196] = t[241] ^ x[151];
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = (t[316] & ~t[317]);
  assign t[235] = (t[318] & ~t[319]);
  assign t[236] = (t[320] & ~t[321]);
  assign t[237] = (t[322] & ~t[323]);
  assign t[238] = (t[324] & ~t[325]);
  assign t[239] = (t[326] & ~t[327]);
  assign t[23] = ~(t[110]);
  assign t[240] = (t[328] & ~t[329]);
  assign t[241] = (t[330] & ~t[331]);
  assign t[242] = t[332] ^ x[2];
  assign t[243] = t[333] ^ x[1];
  assign t[244] = t[334] ^ x[8];
  assign t[245] = t[335] ^ x[7];
  assign t[246] = t[336] ^ x[11];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[14];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[340] ^ x[17];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[22];
  assign t[253] = t[343] ^ x[21];
  assign t[254] = t[344] ^ x[27];
  assign t[255] = t[345] ^ x[26];
  assign t[256] = t[346] ^ x[32];
  assign t[257] = t[347] ^ x[31];
  assign t[258] = t[348] ^ x[35];
  assign t[259] = t[349] ^ x[34];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[38];
  assign t[261] = t[351] ^ x[37];
  assign t[262] = t[352] ^ x[41];
  assign t[263] = t[353] ^ x[40];
  assign t[264] = t[354] ^ x[46];
  assign t[265] = t[355] ^ x[45];
  assign t[266] = t[356] ^ x[51];
  assign t[267] = t[357] ^ x[50];
  assign t[268] = t[358] ^ x[54];
  assign t[269] = t[359] ^ x[53];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[57];
  assign t[271] = t[361] ^ x[56];
  assign t[272] = t[362] ^ x[60];
  assign t[273] = t[363] ^ x[59];
  assign t[274] = t[364] ^ x[65];
  assign t[275] = t[365] ^ x[64];
  assign t[276] = t[366] ^ x[70];
  assign t[277] = t[367] ^ x[69];
  assign t[278] = t[368] ^ x[73];
  assign t[279] = t[369] ^ x[72];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[76];
  assign t[281] = t[371] ^ x[75];
  assign t[282] = t[372] ^ x[79];
  assign t[283] = t[373] ^ x[78];
  assign t[284] = t[374] ^ x[82];
  assign t[285] = t[375] ^ x[81];
  assign t[286] = t[376] ^ x[85];
  assign t[287] = t[377] ^ x[84];
  assign t[288] = t[378] ^ x[88];
  assign t[289] = t[379] ^ x[87];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[91];
  assign t[291] = t[381] ^ x[90];
  assign t[292] = t[382] ^ x[94];
  assign t[293] = t[383] ^ x[93];
  assign t[294] = t[384] ^ x[97];
  assign t[295] = t[385] ^ x[96];
  assign t[296] = t[386] ^ x[100];
  assign t[297] = t[387] ^ x[99];
  assign t[298] = t[388] ^ x[103];
  assign t[299] = t[389] ^ x[102];
  assign t[29] = t[46] | t[112];
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[106];
  assign t[301] = t[391] ^ x[105];
  assign t[302] = t[392] ^ x[109];
  assign t[303] = t[393] ^ x[108];
  assign t[304] = t[394] ^ x[112];
  assign t[305] = t[395] ^ x[111];
  assign t[306] = t[396] ^ x[115];
  assign t[307] = t[397] ^ x[114];
  assign t[308] = t[398] ^ x[118];
  assign t[309] = t[399] ^ x[117];
  assign t[30] = t[16] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[121];
  assign t[311] = t[401] ^ x[120];
  assign t[312] = t[402] ^ x[124];
  assign t[313] = t[403] ^ x[123];
  assign t[314] = t[404] ^ x[127];
  assign t[315] = t[405] ^ x[126];
  assign t[316] = t[406] ^ x[130];
  assign t[317] = t[407] ^ x[129];
  assign t[318] = t[408] ^ x[133];
  assign t[319] = t[409] ^ x[132];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[410] ^ x[136];
  assign t[321] = t[411] ^ x[135];
  assign t[322] = t[412] ^ x[139];
  assign t[323] = t[413] ^ x[138];
  assign t[324] = t[414] ^ x[142];
  assign t[325] = t[415] ^ x[141];
  assign t[326] = t[416] ^ x[145];
  assign t[327] = t[417] ^ x[144];
  assign t[328] = t[418] ^ x[148];
  assign t[329] = t[419] ^ x[147];
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = t[420] ^ x[151];
  assign t[331] = t[421] ^ x[150];
  assign t[332] = (x[0]);
  assign t[333] = (x[0]);
  assign t[334] = (x[6]);
  assign t[335] = (x[6]);
  assign t[336] = (x[9]);
  assign t[337] = (x[9]);
  assign t[338] = (x[12]);
  assign t[339] = (x[12]);
  assign t[33] = t[51] ^ t[40];
  assign t[340] = (x[15]);
  assign t[341] = (x[15]);
  assign t[342] = (x[20]);
  assign t[343] = (x[20]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[30]);
  assign t[347] = (x[30]);
  assign t[348] = (x[33]);
  assign t[349] = (x[33]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[36]);
  assign t[351] = (x[36]);
  assign t[352] = (x[39]);
  assign t[353] = (x[39]);
  assign t[354] = (x[44]);
  assign t[355] = (x[44]);
  assign t[356] = (x[49]);
  assign t[357] = (x[49]);
  assign t[358] = (x[52]);
  assign t[359] = (x[52]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[55]);
  assign t[361] = (x[55]);
  assign t[362] = (x[58]);
  assign t[363] = (x[58]);
  assign t[364] = (x[63]);
  assign t[365] = (x[63]);
  assign t[366] = (x[68]);
  assign t[367] = (x[68]);
  assign t[368] = (x[71]);
  assign t[369] = (x[71]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[74]);
  assign t[371] = (x[74]);
  assign t[372] = (x[77]);
  assign t[373] = (x[77]);
  assign t[374] = (x[80]);
  assign t[375] = (x[80]);
  assign t[376] = (x[83]);
  assign t[377] = (x[83]);
  assign t[378] = (x[86]);
  assign t[379] = (x[86]);
  assign t[37] = t[58] | t[113];
  assign t[380] = (x[89]);
  assign t[381] = (x[89]);
  assign t[382] = (x[92]);
  assign t[383] = (x[92]);
  assign t[384] = (x[95]);
  assign t[385] = (x[95]);
  assign t[386] = (x[98]);
  assign t[387] = (x[98]);
  assign t[388] = (x[101]);
  assign t[389] = (x[101]);
  assign t[38] = t[110] ? x[29] : x[28];
  assign t[390] = (x[104]);
  assign t[391] = (x[104]);
  assign t[392] = (x[107]);
  assign t[393] = (x[107]);
  assign t[394] = (x[110]);
  assign t[395] = (x[110]);
  assign t[396] = (x[113]);
  assign t[397] = (x[113]);
  assign t[398] = (x[116]);
  assign t[399] = (x[116]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[119]);
  assign t[401] = (x[119]);
  assign t[402] = (x[122]);
  assign t[403] = (x[122]);
  assign t[404] = (x[125]);
  assign t[405] = (x[125]);
  assign t[406] = (x[128]);
  assign t[407] = (x[128]);
  assign t[408] = (x[131]);
  assign t[409] = (x[131]);
  assign t[40] = ~(t[61] & t[62]);
  assign t[410] = (x[134]);
  assign t[411] = (x[134]);
  assign t[412] = (x[137]);
  assign t[413] = (x[137]);
  assign t[414] = (x[140]);
  assign t[415] = (x[140]);
  assign t[416] = (x[143]);
  assign t[417] = (x[143]);
  assign t[418] = (x[146]);
  assign t[419] = (x[146]);
  assign t[41] = t[63] ^ t[64];
  assign t[420] = (x[149]);
  assign t[421] = (x[149]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[114]);
  assign t[45] = ~(t[115]);
  assign t[46] = ~(t[68] | t[44]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[116];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[74] | t[117];
  assign t[51] = t[75] ? x[43] : x[42];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[118];
  assign t[54] = t[75] ? x[48] : x[47];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[119]);
  assign t[57] = ~(t[120]);
  assign t[58] = ~(t[81] | t[56]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[84] | t[121];
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = t[87] | t[122];
  assign t[63] = t[110] ? x[62] : x[61];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = t[92] | t[123];
  assign t[67] = t[110] ? x[67] : x[66];
  assign t[68] = ~(t[124]);
  assign t[69] = ~(t[125]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[93] | t[69]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[94] | t[72]);
  assign t[75] = ~(t[23]);
  assign t[76] = ~(t[129]);
  assign t[77] = ~(t[130]);
  assign t[78] = ~(t[95] | t[76]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = ~(t[108] & t[109]);
  assign t[80] = t[98] | t[131];
  assign t[81] = ~(t[132]);
  assign t[82] = ~(t[133]);
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[135]);
  assign t[86] = ~(t[136]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[137];
  assign t[8] = ~(t[110] & t[111]);
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[141]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[105] | t[96]);
  assign t[99] = ~(t[145]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind156(x, y);
 input [97:0] x;
 output y;

 wire [339:0] t;
  assign t[0] = t[1] ? t[2] : t[137];
  assign t[100] = ~(t[161]);
  assign t[101] = ~(t[154] | t[155]);
  assign t[102] = ~(t[162]);
  assign t[103] = ~(t[163]);
  assign t[104] = ~(t[119] | t[120]);
  assign t[105] = ~(t[121] | t[57]);
  assign t[106] = ~(x[4] | t[122]);
  assign t[107] = ~(t[123] & t[141]);
  assign t[108] = ~(t[124] & t[83]);
  assign t[109] = ~(t[123] & t[83]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = ~(t[124] & t[141]);
  assign t[111] = ~(x[4] & t[125]);
  assign t[112] = ~(t[117]);
  assign t[113] = t[80] | t[126];
  assign t[114] = ~(t[164]);
  assign t[115] = ~(t[159] | t[160]);
  assign t[116] = ~(t[127] & t[128]);
  assign t[117] = ~(t[80] | t[129]);
  assign t[118] = t[55] | t[130];
  assign t[119] = ~(t[165]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = ~(t[162] | t[163]);
  assign t[121] = ~(t[84] | t[131]);
  assign t[122] = ~(t[139]);
  assign t[123] = x[4] & t[139];
  assign t[124] = ~(x[4] | t[139]);
  assign t[125] = ~(t[139] | t[141]);
  assign t[126] = t[138] ? t[111] : t[132];
  assign t[127] = ~(t[133] | t[56]);
  assign t[128] = ~(t[134] & t[135]);
  assign t[129] = t[138] ? t[132] : t[111];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = ~(t[31]);
  assign t[131] = t[138] ? t[82] : t[132];
  assign t[132] = ~(t[106] & t[83]);
  assign t[133] = ~(t[84] | t[136]);
  assign t[134] = t[141] & t[50];
  assign t[135] = t[124] | t[123];
  assign t[136] = t[138] ? t[107] : t[108];
  assign t[137] = (t[166]);
  assign t[138] = (t[167]);
  assign t[139] = (t[168]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (t[169]);
  assign t[141] = (t[170]);
  assign t[142] = (t[171]);
  assign t[143] = (t[172]);
  assign t[144] = (t[173]);
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = t[140] ? x[19] : x[18];
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = t[195] ^ x[2];
  assign t[167] = t[196] ^ x[8];
  assign t[168] = t[197] ^ x[11];
  assign t[169] = t[198] ^ x[14];
  assign t[16] = t[21] | t[22];
  assign t[170] = t[199] ^ x[17];
  assign t[171] = t[200] ^ x[22];
  assign t[172] = t[201] ^ x[25];
  assign t[173] = t[202] ^ x[28];
  assign t[174] = t[203] ^ x[31];
  assign t[175] = t[204] ^ x[36];
  assign t[176] = t[205] ^ x[39];
  assign t[177] = t[206] ^ x[42];
  assign t[178] = t[207] ^ x[45];
  assign t[179] = t[208] ^ x[48];
  assign t[17] = ~(t[23] | t[24]);
  assign t[180] = t[209] ^ x[51];
  assign t[181] = t[210] ^ x[54];
  assign t[182] = t[211] ^ x[57];
  assign t[183] = t[212] ^ x[62];
  assign t[184] = t[213] ^ x[65];
  assign t[185] = t[214] ^ x[68];
  assign t[186] = t[215] ^ x[73];
  assign t[187] = t[216] ^ x[76];
  assign t[188] = t[217] ^ x[79];
  assign t[189] = t[218] ^ x[82];
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = t[219] ^ x[85];
  assign t[191] = t[220] ^ x[88];
  assign t[192] = t[221] ^ x[91];
  assign t[193] = t[222] ^ x[94];
  assign t[194] = t[223] ^ x[97];
  assign t[195] = (t[224] & ~t[225]);
  assign t[196] = (t[226] & ~t[227]);
  assign t[197] = (t[228] & ~t[229]);
  assign t[198] = (t[230] & ~t[231]);
  assign t[199] = (t[232] & ~t[233]);
  assign t[19] = x[4] ? t[28] : t[27];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[234] & ~t[235]);
  assign t[201] = (t[236] & ~t[237]);
  assign t[202] = (t[238] & ~t[239]);
  assign t[203] = (t[240] & ~t[241]);
  assign t[204] = (t[242] & ~t[243]);
  assign t[205] = (t[244] & ~t[245]);
  assign t[206] = (t[246] & ~t[247]);
  assign t[207] = (t[248] & ~t[249]);
  assign t[208] = (t[250] & ~t[251]);
  assign t[209] = (t[252] & ~t[253]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = (t[254] & ~t[255]);
  assign t[211] = (t[256] & ~t[257]);
  assign t[212] = (t[258] & ~t[259]);
  assign t[213] = (t[260] & ~t[261]);
  assign t[214] = (t[262] & ~t[263]);
  assign t[215] = (t[264] & ~t[265]);
  assign t[216] = (t[266] & ~t[267]);
  assign t[217] = (t[268] & ~t[269]);
  assign t[218] = (t[270] & ~t[271]);
  assign t[219] = (t[272] & ~t[273]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[274] & ~t[275]);
  assign t[221] = (t[276] & ~t[277]);
  assign t[222] = (t[278] & ~t[279]);
  assign t[223] = (t[280] & ~t[281]);
  assign t[224] = t[282] ^ x[2];
  assign t[225] = t[283] ^ x[1];
  assign t[226] = t[284] ^ x[8];
  assign t[227] = t[285] ^ x[7];
  assign t[228] = t[286] ^ x[11];
  assign t[229] = t[287] ^ x[10];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[288] ^ x[14];
  assign t[231] = t[289] ^ x[13];
  assign t[232] = t[290] ^ x[17];
  assign t[233] = t[291] ^ x[16];
  assign t[234] = t[292] ^ x[22];
  assign t[235] = t[293] ^ x[21];
  assign t[236] = t[294] ^ x[25];
  assign t[237] = t[295] ^ x[24];
  assign t[238] = t[296] ^ x[28];
  assign t[239] = t[297] ^ x[27];
  assign t[23] = ~(t[35] | t[36]);
  assign t[240] = t[298] ^ x[31];
  assign t[241] = t[299] ^ x[30];
  assign t[242] = t[300] ^ x[36];
  assign t[243] = t[301] ^ x[35];
  assign t[244] = t[302] ^ x[39];
  assign t[245] = t[303] ^ x[38];
  assign t[246] = t[304] ^ x[42];
  assign t[247] = t[305] ^ x[41];
  assign t[248] = t[306] ^ x[45];
  assign t[249] = t[307] ^ x[44];
  assign t[24] = ~(t[142] | t[37]);
  assign t[250] = t[308] ^ x[48];
  assign t[251] = t[309] ^ x[47];
  assign t[252] = t[310] ^ x[51];
  assign t[253] = t[311] ^ x[50];
  assign t[254] = t[312] ^ x[54];
  assign t[255] = t[313] ^ x[53];
  assign t[256] = t[314] ^ x[57];
  assign t[257] = t[315] ^ x[56];
  assign t[258] = t[316] ^ x[62];
  assign t[259] = t[317] ^ x[61];
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = t[318] ^ x[65];
  assign t[261] = t[319] ^ x[64];
  assign t[262] = t[320] ^ x[68];
  assign t[263] = t[321] ^ x[67];
  assign t[264] = t[322] ^ x[73];
  assign t[265] = t[323] ^ x[72];
  assign t[266] = t[324] ^ x[76];
  assign t[267] = t[325] ^ x[75];
  assign t[268] = t[326] ^ x[79];
  assign t[269] = t[327] ^ x[78];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[328] ^ x[82];
  assign t[271] = t[329] ^ x[81];
  assign t[272] = t[330] ^ x[85];
  assign t[273] = t[331] ^ x[84];
  assign t[274] = t[332] ^ x[88];
  assign t[275] = t[333] ^ x[87];
  assign t[276] = t[334] ^ x[91];
  assign t[277] = t[335] ^ x[90];
  assign t[278] = t[336] ^ x[94];
  assign t[279] = t[337] ^ x[93];
  assign t[27] = ~(t[42] | t[43]);
  assign t[280] = t[338] ^ x[97];
  assign t[281] = t[339] ^ x[96];
  assign t[282] = (x[0]);
  assign t[283] = (x[0]);
  assign t[284] = (x[6]);
  assign t[285] = (x[6]);
  assign t[286] = (x[9]);
  assign t[287] = (x[9]);
  assign t[288] = (x[12]);
  assign t[289] = (x[12]);
  assign t[28] = ~(t[44] ^ t[45]);
  assign t[290] = (x[15]);
  assign t[291] = (x[15]);
  assign t[292] = (x[20]);
  assign t[293] = (x[20]);
  assign t[294] = (x[23]);
  assign t[295] = (x[23]);
  assign t[296] = (x[26]);
  assign t[297] = (x[26]);
  assign t[298] = (x[29]);
  assign t[299] = (x[29]);
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[34]);
  assign t[301] = (x[34]);
  assign t[302] = (x[37]);
  assign t[303] = (x[37]);
  assign t[304] = (x[40]);
  assign t[305] = (x[40]);
  assign t[306] = (x[43]);
  assign t[307] = (x[43]);
  assign t[308] = (x[46]);
  assign t[309] = (x[46]);
  assign t[30] = ~(t[48] ^ t[49]);
  assign t[310] = (x[49]);
  assign t[311] = (x[49]);
  assign t[312] = (x[52]);
  assign t[313] = (x[52]);
  assign t[314] = (x[55]);
  assign t[315] = (x[55]);
  assign t[316] = (x[60]);
  assign t[317] = (x[60]);
  assign t[318] = (x[63]);
  assign t[319] = (x[63]);
  assign t[31] = ~(t[50] & t[51]);
  assign t[320] = (x[66]);
  assign t[321] = (x[66]);
  assign t[322] = (x[71]);
  assign t[323] = (x[71]);
  assign t[324] = (x[74]);
  assign t[325] = (x[74]);
  assign t[326] = (x[77]);
  assign t[327] = (x[77]);
  assign t[328] = (x[80]);
  assign t[329] = (x[80]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (x[83]);
  assign t[331] = (x[83]);
  assign t[332] = (x[86]);
  assign t[333] = (x[86]);
  assign t[334] = (x[89]);
  assign t[335] = (x[89]);
  assign t[336] = (x[92]);
  assign t[337] = (x[92]);
  assign t[338] = (x[95]);
  assign t[339] = (x[95]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[143]);
  assign t[36] = ~(t[144]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] | t[61]);
  assign t[39] = ~(t[145] | t[62]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[63] ? x[33] : x[32];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = ~(t[66] | t[67]);
  assign t[43] = ~(t[146] | t[68]);
  assign t[44] = ~(t[69] | t[70]);
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = ~(t[73] | t[74]);
  assign t[47] = ~(t[147] | t[75]);
  assign t[48] = ~(t[76] | t[77]);
  assign t[49] = ~(t[78] ^ t[79]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[80] | t[138]);
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = ~(t[139] | t[83]);
  assign t[53] = t[84] & t[138];
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[84] | t[86]);
  assign t[56] = ~(t[84] | t[87]);
  assign t[57] = ~(t[84] | t[88]);
  assign t[58] = ~(t[148]);
  assign t[59] = ~(t[143] | t[144]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[149]);
  assign t[61] = ~(t[150]);
  assign t[62] = ~(t[89] | t[90]);
  assign t[63] = ~(t[91]);
  assign t[64] = ~(t[21] | t[92]);
  assign t[65] = ~(t[54]);
  assign t[66] = ~(t[151]);
  assign t[67] = ~(t[152]);
  assign t[68] = ~(t[93] | t[94]);
  assign t[69] = ~(t[95] | t[96]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[153] | t[97]);
  assign t[71] = t[140] ? x[59] : x[58];
  assign t[72] = ~(t[98] & t[99]);
  assign t[73] = ~(t[154]);
  assign t[74] = ~(t[155]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[102] | t[103]);
  assign t[77] = ~(t[156] | t[104]);
  assign t[78] = t[140] ? x[70] : x[69];
  assign t[79] = ~(t[98] & t[105]);
  assign t[7] = ~(t[138] & t[139]);
  assign t[80] = ~(t[140]);
  assign t[81] = ~(t[141] & t[106]);
  assign t[82] = ~(x[4] & t[52]);
  assign t[83] = ~(t[141]);
  assign t[84] = ~(t[80]);
  assign t[85] = t[138] ? t[108] : t[107];
  assign t[86] = t[138] ? t[110] : t[109];
  assign t[87] = t[138] ? t[111] : t[81];
  assign t[88] = t[138] ? t[109] : t[110];
  assign t[89] = ~(t[157]);
  assign t[8] = ~(t[140] & t[141]);
  assign t[90] = ~(t[149] | t[150]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[112] & t[113]);
  assign t[93] = ~(t[158]);
  assign t[94] = ~(t[151] | t[152]);
  assign t[95] = ~(t[159]);
  assign t[96] = ~(t[160]);
  assign t[97] = ~(t[114] | t[115]);
  assign t[98] = ~(t[54] | t[116]);
  assign t[99] = ~(t[117] | t[118]);
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [97:0] x;
 output y;

 wire [339:0] t;
  assign t[0] = t[1] ? t[2] : t[137];
  assign t[100] = ~(t[161]);
  assign t[101] = ~(t[154] | t[155]);
  assign t[102] = ~(t[162]);
  assign t[103] = ~(t[163]);
  assign t[104] = ~(t[119] | t[120]);
  assign t[105] = ~(t[121] | t[57]);
  assign t[106] = ~(x[4] | t[122]);
  assign t[107] = ~(t[123] & t[141]);
  assign t[108] = ~(t[124] & t[83]);
  assign t[109] = ~(t[123] & t[83]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = ~(t[124] & t[141]);
  assign t[111] = ~(x[4] & t[125]);
  assign t[112] = ~(t[117]);
  assign t[113] = t[80] | t[126];
  assign t[114] = ~(t[164]);
  assign t[115] = ~(t[159] | t[160]);
  assign t[116] = ~(t[127] & t[128]);
  assign t[117] = ~(t[80] | t[129]);
  assign t[118] = t[55] | t[130];
  assign t[119] = ~(t[165]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = ~(t[162] | t[163]);
  assign t[121] = ~(t[84] | t[131]);
  assign t[122] = ~(t[139]);
  assign t[123] = x[4] & t[139];
  assign t[124] = ~(x[4] | t[139]);
  assign t[125] = ~(t[139] | t[141]);
  assign t[126] = t[138] ? t[111] : t[132];
  assign t[127] = ~(t[133] | t[56]);
  assign t[128] = ~(t[134] & t[135]);
  assign t[129] = t[138] ? t[132] : t[111];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = ~(t[31]);
  assign t[131] = t[138] ? t[82] : t[132];
  assign t[132] = ~(t[106] & t[83]);
  assign t[133] = ~(t[84] | t[136]);
  assign t[134] = t[141] & t[50];
  assign t[135] = t[124] | t[123];
  assign t[136] = t[138] ? t[107] : t[108];
  assign t[137] = (t[166]);
  assign t[138] = (t[167]);
  assign t[139] = (t[168]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (t[169]);
  assign t[141] = (t[170]);
  assign t[142] = (t[171]);
  assign t[143] = (t[172]);
  assign t[144] = (t[173]);
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = t[140] ? x[19] : x[18];
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = t[195] ^ x[2];
  assign t[167] = t[196] ^ x[8];
  assign t[168] = t[197] ^ x[11];
  assign t[169] = t[198] ^ x[14];
  assign t[16] = t[21] | t[22];
  assign t[170] = t[199] ^ x[17];
  assign t[171] = t[200] ^ x[22];
  assign t[172] = t[201] ^ x[25];
  assign t[173] = t[202] ^ x[28];
  assign t[174] = t[203] ^ x[31];
  assign t[175] = t[204] ^ x[36];
  assign t[176] = t[205] ^ x[39];
  assign t[177] = t[206] ^ x[42];
  assign t[178] = t[207] ^ x[45];
  assign t[179] = t[208] ^ x[48];
  assign t[17] = ~(t[23] | t[24]);
  assign t[180] = t[209] ^ x[51];
  assign t[181] = t[210] ^ x[54];
  assign t[182] = t[211] ^ x[57];
  assign t[183] = t[212] ^ x[62];
  assign t[184] = t[213] ^ x[65];
  assign t[185] = t[214] ^ x[68];
  assign t[186] = t[215] ^ x[73];
  assign t[187] = t[216] ^ x[76];
  assign t[188] = t[217] ^ x[79];
  assign t[189] = t[218] ^ x[82];
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = t[219] ^ x[85];
  assign t[191] = t[220] ^ x[88];
  assign t[192] = t[221] ^ x[91];
  assign t[193] = t[222] ^ x[94];
  assign t[194] = t[223] ^ x[97];
  assign t[195] = (t[224] & ~t[225]);
  assign t[196] = (t[226] & ~t[227]);
  assign t[197] = (t[228] & ~t[229]);
  assign t[198] = (t[230] & ~t[231]);
  assign t[199] = (t[232] & ~t[233]);
  assign t[19] = x[4] ? t[28] : t[27];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[234] & ~t[235]);
  assign t[201] = (t[236] & ~t[237]);
  assign t[202] = (t[238] & ~t[239]);
  assign t[203] = (t[240] & ~t[241]);
  assign t[204] = (t[242] & ~t[243]);
  assign t[205] = (t[244] & ~t[245]);
  assign t[206] = (t[246] & ~t[247]);
  assign t[207] = (t[248] & ~t[249]);
  assign t[208] = (t[250] & ~t[251]);
  assign t[209] = (t[252] & ~t[253]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[210] = (t[254] & ~t[255]);
  assign t[211] = (t[256] & ~t[257]);
  assign t[212] = (t[258] & ~t[259]);
  assign t[213] = (t[260] & ~t[261]);
  assign t[214] = (t[262] & ~t[263]);
  assign t[215] = (t[264] & ~t[265]);
  assign t[216] = (t[266] & ~t[267]);
  assign t[217] = (t[268] & ~t[269]);
  assign t[218] = (t[270] & ~t[271]);
  assign t[219] = (t[272] & ~t[273]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[274] & ~t[275]);
  assign t[221] = (t[276] & ~t[277]);
  assign t[222] = (t[278] & ~t[279]);
  assign t[223] = (t[280] & ~t[281]);
  assign t[224] = t[282] ^ x[2];
  assign t[225] = t[283] ^ x[1];
  assign t[226] = t[284] ^ x[8];
  assign t[227] = t[285] ^ x[7];
  assign t[228] = t[286] ^ x[11];
  assign t[229] = t[287] ^ x[10];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[288] ^ x[14];
  assign t[231] = t[289] ^ x[13];
  assign t[232] = t[290] ^ x[17];
  assign t[233] = t[291] ^ x[16];
  assign t[234] = t[292] ^ x[22];
  assign t[235] = t[293] ^ x[21];
  assign t[236] = t[294] ^ x[25];
  assign t[237] = t[295] ^ x[24];
  assign t[238] = t[296] ^ x[28];
  assign t[239] = t[297] ^ x[27];
  assign t[23] = ~(t[35] | t[36]);
  assign t[240] = t[298] ^ x[31];
  assign t[241] = t[299] ^ x[30];
  assign t[242] = t[300] ^ x[36];
  assign t[243] = t[301] ^ x[35];
  assign t[244] = t[302] ^ x[39];
  assign t[245] = t[303] ^ x[38];
  assign t[246] = t[304] ^ x[42];
  assign t[247] = t[305] ^ x[41];
  assign t[248] = t[306] ^ x[45];
  assign t[249] = t[307] ^ x[44];
  assign t[24] = ~(t[142] | t[37]);
  assign t[250] = t[308] ^ x[48];
  assign t[251] = t[309] ^ x[47];
  assign t[252] = t[310] ^ x[51];
  assign t[253] = t[311] ^ x[50];
  assign t[254] = t[312] ^ x[54];
  assign t[255] = t[313] ^ x[53];
  assign t[256] = t[314] ^ x[57];
  assign t[257] = t[315] ^ x[56];
  assign t[258] = t[316] ^ x[62];
  assign t[259] = t[317] ^ x[61];
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = t[318] ^ x[65];
  assign t[261] = t[319] ^ x[64];
  assign t[262] = t[320] ^ x[68];
  assign t[263] = t[321] ^ x[67];
  assign t[264] = t[322] ^ x[73];
  assign t[265] = t[323] ^ x[72];
  assign t[266] = t[324] ^ x[76];
  assign t[267] = t[325] ^ x[75];
  assign t[268] = t[326] ^ x[79];
  assign t[269] = t[327] ^ x[78];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[328] ^ x[82];
  assign t[271] = t[329] ^ x[81];
  assign t[272] = t[330] ^ x[85];
  assign t[273] = t[331] ^ x[84];
  assign t[274] = t[332] ^ x[88];
  assign t[275] = t[333] ^ x[87];
  assign t[276] = t[334] ^ x[91];
  assign t[277] = t[335] ^ x[90];
  assign t[278] = t[336] ^ x[94];
  assign t[279] = t[337] ^ x[93];
  assign t[27] = ~(t[42] | t[43]);
  assign t[280] = t[338] ^ x[97];
  assign t[281] = t[339] ^ x[96];
  assign t[282] = (x[0]);
  assign t[283] = (x[0]);
  assign t[284] = (x[6]);
  assign t[285] = (x[6]);
  assign t[286] = (x[9]);
  assign t[287] = (x[9]);
  assign t[288] = (x[12]);
  assign t[289] = (x[12]);
  assign t[28] = ~(t[44] ^ t[45]);
  assign t[290] = (x[15]);
  assign t[291] = (x[15]);
  assign t[292] = (x[20]);
  assign t[293] = (x[20]);
  assign t[294] = (x[23]);
  assign t[295] = (x[23]);
  assign t[296] = (x[26]);
  assign t[297] = (x[26]);
  assign t[298] = (x[29]);
  assign t[299] = (x[29]);
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[34]);
  assign t[301] = (x[34]);
  assign t[302] = (x[37]);
  assign t[303] = (x[37]);
  assign t[304] = (x[40]);
  assign t[305] = (x[40]);
  assign t[306] = (x[43]);
  assign t[307] = (x[43]);
  assign t[308] = (x[46]);
  assign t[309] = (x[46]);
  assign t[30] = ~(t[48] ^ t[49]);
  assign t[310] = (x[49]);
  assign t[311] = (x[49]);
  assign t[312] = (x[52]);
  assign t[313] = (x[52]);
  assign t[314] = (x[55]);
  assign t[315] = (x[55]);
  assign t[316] = (x[60]);
  assign t[317] = (x[60]);
  assign t[318] = (x[63]);
  assign t[319] = (x[63]);
  assign t[31] = ~(t[50] & t[51]);
  assign t[320] = (x[66]);
  assign t[321] = (x[66]);
  assign t[322] = (x[71]);
  assign t[323] = (x[71]);
  assign t[324] = (x[74]);
  assign t[325] = (x[74]);
  assign t[326] = (x[77]);
  assign t[327] = (x[77]);
  assign t[328] = (x[80]);
  assign t[329] = (x[80]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (x[83]);
  assign t[331] = (x[83]);
  assign t[332] = (x[86]);
  assign t[333] = (x[86]);
  assign t[334] = (x[89]);
  assign t[335] = (x[89]);
  assign t[336] = (x[92]);
  assign t[337] = (x[92]);
  assign t[338] = (x[95]);
  assign t[339] = (x[95]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[143]);
  assign t[36] = ~(t[144]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] | t[61]);
  assign t[39] = ~(t[145] | t[62]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[63] ? x[33] : x[32];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = ~(t[66] | t[67]);
  assign t[43] = ~(t[146] | t[68]);
  assign t[44] = ~(t[69] | t[70]);
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = ~(t[73] | t[74]);
  assign t[47] = ~(t[147] | t[75]);
  assign t[48] = ~(t[76] | t[77]);
  assign t[49] = ~(t[78] ^ t[79]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[80] | t[138]);
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = ~(t[139] | t[83]);
  assign t[53] = t[84] & t[138];
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[84] | t[86]);
  assign t[56] = ~(t[84] | t[87]);
  assign t[57] = ~(t[84] | t[88]);
  assign t[58] = ~(t[148]);
  assign t[59] = ~(t[143] | t[144]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[149]);
  assign t[61] = ~(t[150]);
  assign t[62] = ~(t[89] | t[90]);
  assign t[63] = ~(t[91]);
  assign t[64] = ~(t[21] | t[92]);
  assign t[65] = ~(t[54]);
  assign t[66] = ~(t[151]);
  assign t[67] = ~(t[152]);
  assign t[68] = ~(t[93] | t[94]);
  assign t[69] = ~(t[95] | t[96]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[153] | t[97]);
  assign t[71] = t[140] ? x[59] : x[58];
  assign t[72] = ~(t[98] & t[99]);
  assign t[73] = ~(t[154]);
  assign t[74] = ~(t[155]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[102] | t[103]);
  assign t[77] = ~(t[156] | t[104]);
  assign t[78] = t[140] ? x[70] : x[69];
  assign t[79] = ~(t[98] & t[105]);
  assign t[7] = ~(t[138] & t[139]);
  assign t[80] = ~(t[140]);
  assign t[81] = ~(t[141] & t[106]);
  assign t[82] = ~(x[4] & t[52]);
  assign t[83] = ~(t[141]);
  assign t[84] = ~(t[80]);
  assign t[85] = t[138] ? t[108] : t[107];
  assign t[86] = t[138] ? t[110] : t[109];
  assign t[87] = t[138] ? t[111] : t[81];
  assign t[88] = t[138] ? t[109] : t[110];
  assign t[89] = ~(t[157]);
  assign t[8] = ~(t[140] & t[141]);
  assign t[90] = ~(t[149] | t[150]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[112] & t[113]);
  assign t[93] = ~(t[158]);
  assign t[94] = ~(t[151] | t[152]);
  assign t[95] = ~(t[159]);
  assign t[96] = ~(t[160]);
  assign t[97] = ~(t[114] | t[115]);
  assign t[98] = ~(t[54] | t[116]);
  assign t[99] = ~(t[117] | t[118]);
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [79:0] x;
 output y;

 wire [221:0] t;
  assign t[0] = t[1] ? t[2] : t[61];
  assign t[100] = t[123] ^ x[61];
  assign t[101] = t[124] ^ x[64];
  assign t[102] = t[125] ^ x[67];
  assign t[103] = t[126] ^ x[70];
  assign t[104] = t[127] ^ x[73];
  assign t[105] = t[128] ^ x[76];
  assign t[106] = t[129] ^ x[79];
  assign t[107] = (t[130] & ~t[131]);
  assign t[108] = (t[132] & ~t[133]);
  assign t[109] = (t[134] & ~t[135]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = (t[136] & ~t[137]);
  assign t[111] = (t[138] & ~t[139]);
  assign t[112] = (t[140] & ~t[141]);
  assign t[113] = (t[142] & ~t[143]);
  assign t[114] = (t[144] & ~t[145]);
  assign t[115] = (t[146] & ~t[147]);
  assign t[116] = (t[148] & ~t[149]);
  assign t[117] = (t[150] & ~t[151]);
  assign t[118] = (t[152] & ~t[153]);
  assign t[119] = (t[154] & ~t[155]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[156] & ~t[157]);
  assign t[121] = (t[158] & ~t[159]);
  assign t[122] = (t[160] & ~t[161]);
  assign t[123] = (t[162] & ~t[163]);
  assign t[124] = (t[164] & ~t[165]);
  assign t[125] = (t[166] & ~t[167]);
  assign t[126] = (t[168] & ~t[169]);
  assign t[127] = (t[170] & ~t[171]);
  assign t[128] = (t[172] & ~t[173]);
  assign t[129] = (t[174] & ~t[175]);
  assign t[12] = t[64] ? x[19] : x[18];
  assign t[130] = t[176] ^ x[2];
  assign t[131] = t[177] ^ x[1];
  assign t[132] = t[178] ^ x[8];
  assign t[133] = t[179] ^ x[7];
  assign t[134] = t[180] ^ x[11];
  assign t[135] = t[181] ^ x[10];
  assign t[136] = t[182] ^ x[14];
  assign t[137] = t[183] ^ x[13];
  assign t[138] = t[184] ^ x[17];
  assign t[139] = t[185] ^ x[16];
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = t[186] ^ x[22];
  assign t[141] = t[187] ^ x[21];
  assign t[142] = t[188] ^ x[25];
  assign t[143] = t[189] ^ x[24];
  assign t[144] = t[190] ^ x[30];
  assign t[145] = t[191] ^ x[29];
  assign t[146] = t[192] ^ x[33];
  assign t[147] = t[193] ^ x[32];
  assign t[148] = t[194] ^ x[36];
  assign t[149] = t[195] ^ x[35];
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = t[196] ^ x[39];
  assign t[151] = t[197] ^ x[38];
  assign t[152] = t[198] ^ x[42];
  assign t[153] = t[199] ^ x[41];
  assign t[154] = t[200] ^ x[47];
  assign t[155] = t[201] ^ x[46];
  assign t[156] = t[202] ^ x[50];
  assign t[157] = t[203] ^ x[49];
  assign t[158] = t[204] ^ x[55];
  assign t[159] = t[205] ^ x[54];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[206] ^ x[58];
  assign t[161] = t[207] ^ x[57];
  assign t[162] = t[208] ^ x[61];
  assign t[163] = t[209] ^ x[60];
  assign t[164] = t[210] ^ x[64];
  assign t[165] = t[211] ^ x[63];
  assign t[166] = t[212] ^ x[67];
  assign t[167] = t[213] ^ x[66];
  assign t[168] = t[214] ^ x[70];
  assign t[169] = t[215] ^ x[69];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[216] ^ x[73];
  assign t[171] = t[217] ^ x[72];
  assign t[172] = t[218] ^ x[76];
  assign t[173] = t[219] ^ x[75];
  assign t[174] = t[220] ^ x[79];
  assign t[175] = t[221] ^ x[78];
  assign t[176] = (x[0]);
  assign t[177] = (x[0]);
  assign t[178] = (x[6]);
  assign t[179] = (x[6]);
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = (x[9]);
  assign t[181] = (x[9]);
  assign t[182] = (x[12]);
  assign t[183] = (x[12]);
  assign t[184] = (x[15]);
  assign t[185] = (x[15]);
  assign t[186] = (x[20]);
  assign t[187] = (x[20]);
  assign t[188] = (x[23]);
  assign t[189] = (x[23]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[28]);
  assign t[191] = (x[28]);
  assign t[192] = (x[31]);
  assign t[193] = (x[31]);
  assign t[194] = (x[34]);
  assign t[195] = (x[34]);
  assign t[196] = (x[37]);
  assign t[197] = (x[37]);
  assign t[198] = (x[40]);
  assign t[199] = (x[40]);
  assign t[19] = ~(t[66] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (x[45]);
  assign t[201] = (x[45]);
  assign t[202] = (x[48]);
  assign t[203] = (x[48]);
  assign t[204] = (x[53]);
  assign t[205] = (x[53]);
  assign t[206] = (x[56]);
  assign t[207] = (x[56]);
  assign t[208] = (x[59]);
  assign t[209] = (x[59]);
  assign t[20] = ~(t[67] & t[28]);
  assign t[210] = (x[62]);
  assign t[211] = (x[62]);
  assign t[212] = (x[65]);
  assign t[213] = (x[65]);
  assign t[214] = (x[68]);
  assign t[215] = (x[68]);
  assign t[216] = (x[71]);
  assign t[217] = (x[71]);
  assign t[218] = (x[74]);
  assign t[219] = (x[74]);
  assign t[21] = t[64] ? x[27] : x[26];
  assign t[220] = (x[77]);
  assign t[221] = (x[77]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[35] & t[36]);
  assign t[26] = t[37] ^ t[38];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[68] & t[39]);
  assign t[29] = ~(t[69] & t[40]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[70] & t[41]);
  assign t[31] = ~(t[71] & t[42]);
  assign t[32] = ~(t[72] & t[43]);
  assign t[33] = t[64] ? x[44] : x[43];
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[73] & t[46]);
  assign t[36] = ~(t[74] & t[47]);
  assign t[37] = t[48] ? x[52] : x[51];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[66]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[75]);
  assign t[41] = ~(t[75] & t[51]);
  assign t[42] = ~(t[76]);
  assign t[43] = ~(t[76] & t[52]);
  assign t[44] = ~(t[77] & t[53]);
  assign t[45] = ~(t[78] & t[54]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[55]);
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[69]);
  assign t[52] = ~(t[71]);
  assign t[53] = ~(t[82]);
  assign t[54] = ~(t[82] & t[59]);
  assign t[55] = ~(t[73]);
  assign t[56] = ~(t[64]);
  assign t[57] = ~(t[83]);
  assign t[58] = ~(t[83] & t[60]);
  assign t[59] = ~(t[77]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[80]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = (t[86]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = ~(t[62] & t[63]);
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = t[107] ^ x[2];
  assign t[85] = t[108] ^ x[8];
  assign t[86] = t[109] ^ x[11];
  assign t[87] = t[110] ^ x[14];
  assign t[88] = t[111] ^ x[17];
  assign t[89] = t[112] ^ x[22];
  assign t[8] = ~(t[64] & t[65]);
  assign t[90] = t[113] ^ x[25];
  assign t[91] = t[114] ^ x[30];
  assign t[92] = t[115] ^ x[33];
  assign t[93] = t[116] ^ x[36];
  assign t[94] = t[117] ^ x[39];
  assign t[95] = t[118] ^ x[42];
  assign t[96] = t[119] ^ x[47];
  assign t[97] = t[120] ^ x[50];
  assign t[98] = t[121] ^ x[55];
  assign t[99] = t[122] ^ x[58];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [79:0] x;
 output y;

 wire [221:0] t;
  assign t[0] = t[1] ? t[2] : t[61];
  assign t[100] = t[123] ^ x[61];
  assign t[101] = t[124] ^ x[64];
  assign t[102] = t[125] ^ x[67];
  assign t[103] = t[126] ^ x[70];
  assign t[104] = t[127] ^ x[73];
  assign t[105] = t[128] ^ x[76];
  assign t[106] = t[129] ^ x[79];
  assign t[107] = (t[130] & ~t[131]);
  assign t[108] = (t[132] & ~t[133]);
  assign t[109] = (t[134] & ~t[135]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = (t[136] & ~t[137]);
  assign t[111] = (t[138] & ~t[139]);
  assign t[112] = (t[140] & ~t[141]);
  assign t[113] = (t[142] & ~t[143]);
  assign t[114] = (t[144] & ~t[145]);
  assign t[115] = (t[146] & ~t[147]);
  assign t[116] = (t[148] & ~t[149]);
  assign t[117] = (t[150] & ~t[151]);
  assign t[118] = (t[152] & ~t[153]);
  assign t[119] = (t[154] & ~t[155]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[156] & ~t[157]);
  assign t[121] = (t[158] & ~t[159]);
  assign t[122] = (t[160] & ~t[161]);
  assign t[123] = (t[162] & ~t[163]);
  assign t[124] = (t[164] & ~t[165]);
  assign t[125] = (t[166] & ~t[167]);
  assign t[126] = (t[168] & ~t[169]);
  assign t[127] = (t[170] & ~t[171]);
  assign t[128] = (t[172] & ~t[173]);
  assign t[129] = (t[174] & ~t[175]);
  assign t[12] = t[64] ? x[19] : x[18];
  assign t[130] = t[176] ^ x[2];
  assign t[131] = t[177] ^ x[1];
  assign t[132] = t[178] ^ x[8];
  assign t[133] = t[179] ^ x[7];
  assign t[134] = t[180] ^ x[11];
  assign t[135] = t[181] ^ x[10];
  assign t[136] = t[182] ^ x[14];
  assign t[137] = t[183] ^ x[13];
  assign t[138] = t[184] ^ x[17];
  assign t[139] = t[185] ^ x[16];
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = t[186] ^ x[22];
  assign t[141] = t[187] ^ x[21];
  assign t[142] = t[188] ^ x[25];
  assign t[143] = t[189] ^ x[24];
  assign t[144] = t[190] ^ x[30];
  assign t[145] = t[191] ^ x[29];
  assign t[146] = t[192] ^ x[33];
  assign t[147] = t[193] ^ x[32];
  assign t[148] = t[194] ^ x[36];
  assign t[149] = t[195] ^ x[35];
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = t[196] ^ x[39];
  assign t[151] = t[197] ^ x[38];
  assign t[152] = t[198] ^ x[42];
  assign t[153] = t[199] ^ x[41];
  assign t[154] = t[200] ^ x[47];
  assign t[155] = t[201] ^ x[46];
  assign t[156] = t[202] ^ x[50];
  assign t[157] = t[203] ^ x[49];
  assign t[158] = t[204] ^ x[55];
  assign t[159] = t[205] ^ x[54];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[206] ^ x[58];
  assign t[161] = t[207] ^ x[57];
  assign t[162] = t[208] ^ x[61];
  assign t[163] = t[209] ^ x[60];
  assign t[164] = t[210] ^ x[64];
  assign t[165] = t[211] ^ x[63];
  assign t[166] = t[212] ^ x[67];
  assign t[167] = t[213] ^ x[66];
  assign t[168] = t[214] ^ x[70];
  assign t[169] = t[215] ^ x[69];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[216] ^ x[73];
  assign t[171] = t[217] ^ x[72];
  assign t[172] = t[218] ^ x[76];
  assign t[173] = t[219] ^ x[75];
  assign t[174] = t[220] ^ x[79];
  assign t[175] = t[221] ^ x[78];
  assign t[176] = (x[0]);
  assign t[177] = (x[0]);
  assign t[178] = (x[6]);
  assign t[179] = (x[6]);
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = (x[9]);
  assign t[181] = (x[9]);
  assign t[182] = (x[12]);
  assign t[183] = (x[12]);
  assign t[184] = (x[15]);
  assign t[185] = (x[15]);
  assign t[186] = (x[20]);
  assign t[187] = (x[20]);
  assign t[188] = (x[23]);
  assign t[189] = (x[23]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[28]);
  assign t[191] = (x[28]);
  assign t[192] = (x[31]);
  assign t[193] = (x[31]);
  assign t[194] = (x[34]);
  assign t[195] = (x[34]);
  assign t[196] = (x[37]);
  assign t[197] = (x[37]);
  assign t[198] = (x[40]);
  assign t[199] = (x[40]);
  assign t[19] = ~(t[66] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (x[45]);
  assign t[201] = (x[45]);
  assign t[202] = (x[48]);
  assign t[203] = (x[48]);
  assign t[204] = (x[53]);
  assign t[205] = (x[53]);
  assign t[206] = (x[56]);
  assign t[207] = (x[56]);
  assign t[208] = (x[59]);
  assign t[209] = (x[59]);
  assign t[20] = ~(t[67] & t[28]);
  assign t[210] = (x[62]);
  assign t[211] = (x[62]);
  assign t[212] = (x[65]);
  assign t[213] = (x[65]);
  assign t[214] = (x[68]);
  assign t[215] = (x[68]);
  assign t[216] = (x[71]);
  assign t[217] = (x[71]);
  assign t[218] = (x[74]);
  assign t[219] = (x[74]);
  assign t[21] = t[64] ? x[27] : x[26];
  assign t[220] = (x[77]);
  assign t[221] = (x[77]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[35] & t[36]);
  assign t[26] = t[37] ^ t[38];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[68] & t[39]);
  assign t[29] = ~(t[69] & t[40]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[70] & t[41]);
  assign t[31] = ~(t[71] & t[42]);
  assign t[32] = ~(t[72] & t[43]);
  assign t[33] = t[64] ? x[44] : x[43];
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[73] & t[46]);
  assign t[36] = ~(t[74] & t[47]);
  assign t[37] = t[48] ? x[52] : x[51];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[66]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[75]);
  assign t[41] = ~(t[75] & t[51]);
  assign t[42] = ~(t[76]);
  assign t[43] = ~(t[76] & t[52]);
  assign t[44] = ~(t[77] & t[53]);
  assign t[45] = ~(t[78] & t[54]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[55]);
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[69]);
  assign t[52] = ~(t[71]);
  assign t[53] = ~(t[82]);
  assign t[54] = ~(t[82] & t[59]);
  assign t[55] = ~(t[73]);
  assign t[56] = ~(t[64]);
  assign t[57] = ~(t[83]);
  assign t[58] = ~(t[83] & t[60]);
  assign t[59] = ~(t[77]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[80]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = (t[86]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = ~(t[62] & t[63]);
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = t[107] ^ x[2];
  assign t[85] = t[108] ^ x[8];
  assign t[86] = t[109] ^ x[11];
  assign t[87] = t[110] ^ x[14];
  assign t[88] = t[111] ^ x[17];
  assign t[89] = t[112] ^ x[22];
  assign t[8] = ~(t[64] & t[65]);
  assign t[90] = t[113] ^ x[25];
  assign t[91] = t[114] ^ x[30];
  assign t[92] = t[115] ^ x[33];
  assign t[93] = t[116] ^ x[36];
  assign t[94] = t[117] ^ x[39];
  assign t[95] = t[118] ^ x[42];
  assign t[96] = t[119] ^ x[47];
  assign t[97] = t[120] ^ x[50];
  assign t[98] = t[121] ^ x[55];
  assign t[99] = t[122] ^ x[58];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [97:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = t[131] ^ x[2];
  assign t[103] = t[132] ^ x[8];
  assign t[104] = t[133] ^ x[11];
  assign t[105] = t[134] ^ x[14];
  assign t[106] = t[135] ^ x[17];
  assign t[107] = t[136] ^ x[22];
  assign t[108] = t[137] ^ x[27];
  assign t[109] = t[138] ^ x[30];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[33];
  assign t[111] = t[140] ^ x[36];
  assign t[112] = t[141] ^ x[41];
  assign t[113] = t[142] ^ x[46];
  assign t[114] = t[143] ^ x[49];
  assign t[115] = t[144] ^ x[52];
  assign t[116] = t[145] ^ x[55];
  assign t[117] = t[146] ^ x[58];
  assign t[118] = t[147] ^ x[61];
  assign t[119] = t[148] ^ x[64];
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[149] ^ x[67];
  assign t[121] = t[150] ^ x[70];
  assign t[122] = t[151] ^ x[73];
  assign t[123] = t[152] ^ x[76];
  assign t[124] = t[153] ^ x[79];
  assign t[125] = t[154] ^ x[82];
  assign t[126] = t[155] ^ x[85];
  assign t[127] = t[156] ^ x[88];
  assign t[128] = t[157] ^ x[91];
  assign t[129] = t[158] ^ x[94];
  assign t[12] = t[76] ? x[18] : x[19];
  assign t[130] = t[159] ^ x[97];
  assign t[131] = (t[160] & ~t[161]);
  assign t[132] = (t[162] & ~t[163]);
  assign t[133] = (t[164] & ~t[165]);
  assign t[134] = (t[166] & ~t[167]);
  assign t[135] = (t[168] & ~t[169]);
  assign t[136] = (t[170] & ~t[171]);
  assign t[137] = (t[172] & ~t[173]);
  assign t[138] = (t[174] & ~t[175]);
  assign t[139] = (t[176] & ~t[177]);
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = (t[178] & ~t[179]);
  assign t[141] = (t[180] & ~t[181]);
  assign t[142] = (t[182] & ~t[183]);
  assign t[143] = (t[184] & ~t[185]);
  assign t[144] = (t[186] & ~t[187]);
  assign t[145] = (t[188] & ~t[189]);
  assign t[146] = (t[190] & ~t[191]);
  assign t[147] = (t[192] & ~t[193]);
  assign t[148] = (t[194] & ~t[195]);
  assign t[149] = (t[196] & ~t[197]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (t[198] & ~t[199]);
  assign t[151] = (t[200] & ~t[201]);
  assign t[152] = (t[202] & ~t[203]);
  assign t[153] = (t[204] & ~t[205]);
  assign t[154] = (t[206] & ~t[207]);
  assign t[155] = (t[208] & ~t[209]);
  assign t[156] = (t[210] & ~t[211]);
  assign t[157] = (t[212] & ~t[213]);
  assign t[158] = (t[214] & ~t[215]);
  assign t[159] = (t[216] & ~t[217]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[218] ^ x[2];
  assign t[161] = t[219] ^ x[1];
  assign t[162] = t[220] ^ x[8];
  assign t[163] = t[221] ^ x[7];
  assign t[164] = t[222] ^ x[11];
  assign t[165] = t[223] ^ x[10];
  assign t[166] = t[224] ^ x[14];
  assign t[167] = t[225] ^ x[13];
  assign t[168] = t[226] ^ x[17];
  assign t[169] = t[227] ^ x[16];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[228] ^ x[22];
  assign t[171] = t[229] ^ x[21];
  assign t[172] = t[230] ^ x[27];
  assign t[173] = t[231] ^ x[26];
  assign t[174] = t[232] ^ x[30];
  assign t[175] = t[233] ^ x[29];
  assign t[176] = t[234] ^ x[33];
  assign t[177] = t[235] ^ x[32];
  assign t[178] = t[236] ^ x[36];
  assign t[179] = t[237] ^ x[35];
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = t[238] ^ x[41];
  assign t[181] = t[239] ^ x[40];
  assign t[182] = t[240] ^ x[46];
  assign t[183] = t[241] ^ x[45];
  assign t[184] = t[242] ^ x[49];
  assign t[185] = t[243] ^ x[48];
  assign t[186] = t[244] ^ x[52];
  assign t[187] = t[245] ^ x[51];
  assign t[188] = t[246] ^ x[55];
  assign t[189] = t[247] ^ x[54];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[248] ^ x[58];
  assign t[191] = t[249] ^ x[57];
  assign t[192] = t[250] ^ x[61];
  assign t[193] = t[251] ^ x[60];
  assign t[194] = t[252] ^ x[64];
  assign t[195] = t[253] ^ x[63];
  assign t[196] = t[254] ^ x[67];
  assign t[197] = t[255] ^ x[66];
  assign t[198] = t[256] ^ x[70];
  assign t[199] = t[257] ^ x[69];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[258] ^ x[73];
  assign t[201] = t[259] ^ x[72];
  assign t[202] = t[260] ^ x[76];
  assign t[203] = t[261] ^ x[75];
  assign t[204] = t[262] ^ x[79];
  assign t[205] = t[263] ^ x[78];
  assign t[206] = t[264] ^ x[82];
  assign t[207] = t[265] ^ x[81];
  assign t[208] = t[266] ^ x[85];
  assign t[209] = t[267] ^ x[84];
  assign t[20] = ~(t[29] & t[78]);
  assign t[210] = t[268] ^ x[88];
  assign t[211] = t[269] ^ x[87];
  assign t[212] = t[270] ^ x[91];
  assign t[213] = t[271] ^ x[90];
  assign t[214] = t[272] ^ x[94];
  assign t[215] = t[273] ^ x[93];
  assign t[216] = t[274] ^ x[97];
  assign t[217] = t[275] ^ x[96];
  assign t[218] = (x[0]);
  assign t[219] = (x[0]);
  assign t[21] = t[76] ? x[24] : x[23];
  assign t[220] = (x[6]);
  assign t[221] = (x[6]);
  assign t[222] = (x[9]);
  assign t[223] = (x[9]);
  assign t[224] = (x[12]);
  assign t[225] = (x[12]);
  assign t[226] = (x[15]);
  assign t[227] = (x[15]);
  assign t[228] = (x[20]);
  assign t[229] = (x[20]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[25]);
  assign t[231] = (x[25]);
  assign t[232] = (x[28]);
  assign t[233] = (x[28]);
  assign t[234] = (x[31]);
  assign t[235] = (x[31]);
  assign t[236] = (x[34]);
  assign t[237] = (x[34]);
  assign t[238] = (x[39]);
  assign t[239] = (x[39]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[240] = (x[44]);
  assign t[241] = (x[44]);
  assign t[242] = (x[47]);
  assign t[243] = (x[47]);
  assign t[244] = (x[50]);
  assign t[245] = (x[50]);
  assign t[246] = (x[53]);
  assign t[247] = (x[53]);
  assign t[248] = (x[56]);
  assign t[249] = (x[56]);
  assign t[24] = t[34] ^ t[35];
  assign t[250] = (x[59]);
  assign t[251] = (x[59]);
  assign t[252] = (x[62]);
  assign t[253] = (x[62]);
  assign t[254] = (x[65]);
  assign t[255] = (x[65]);
  assign t[256] = (x[68]);
  assign t[257] = (x[68]);
  assign t[258] = (x[71]);
  assign t[259] = (x[71]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[260] = (x[74]);
  assign t[261] = (x[74]);
  assign t[262] = (x[77]);
  assign t[263] = (x[77]);
  assign t[264] = (x[80]);
  assign t[265] = (x[80]);
  assign t[266] = (x[83]);
  assign t[267] = (x[83]);
  assign t[268] = (x[86]);
  assign t[269] = (x[86]);
  assign t[26] = t[38] ^ t[39];
  assign t[270] = (x[89]);
  assign t[271] = (x[89]);
  assign t[272] = (x[92]);
  assign t[273] = (x[92]);
  assign t[274] = (x[95]);
  assign t[275] = (x[95]);
  assign t[27] = ~(t[79]);
  assign t[28] = ~(t[80]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = ~(t[44] & t[81]);
  assign t[32] = ~(t[45] & t[46]);
  assign t[33] = ~(t[47] & t[82]);
  assign t[34] = t[76] ? x[38] : x[37];
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[52] & t[83]);
  assign t[38] = t[53] ? x[43] : x[42];
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[80] & t[79]);
  assign t[41] = ~(t[84]);
  assign t[42] = ~(t[85]);
  assign t[43] = ~(t[86]);
  assign t[44] = ~(t[56] & t[57]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[58] & t[59]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[62] & t[89]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[90]);
  assign t[51] = ~(t[91]);
  assign t[52] = ~(t[63] & t[64]);
  assign t[53] = ~(t[65]);
  assign t[54] = ~(t[66] & t[67]);
  assign t[55] = ~(t[68] & t[92]);
  assign t[56] = ~(t[86] & t[85]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[88] & t[87]);
  assign t[59] = ~(t[94]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[69] & t[70]);
  assign t[63] = ~(t[91] & t[90]);
  assign t[64] = ~(t[97]);
  assign t[65] = ~(t[76]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[99]);
  assign t[68] = ~(t[71] & t[72]);
  assign t[69] = ~(t[96] & t[95]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[100]);
  assign t[71] = ~(t[99] & t[98]);
  assign t[72] = ~(t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[74] & t[75]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[76] & t[77]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind161(x, y);
 input [97:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = t[131] ^ x[2];
  assign t[103] = t[132] ^ x[8];
  assign t[104] = t[133] ^ x[11];
  assign t[105] = t[134] ^ x[14];
  assign t[106] = t[135] ^ x[17];
  assign t[107] = t[136] ^ x[22];
  assign t[108] = t[137] ^ x[27];
  assign t[109] = t[138] ^ x[30];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[33];
  assign t[111] = t[140] ^ x[36];
  assign t[112] = t[141] ^ x[41];
  assign t[113] = t[142] ^ x[46];
  assign t[114] = t[143] ^ x[49];
  assign t[115] = t[144] ^ x[52];
  assign t[116] = t[145] ^ x[55];
  assign t[117] = t[146] ^ x[58];
  assign t[118] = t[147] ^ x[61];
  assign t[119] = t[148] ^ x[64];
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[149] ^ x[67];
  assign t[121] = t[150] ^ x[70];
  assign t[122] = t[151] ^ x[73];
  assign t[123] = t[152] ^ x[76];
  assign t[124] = t[153] ^ x[79];
  assign t[125] = t[154] ^ x[82];
  assign t[126] = t[155] ^ x[85];
  assign t[127] = t[156] ^ x[88];
  assign t[128] = t[157] ^ x[91];
  assign t[129] = t[158] ^ x[94];
  assign t[12] = t[76] ? x[18] : x[19];
  assign t[130] = t[159] ^ x[97];
  assign t[131] = (t[160] & ~t[161]);
  assign t[132] = (t[162] & ~t[163]);
  assign t[133] = (t[164] & ~t[165]);
  assign t[134] = (t[166] & ~t[167]);
  assign t[135] = (t[168] & ~t[169]);
  assign t[136] = (t[170] & ~t[171]);
  assign t[137] = (t[172] & ~t[173]);
  assign t[138] = (t[174] & ~t[175]);
  assign t[139] = (t[176] & ~t[177]);
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = (t[178] & ~t[179]);
  assign t[141] = (t[180] & ~t[181]);
  assign t[142] = (t[182] & ~t[183]);
  assign t[143] = (t[184] & ~t[185]);
  assign t[144] = (t[186] & ~t[187]);
  assign t[145] = (t[188] & ~t[189]);
  assign t[146] = (t[190] & ~t[191]);
  assign t[147] = (t[192] & ~t[193]);
  assign t[148] = (t[194] & ~t[195]);
  assign t[149] = (t[196] & ~t[197]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (t[198] & ~t[199]);
  assign t[151] = (t[200] & ~t[201]);
  assign t[152] = (t[202] & ~t[203]);
  assign t[153] = (t[204] & ~t[205]);
  assign t[154] = (t[206] & ~t[207]);
  assign t[155] = (t[208] & ~t[209]);
  assign t[156] = (t[210] & ~t[211]);
  assign t[157] = (t[212] & ~t[213]);
  assign t[158] = (t[214] & ~t[215]);
  assign t[159] = (t[216] & ~t[217]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[218] ^ x[2];
  assign t[161] = t[219] ^ x[1];
  assign t[162] = t[220] ^ x[8];
  assign t[163] = t[221] ^ x[7];
  assign t[164] = t[222] ^ x[11];
  assign t[165] = t[223] ^ x[10];
  assign t[166] = t[224] ^ x[14];
  assign t[167] = t[225] ^ x[13];
  assign t[168] = t[226] ^ x[17];
  assign t[169] = t[227] ^ x[16];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[228] ^ x[22];
  assign t[171] = t[229] ^ x[21];
  assign t[172] = t[230] ^ x[27];
  assign t[173] = t[231] ^ x[26];
  assign t[174] = t[232] ^ x[30];
  assign t[175] = t[233] ^ x[29];
  assign t[176] = t[234] ^ x[33];
  assign t[177] = t[235] ^ x[32];
  assign t[178] = t[236] ^ x[36];
  assign t[179] = t[237] ^ x[35];
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = t[238] ^ x[41];
  assign t[181] = t[239] ^ x[40];
  assign t[182] = t[240] ^ x[46];
  assign t[183] = t[241] ^ x[45];
  assign t[184] = t[242] ^ x[49];
  assign t[185] = t[243] ^ x[48];
  assign t[186] = t[244] ^ x[52];
  assign t[187] = t[245] ^ x[51];
  assign t[188] = t[246] ^ x[55];
  assign t[189] = t[247] ^ x[54];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[248] ^ x[58];
  assign t[191] = t[249] ^ x[57];
  assign t[192] = t[250] ^ x[61];
  assign t[193] = t[251] ^ x[60];
  assign t[194] = t[252] ^ x[64];
  assign t[195] = t[253] ^ x[63];
  assign t[196] = t[254] ^ x[67];
  assign t[197] = t[255] ^ x[66];
  assign t[198] = t[256] ^ x[70];
  assign t[199] = t[257] ^ x[69];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[258] ^ x[73];
  assign t[201] = t[259] ^ x[72];
  assign t[202] = t[260] ^ x[76];
  assign t[203] = t[261] ^ x[75];
  assign t[204] = t[262] ^ x[79];
  assign t[205] = t[263] ^ x[78];
  assign t[206] = t[264] ^ x[82];
  assign t[207] = t[265] ^ x[81];
  assign t[208] = t[266] ^ x[85];
  assign t[209] = t[267] ^ x[84];
  assign t[20] = ~(t[29] & t[78]);
  assign t[210] = t[268] ^ x[88];
  assign t[211] = t[269] ^ x[87];
  assign t[212] = t[270] ^ x[91];
  assign t[213] = t[271] ^ x[90];
  assign t[214] = t[272] ^ x[94];
  assign t[215] = t[273] ^ x[93];
  assign t[216] = t[274] ^ x[97];
  assign t[217] = t[275] ^ x[96];
  assign t[218] = (x[0]);
  assign t[219] = (x[0]);
  assign t[21] = t[76] ? x[24] : x[23];
  assign t[220] = (x[6]);
  assign t[221] = (x[6]);
  assign t[222] = (x[9]);
  assign t[223] = (x[9]);
  assign t[224] = (x[12]);
  assign t[225] = (x[12]);
  assign t[226] = (x[15]);
  assign t[227] = (x[15]);
  assign t[228] = (x[20]);
  assign t[229] = (x[20]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[25]);
  assign t[231] = (x[25]);
  assign t[232] = (x[28]);
  assign t[233] = (x[28]);
  assign t[234] = (x[31]);
  assign t[235] = (x[31]);
  assign t[236] = (x[34]);
  assign t[237] = (x[34]);
  assign t[238] = (x[39]);
  assign t[239] = (x[39]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[240] = (x[44]);
  assign t[241] = (x[44]);
  assign t[242] = (x[47]);
  assign t[243] = (x[47]);
  assign t[244] = (x[50]);
  assign t[245] = (x[50]);
  assign t[246] = (x[53]);
  assign t[247] = (x[53]);
  assign t[248] = (x[56]);
  assign t[249] = (x[56]);
  assign t[24] = t[34] ^ t[35];
  assign t[250] = (x[59]);
  assign t[251] = (x[59]);
  assign t[252] = (x[62]);
  assign t[253] = (x[62]);
  assign t[254] = (x[65]);
  assign t[255] = (x[65]);
  assign t[256] = (x[68]);
  assign t[257] = (x[68]);
  assign t[258] = (x[71]);
  assign t[259] = (x[71]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[260] = (x[74]);
  assign t[261] = (x[74]);
  assign t[262] = (x[77]);
  assign t[263] = (x[77]);
  assign t[264] = (x[80]);
  assign t[265] = (x[80]);
  assign t[266] = (x[83]);
  assign t[267] = (x[83]);
  assign t[268] = (x[86]);
  assign t[269] = (x[86]);
  assign t[26] = t[38] ^ t[39];
  assign t[270] = (x[89]);
  assign t[271] = (x[89]);
  assign t[272] = (x[92]);
  assign t[273] = (x[92]);
  assign t[274] = (x[95]);
  assign t[275] = (x[95]);
  assign t[27] = ~(t[79]);
  assign t[28] = ~(t[80]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = ~(t[44] & t[81]);
  assign t[32] = ~(t[45] & t[46]);
  assign t[33] = ~(t[47] & t[82]);
  assign t[34] = t[76] ? x[38] : x[37];
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[52] & t[83]);
  assign t[38] = t[53] ? x[43] : x[42];
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[80] & t[79]);
  assign t[41] = ~(t[84]);
  assign t[42] = ~(t[85]);
  assign t[43] = ~(t[86]);
  assign t[44] = ~(t[56] & t[57]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[58] & t[59]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[62] & t[89]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[90]);
  assign t[51] = ~(t[91]);
  assign t[52] = ~(t[63] & t[64]);
  assign t[53] = ~(t[65]);
  assign t[54] = ~(t[66] & t[67]);
  assign t[55] = ~(t[68] & t[92]);
  assign t[56] = ~(t[86] & t[85]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[88] & t[87]);
  assign t[59] = ~(t[94]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[69] & t[70]);
  assign t[63] = ~(t[91] & t[90]);
  assign t[64] = ~(t[97]);
  assign t[65] = ~(t[76]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[99]);
  assign t[68] = ~(t[71] & t[72]);
  assign t[69] = ~(t[96] & t[95]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[100]);
  assign t[71] = ~(t[99] & t[98]);
  assign t[72] = ~(t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[74] & t[75]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[76] & t[77]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [97:0] x;
 output y;

 wire [269:0] t;
  assign t[0] = t[1] ? t[2] : t[67];
  assign t[100] = t[129] ^ x[17];
  assign t[101] = t[130] ^ x[22];
  assign t[102] = t[131] ^ x[27];
  assign t[103] = t[132] ^ x[30];
  assign t[104] = t[133] ^ x[33];
  assign t[105] = t[134] ^ x[36];
  assign t[106] = t[135] ^ x[41];
  assign t[107] = t[136] ^ x[46];
  assign t[108] = t[137] ^ x[49];
  assign t[109] = t[138] ^ x[52];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[55];
  assign t[111] = t[140] ^ x[58];
  assign t[112] = t[141] ^ x[61];
  assign t[113] = t[142] ^ x[64];
  assign t[114] = t[143] ^ x[67];
  assign t[115] = t[144] ^ x[70];
  assign t[116] = t[145] ^ x[73];
  assign t[117] = t[146] ^ x[76];
  assign t[118] = t[147] ^ x[79];
  assign t[119] = t[148] ^ x[82];
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[149] ^ x[85];
  assign t[121] = t[150] ^ x[88];
  assign t[122] = t[151] ^ x[91];
  assign t[123] = t[152] ^ x[94];
  assign t[124] = t[153] ^ x[97];
  assign t[125] = (t[154] & ~t[155]);
  assign t[126] = (t[156] & ~t[157]);
  assign t[127] = (t[158] & ~t[159]);
  assign t[128] = (t[160] & ~t[161]);
  assign t[129] = (t[162] & ~t[163]);
  assign t[12] = t[70] ? x[18] : x[19];
  assign t[130] = (t[164] & ~t[165]);
  assign t[131] = (t[166] & ~t[167]);
  assign t[132] = (t[168] & ~t[169]);
  assign t[133] = (t[170] & ~t[171]);
  assign t[134] = (t[172] & ~t[173]);
  assign t[135] = (t[174] & ~t[175]);
  assign t[136] = (t[176] & ~t[177]);
  assign t[137] = (t[178] & ~t[179]);
  assign t[138] = (t[180] & ~t[181]);
  assign t[139] = (t[182] & ~t[183]);
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = (t[184] & ~t[185]);
  assign t[141] = (t[186] & ~t[187]);
  assign t[142] = (t[188] & ~t[189]);
  assign t[143] = (t[190] & ~t[191]);
  assign t[144] = (t[192] & ~t[193]);
  assign t[145] = (t[194] & ~t[195]);
  assign t[146] = (t[196] & ~t[197]);
  assign t[147] = (t[198] & ~t[199]);
  assign t[148] = (t[200] & ~t[201]);
  assign t[149] = (t[202] & ~t[203]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (t[204] & ~t[205]);
  assign t[151] = (t[206] & ~t[207]);
  assign t[152] = (t[208] & ~t[209]);
  assign t[153] = (t[210] & ~t[211]);
  assign t[154] = t[212] ^ x[2];
  assign t[155] = t[213] ^ x[1];
  assign t[156] = t[214] ^ x[8];
  assign t[157] = t[215] ^ x[7];
  assign t[158] = t[216] ^ x[11];
  assign t[159] = t[217] ^ x[10];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[218] ^ x[14];
  assign t[161] = t[219] ^ x[13];
  assign t[162] = t[220] ^ x[17];
  assign t[163] = t[221] ^ x[16];
  assign t[164] = t[222] ^ x[22];
  assign t[165] = t[223] ^ x[21];
  assign t[166] = t[224] ^ x[27];
  assign t[167] = t[225] ^ x[26];
  assign t[168] = t[226] ^ x[30];
  assign t[169] = t[227] ^ x[29];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[228] ^ x[33];
  assign t[171] = t[229] ^ x[32];
  assign t[172] = t[230] ^ x[36];
  assign t[173] = t[231] ^ x[35];
  assign t[174] = t[232] ^ x[41];
  assign t[175] = t[233] ^ x[40];
  assign t[176] = t[234] ^ x[46];
  assign t[177] = t[235] ^ x[45];
  assign t[178] = t[236] ^ x[49];
  assign t[179] = t[237] ^ x[48];
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = t[238] ^ x[52];
  assign t[181] = t[239] ^ x[51];
  assign t[182] = t[240] ^ x[55];
  assign t[183] = t[241] ^ x[54];
  assign t[184] = t[242] ^ x[58];
  assign t[185] = t[243] ^ x[57];
  assign t[186] = t[244] ^ x[61];
  assign t[187] = t[245] ^ x[60];
  assign t[188] = t[246] ^ x[64];
  assign t[189] = t[247] ^ x[63];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[248] ^ x[67];
  assign t[191] = t[249] ^ x[66];
  assign t[192] = t[250] ^ x[70];
  assign t[193] = t[251] ^ x[69];
  assign t[194] = t[252] ^ x[73];
  assign t[195] = t[253] ^ x[72];
  assign t[196] = t[254] ^ x[76];
  assign t[197] = t[255] ^ x[75];
  assign t[198] = t[256] ^ x[79];
  assign t[199] = t[257] ^ x[78];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[258] ^ x[82];
  assign t[201] = t[259] ^ x[81];
  assign t[202] = t[260] ^ x[85];
  assign t[203] = t[261] ^ x[84];
  assign t[204] = t[262] ^ x[88];
  assign t[205] = t[263] ^ x[87];
  assign t[206] = t[264] ^ x[91];
  assign t[207] = t[265] ^ x[90];
  assign t[208] = t[266] ^ x[94];
  assign t[209] = t[267] ^ x[93];
  assign t[20] = t[29] | t[72];
  assign t[210] = t[268] ^ x[97];
  assign t[211] = t[269] ^ x[96];
  assign t[212] = (x[0]);
  assign t[213] = (x[0]);
  assign t[214] = (x[6]);
  assign t[215] = (x[6]);
  assign t[216] = (x[9]);
  assign t[217] = (x[9]);
  assign t[218] = (x[12]);
  assign t[219] = (x[12]);
  assign t[21] = t[70] ? x[24] : x[23];
  assign t[220] = (x[15]);
  assign t[221] = (x[15]);
  assign t[222] = (x[20]);
  assign t[223] = (x[20]);
  assign t[224] = (x[25]);
  assign t[225] = (x[25]);
  assign t[226] = (x[28]);
  assign t[227] = (x[28]);
  assign t[228] = (x[31]);
  assign t[229] = (x[31]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[34]);
  assign t[231] = (x[34]);
  assign t[232] = (x[39]);
  assign t[233] = (x[39]);
  assign t[234] = (x[44]);
  assign t[235] = (x[44]);
  assign t[236] = (x[47]);
  assign t[237] = (x[47]);
  assign t[238] = (x[50]);
  assign t[239] = (x[50]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[240] = (x[53]);
  assign t[241] = (x[53]);
  assign t[242] = (x[56]);
  assign t[243] = (x[56]);
  assign t[244] = (x[59]);
  assign t[245] = (x[59]);
  assign t[246] = (x[62]);
  assign t[247] = (x[62]);
  assign t[248] = (x[65]);
  assign t[249] = (x[65]);
  assign t[24] = t[34] ^ t[35];
  assign t[250] = (x[68]);
  assign t[251] = (x[68]);
  assign t[252] = (x[71]);
  assign t[253] = (x[71]);
  assign t[254] = (x[74]);
  assign t[255] = (x[74]);
  assign t[256] = (x[77]);
  assign t[257] = (x[77]);
  assign t[258] = (x[80]);
  assign t[259] = (x[80]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[260] = (x[83]);
  assign t[261] = (x[83]);
  assign t[262] = (x[86]);
  assign t[263] = (x[86]);
  assign t[264] = (x[89]);
  assign t[265] = (x[89]);
  assign t[266] = (x[92]);
  assign t[267] = (x[92]);
  assign t[268] = (x[95]);
  assign t[269] = (x[95]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = ~(t[73]);
  assign t[28] = ~(t[74]);
  assign t[29] = ~(t[40] | t[27]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[41] & t[42]);
  assign t[31] = t[43] | t[75];
  assign t[32] = ~(t[44] & t[45]);
  assign t[33] = t[46] | t[76];
  assign t[34] = t[70] ? x[38] : x[37];
  assign t[35] = ~(t[47] & t[48]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = t[51] | t[77];
  assign t[38] = t[52] ? x[43] : x[42];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[78]);
  assign t[41] = ~(t[79]);
  assign t[42] = ~(t[80]);
  assign t[43] = ~(t[55] | t[41]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[56] | t[44]);
  assign t[47] = ~(t[57] & t[58]);
  assign t[48] = t[59] | t[83];
  assign t[49] = ~(t[84]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[85]);
  assign t[51] = ~(t[60] | t[49]);
  assign t[52] = ~(t[61]);
  assign t[53] = ~(t[62] & t[63]);
  assign t[54] = t[64] | t[86];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[89]);
  assign t[58] = ~(t[90]);
  assign t[59] = ~(t[65] | t[57]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[70]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[66] | t[62]);
  assign t[65] = ~(t[94]);
  assign t[66] = ~(t[95]);
  assign t[67] = (t[96]);
  assign t[68] = (t[97]);
  assign t[69] = (t[98]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[68] & t[69]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[70] & t[71]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = t[125] ^ x[2];
  assign t[97] = t[126] ^ x[8];
  assign t[98] = t[127] ^ x[11];
  assign t[99] = t[128] ^ x[14];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [97:0] x;
 output y;

 wire [269:0] t;
  assign t[0] = t[1] ? t[2] : t[67];
  assign t[100] = t[129] ^ x[17];
  assign t[101] = t[130] ^ x[22];
  assign t[102] = t[131] ^ x[27];
  assign t[103] = t[132] ^ x[30];
  assign t[104] = t[133] ^ x[33];
  assign t[105] = t[134] ^ x[36];
  assign t[106] = t[135] ^ x[41];
  assign t[107] = t[136] ^ x[46];
  assign t[108] = t[137] ^ x[49];
  assign t[109] = t[138] ^ x[52];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[55];
  assign t[111] = t[140] ^ x[58];
  assign t[112] = t[141] ^ x[61];
  assign t[113] = t[142] ^ x[64];
  assign t[114] = t[143] ^ x[67];
  assign t[115] = t[144] ^ x[70];
  assign t[116] = t[145] ^ x[73];
  assign t[117] = t[146] ^ x[76];
  assign t[118] = t[147] ^ x[79];
  assign t[119] = t[148] ^ x[82];
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[149] ^ x[85];
  assign t[121] = t[150] ^ x[88];
  assign t[122] = t[151] ^ x[91];
  assign t[123] = t[152] ^ x[94];
  assign t[124] = t[153] ^ x[97];
  assign t[125] = (t[154] & ~t[155]);
  assign t[126] = (t[156] & ~t[157]);
  assign t[127] = (t[158] & ~t[159]);
  assign t[128] = (t[160] & ~t[161]);
  assign t[129] = (t[162] & ~t[163]);
  assign t[12] = t[70] ? x[18] : x[19];
  assign t[130] = (t[164] & ~t[165]);
  assign t[131] = (t[166] & ~t[167]);
  assign t[132] = (t[168] & ~t[169]);
  assign t[133] = (t[170] & ~t[171]);
  assign t[134] = (t[172] & ~t[173]);
  assign t[135] = (t[174] & ~t[175]);
  assign t[136] = (t[176] & ~t[177]);
  assign t[137] = (t[178] & ~t[179]);
  assign t[138] = (t[180] & ~t[181]);
  assign t[139] = (t[182] & ~t[183]);
  assign t[13] = x[4] ? t[16] : t[15];
  assign t[140] = (t[184] & ~t[185]);
  assign t[141] = (t[186] & ~t[187]);
  assign t[142] = (t[188] & ~t[189]);
  assign t[143] = (t[190] & ~t[191]);
  assign t[144] = (t[192] & ~t[193]);
  assign t[145] = (t[194] & ~t[195]);
  assign t[146] = (t[196] & ~t[197]);
  assign t[147] = (t[198] & ~t[199]);
  assign t[148] = (t[200] & ~t[201]);
  assign t[149] = (t[202] & ~t[203]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (t[204] & ~t[205]);
  assign t[151] = (t[206] & ~t[207]);
  assign t[152] = (t[208] & ~t[209]);
  assign t[153] = (t[210] & ~t[211]);
  assign t[154] = t[212] ^ x[2];
  assign t[155] = t[213] ^ x[1];
  assign t[156] = t[214] ^ x[8];
  assign t[157] = t[215] ^ x[7];
  assign t[158] = t[216] ^ x[11];
  assign t[159] = t[217] ^ x[10];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[218] ^ x[14];
  assign t[161] = t[219] ^ x[13];
  assign t[162] = t[220] ^ x[17];
  assign t[163] = t[221] ^ x[16];
  assign t[164] = t[222] ^ x[22];
  assign t[165] = t[223] ^ x[21];
  assign t[166] = t[224] ^ x[27];
  assign t[167] = t[225] ^ x[26];
  assign t[168] = t[226] ^ x[30];
  assign t[169] = t[227] ^ x[29];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[228] ^ x[33];
  assign t[171] = t[229] ^ x[32];
  assign t[172] = t[230] ^ x[36];
  assign t[173] = t[231] ^ x[35];
  assign t[174] = t[232] ^ x[41];
  assign t[175] = t[233] ^ x[40];
  assign t[176] = t[234] ^ x[46];
  assign t[177] = t[235] ^ x[45];
  assign t[178] = t[236] ^ x[49];
  assign t[179] = t[237] ^ x[48];
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = t[238] ^ x[52];
  assign t[181] = t[239] ^ x[51];
  assign t[182] = t[240] ^ x[55];
  assign t[183] = t[241] ^ x[54];
  assign t[184] = t[242] ^ x[58];
  assign t[185] = t[243] ^ x[57];
  assign t[186] = t[244] ^ x[61];
  assign t[187] = t[245] ^ x[60];
  assign t[188] = t[246] ^ x[64];
  assign t[189] = t[247] ^ x[63];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[248] ^ x[67];
  assign t[191] = t[249] ^ x[66];
  assign t[192] = t[250] ^ x[70];
  assign t[193] = t[251] ^ x[69];
  assign t[194] = t[252] ^ x[73];
  assign t[195] = t[253] ^ x[72];
  assign t[196] = t[254] ^ x[76];
  assign t[197] = t[255] ^ x[75];
  assign t[198] = t[256] ^ x[79];
  assign t[199] = t[257] ^ x[78];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[258] ^ x[82];
  assign t[201] = t[259] ^ x[81];
  assign t[202] = t[260] ^ x[85];
  assign t[203] = t[261] ^ x[84];
  assign t[204] = t[262] ^ x[88];
  assign t[205] = t[263] ^ x[87];
  assign t[206] = t[264] ^ x[91];
  assign t[207] = t[265] ^ x[90];
  assign t[208] = t[266] ^ x[94];
  assign t[209] = t[267] ^ x[93];
  assign t[20] = t[29] | t[72];
  assign t[210] = t[268] ^ x[97];
  assign t[211] = t[269] ^ x[96];
  assign t[212] = (x[0]);
  assign t[213] = (x[0]);
  assign t[214] = (x[6]);
  assign t[215] = (x[6]);
  assign t[216] = (x[9]);
  assign t[217] = (x[9]);
  assign t[218] = (x[12]);
  assign t[219] = (x[12]);
  assign t[21] = t[70] ? x[24] : x[23];
  assign t[220] = (x[15]);
  assign t[221] = (x[15]);
  assign t[222] = (x[20]);
  assign t[223] = (x[20]);
  assign t[224] = (x[25]);
  assign t[225] = (x[25]);
  assign t[226] = (x[28]);
  assign t[227] = (x[28]);
  assign t[228] = (x[31]);
  assign t[229] = (x[31]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[34]);
  assign t[231] = (x[34]);
  assign t[232] = (x[39]);
  assign t[233] = (x[39]);
  assign t[234] = (x[44]);
  assign t[235] = (x[44]);
  assign t[236] = (x[47]);
  assign t[237] = (x[47]);
  assign t[238] = (x[50]);
  assign t[239] = (x[50]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[240] = (x[53]);
  assign t[241] = (x[53]);
  assign t[242] = (x[56]);
  assign t[243] = (x[56]);
  assign t[244] = (x[59]);
  assign t[245] = (x[59]);
  assign t[246] = (x[62]);
  assign t[247] = (x[62]);
  assign t[248] = (x[65]);
  assign t[249] = (x[65]);
  assign t[24] = t[34] ^ t[35];
  assign t[250] = (x[68]);
  assign t[251] = (x[68]);
  assign t[252] = (x[71]);
  assign t[253] = (x[71]);
  assign t[254] = (x[74]);
  assign t[255] = (x[74]);
  assign t[256] = (x[77]);
  assign t[257] = (x[77]);
  assign t[258] = (x[80]);
  assign t[259] = (x[80]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[260] = (x[83]);
  assign t[261] = (x[83]);
  assign t[262] = (x[86]);
  assign t[263] = (x[86]);
  assign t[264] = (x[89]);
  assign t[265] = (x[89]);
  assign t[266] = (x[92]);
  assign t[267] = (x[92]);
  assign t[268] = (x[95]);
  assign t[269] = (x[95]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = ~(t[73]);
  assign t[28] = ~(t[74]);
  assign t[29] = ~(t[40] | t[27]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[30] = ~(t[41] & t[42]);
  assign t[31] = t[43] | t[75];
  assign t[32] = ~(t[44] & t[45]);
  assign t[33] = t[46] | t[76];
  assign t[34] = t[70] ? x[38] : x[37];
  assign t[35] = ~(t[47] & t[48]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = t[51] | t[77];
  assign t[38] = t[52] ? x[43] : x[42];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[78]);
  assign t[41] = ~(t[79]);
  assign t[42] = ~(t[80]);
  assign t[43] = ~(t[55] | t[41]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[56] | t[44]);
  assign t[47] = ~(t[57] & t[58]);
  assign t[48] = t[59] | t[83];
  assign t[49] = ~(t[84]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[85]);
  assign t[51] = ~(t[60] | t[49]);
  assign t[52] = ~(t[61]);
  assign t[53] = ~(t[62] & t[63]);
  assign t[54] = t[64] | t[86];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[89]);
  assign t[58] = ~(t[90]);
  assign t[59] = ~(t[65] | t[57]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[70]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[66] | t[62]);
  assign t[65] = ~(t[94]);
  assign t[66] = ~(t[95]);
  assign t[67] = (t[96]);
  assign t[68] = (t[97]);
  assign t[69] = (t[98]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[68] & t[69]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[70] & t[71]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = t[125] ^ x[2];
  assign t[97] = t[126] ^ x[8];
  assign t[98] = t[127] ^ x[11];
  assign t[99] = t[128] ^ x[14];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[224]);
  assign t[101] = ~(t[213] | t[214]);
  assign t[102] = ~(t[138] & t[140]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[141] | t[142]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[227] | t[145]);
  assign t[108] = t[204] ? x[95] : x[94];
  assign t[109] = ~(t[146] & t[147]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[228]);
  assign t[111] = ~(t[229]);
  assign t[112] = ~(t[148] | t[149]);
  assign t[113] = ~(t[150] | t[151]);
  assign t[114] = ~(t[230] | t[152]);
  assign t[115] = t[204] ? x[106] : x[105];
  assign t[116] = ~(t[146] & t[153]);
  assign t[117] = ~(t[122] | t[202]);
  assign t[118] = ~(t[154] & t[155]);
  assign t[119] = ~(t[203] | t[156]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[80] & t[202];
  assign t[121] = ~(t[122] | t[157]);
  assign t[122] = ~(t[204]);
  assign t[123] = t[202] ? t[159] : t[158];
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[161] & t[156]);
  assign t[126] = ~(t[231]);
  assign t[127] = ~(t[218] | t[219]);
  assign t[128] = ~(t[162] & t[163]);
  assign t[129] = ~(t[164] & t[79]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = ~(t[80] | t[165]);
  assign t[131] = ~(t[80] | t[166]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[220] | t[221]);
  assign t[134] = ~(t[130] | t[167]);
  assign t[135] = ~(t[168] | t[169]);
  assign t[136] = ~(t[233]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[49] | t[170]);
  assign t[139] = ~(t[171] | t[172]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = ~(t[167] | t[131]);
  assign t[141] = ~(t[234]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[235]);
  assign t[144] = ~(t[236]);
  assign t[145] = ~(t[173] | t[174]);
  assign t[146] = ~(t[49] | t[175]);
  assign t[147] = ~(t[121] | t[176]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = ~(t[238]);
  assign t[151] = ~(t[239]);
  assign t[152] = ~(t[177] | t[178]);
  assign t[153] = ~(t[179] | t[131]);
  assign t[154] = ~(t[205] & t[180]);
  assign t[155] = ~(x[4] & t[119]);
  assign t[156] = ~(t[205]);
  assign t[157] = t[202] ? t[158] : t[159];
  assign t[158] = ~(t[180] & t[156]);
  assign t[159] = ~(x[4] & t[181]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = x[4] & t[203];
  assign t[161] = ~(x[4] | t[203]);
  assign t[162] = ~(t[171] | t[182]);
  assign t[163] = ~(t[122] & t[183]);
  assign t[164] = ~(t[184] & t[185]);
  assign t[165] = t[202] ? t[124] : t[125];
  assign t[166] = t[202] ? t[187] : t[186];
  assign t[167] = ~(t[80] | t[188]);
  assign t[168] = t[172] | t[189];
  assign t[169] = ~(t[190] & t[79]);
  assign t[16] = x[4] ? t[25] : t[24];
  assign t[170] = ~(t[80] | t[191]);
  assign t[171] = ~(t[122] | t[192]);
  assign t[172] = ~(t[193] & t[77]);
  assign t[173] = ~(t[240]);
  assign t[174] = ~(t[235] | t[236]);
  assign t[175] = ~(t[134] & t[164]);
  assign t[176] = t[170] | t[194];
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[238] | t[239]);
  assign t[179] = ~(t[80] | t[195]);
  assign t[17] = ~(t[26] ^ t[27]);
  assign t[180] = ~(x[4] | t[196]);
  assign t[181] = ~(t[203] | t[205]);
  assign t[182] = ~(t[80] | t[197]);
  assign t[183] = ~(t[159] & t[154]);
  assign t[184] = t[205] & t[117];
  assign t[185] = t[161] | t[160];
  assign t[186] = ~(t[161] & t[205]);
  assign t[187] = ~(t[160] & t[156]);
  assign t[188] = t[202] ? t[159] : t[154];
  assign t[189] = ~(t[80] | t[198]);
  assign t[18] = t[28] ? x[18] : x[19];
  assign t[190] = ~(t[194] | t[179]);
  assign t[191] = t[202] ? t[186] : t[187];
  assign t[192] = t[202] ? t[125] : t[187];
  assign t[193] = ~(t[199] | t[121]);
  assign t[194] = ~(t[76]);
  assign t[195] = t[202] ? t[155] : t[158];
  assign t[196] = ~(t[203]);
  assign t[197] = t[202] ? t[158] : t[155];
  assign t[198] = t[202] ? t[154] : t[159];
  assign t[199] = ~(t[122] | t[200]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[202] ? t[187] : t[125];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = ~(t[31] | t[32]);
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[33] ^ t[34]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = x[4] ? t[36] : t[35];
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = x[4] ? t[38] : t[37];
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[8];
  assign t[244] = t[285] ^ x[11];
  assign t[245] = t[286] ^ x[14];
  assign t[246] = t[287] ^ x[17];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = ~(t[39] | t[40]);
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[34];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = ~(t[24] ^ t[41]);
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[68];
  assign t[262] = t[303] ^ x[71];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[79];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[98];
  assign t[26] = x[4] ? t[43] : t[42];
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = ~(t[46]);
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[8];
  assign t[327] = t[409] ^ x[7];
  assign t[328] = t[410] ^ x[11];
  assign t[329] = t[411] ^ x[10];
  assign t[32] = ~(t[206] | t[52]);
  assign t[330] = t[412] ^ x[14];
  assign t[331] = t[413] ^ x[13];
  assign t[332] = t[414] ^ x[17];
  assign t[333] = t[415] ^ x[16];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[34];
  assign t[343] = t[425] ^ x[33];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[68];
  assign t[363] = t[445] ^ x[67];
  assign t[364] = t[446] ^ x[71];
  assign t[365] = t[447] ^ x[70];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[79];
  assign t[369] = t[451] ^ x[78];
  assign t[36] = ~(t[44] ^ t[59]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[98];
  assign t[379] = t[461] ^ x[97];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[35] ^ t[62]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[6]);
  assign t[409] = (x[6]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[9]);
  assign t[411] = (x[9]);
  assign t[412] = (x[12]);
  assign t[413] = (x[12]);
  assign t[414] = (x[15]);
  assign t[415] = (x[15]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[66] ^ t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[32]);
  assign t[425] = (x[32]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[66]);
  assign t[445] = (x[66]);
  assign t[446] = (x[69]);
  assign t[447] = (x[69]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[77]);
  assign t[451] = (x[77]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = (x[96]);
  assign t[461] = (x[96]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[204]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[78] & t[79]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[208]);
  assign t[51] = ~(t[209]);
  assign t[52] = ~(t[82] | t[83]);
  assign t[53] = ~(t[84] | t[85]);
  assign t[54] = ~(t[210] | t[86]);
  assign t[55] = t[87] ? x[36] : x[35];
  assign t[56] = ~(t[88] & t[89]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[58] = ~(t[211] | t[92]);
  assign t[59] = ~(t[93] ^ t[94]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[212] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[213]);
  assign t[64] = ~(t[214]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = t[204] ? x[50] : x[49];
  assign t[67] = t[47] | t[102];
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[215] | t[105]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[108] ^ t[109]);
  assign t[72] = ~(t[110] | t[111]);
  assign t[73] = ~(t[216] | t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117] & t[118]);
  assign t[77] = ~(t[119] & t[120]);
  assign t[78] = ~(t[121]);
  assign t[79] = t[122] | t[123];
  assign t[7] = ~(t[202] & t[203]);
  assign t[80] = ~(t[122]);
  assign t[81] = t[202] ? t[125] : t[124];
  assign t[82] = ~(t[217]);
  assign t[83] = ~(t[208] | t[209]);
  assign t[84] = ~(t[218]);
  assign t[85] = ~(t[219]);
  assign t[86] = ~(t[126] | t[127]);
  assign t[87] = ~(t[46]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = ~(t[204] & t[205]);
  assign t[90] = ~(t[220]);
  assign t[91] = ~(t[221]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = t[87] ? x[73] : x[72];
  assign t[94] = ~(t[134] & t[135]);
  assign t[95] = ~(t[222]);
  assign t[96] = ~(t[223]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[87] ? x[81] : x[80];
  assign t[99] = ~(t[138] & t[139]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[224]);
  assign t[101] = ~(t[213] | t[214]);
  assign t[102] = ~(t[138] & t[140]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[141] | t[142]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[227] | t[145]);
  assign t[108] = t[204] ? x[95] : x[94];
  assign t[109] = ~(t[146] & t[147]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[228]);
  assign t[111] = ~(t[229]);
  assign t[112] = ~(t[148] | t[149]);
  assign t[113] = ~(t[150] | t[151]);
  assign t[114] = ~(t[230] | t[152]);
  assign t[115] = t[204] ? x[106] : x[105];
  assign t[116] = ~(t[146] & t[153]);
  assign t[117] = ~(t[122] | t[202]);
  assign t[118] = ~(t[154] & t[155]);
  assign t[119] = ~(t[203] | t[156]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = t[80] & t[202];
  assign t[121] = ~(t[122] | t[157]);
  assign t[122] = ~(t[204]);
  assign t[123] = t[202] ? t[159] : t[158];
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[161] & t[156]);
  assign t[126] = ~(t[231]);
  assign t[127] = ~(t[218] | t[219]);
  assign t[128] = ~(t[162] & t[163]);
  assign t[129] = ~(t[164] & t[79]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = ~(t[80] | t[165]);
  assign t[131] = ~(t[80] | t[166]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[220] | t[221]);
  assign t[134] = ~(t[130] | t[167]);
  assign t[135] = ~(t[168] | t[169]);
  assign t[136] = ~(t[233]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[49] | t[170]);
  assign t[139] = ~(t[171] | t[172]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = ~(t[167] | t[131]);
  assign t[141] = ~(t[234]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[235]);
  assign t[144] = ~(t[236]);
  assign t[145] = ~(t[173] | t[174]);
  assign t[146] = ~(t[49] | t[175]);
  assign t[147] = ~(t[121] | t[176]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = ~(t[238]);
  assign t[151] = ~(t[239]);
  assign t[152] = ~(t[177] | t[178]);
  assign t[153] = ~(t[179] | t[131]);
  assign t[154] = ~(t[205] & t[180]);
  assign t[155] = ~(x[4] & t[119]);
  assign t[156] = ~(t[205]);
  assign t[157] = t[202] ? t[158] : t[159];
  assign t[158] = ~(t[180] & t[156]);
  assign t[159] = ~(x[4] & t[181]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = x[4] & t[203];
  assign t[161] = ~(x[4] | t[203]);
  assign t[162] = ~(t[171] | t[182]);
  assign t[163] = ~(t[122] & t[183]);
  assign t[164] = ~(t[184] & t[185]);
  assign t[165] = t[202] ? t[124] : t[125];
  assign t[166] = t[202] ? t[187] : t[186];
  assign t[167] = ~(t[80] | t[188]);
  assign t[168] = t[172] | t[189];
  assign t[169] = ~(t[190] & t[79]);
  assign t[16] = x[4] ? t[25] : t[24];
  assign t[170] = ~(t[80] | t[191]);
  assign t[171] = ~(t[122] | t[192]);
  assign t[172] = ~(t[193] & t[77]);
  assign t[173] = ~(t[240]);
  assign t[174] = ~(t[235] | t[236]);
  assign t[175] = ~(t[134] & t[164]);
  assign t[176] = t[170] | t[194];
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[238] | t[239]);
  assign t[179] = ~(t[80] | t[195]);
  assign t[17] = ~(t[26] ^ t[27]);
  assign t[180] = ~(x[4] | t[196]);
  assign t[181] = ~(t[203] | t[205]);
  assign t[182] = ~(t[80] | t[197]);
  assign t[183] = ~(t[159] & t[154]);
  assign t[184] = t[205] & t[117];
  assign t[185] = t[161] | t[160];
  assign t[186] = ~(t[161] & t[205]);
  assign t[187] = ~(t[160] & t[156]);
  assign t[188] = t[202] ? t[159] : t[154];
  assign t[189] = ~(t[80] | t[198]);
  assign t[18] = t[28] ? x[18] : x[19];
  assign t[190] = ~(t[194] | t[179]);
  assign t[191] = t[202] ? t[186] : t[187];
  assign t[192] = t[202] ? t[125] : t[187];
  assign t[193] = ~(t[199] | t[121]);
  assign t[194] = ~(t[76]);
  assign t[195] = t[202] ? t[155] : t[158];
  assign t[196] = ~(t[203]);
  assign t[197] = t[202] ? t[158] : t[155];
  assign t[198] = t[202] ? t[154] : t[159];
  assign t[199] = ~(t[122] | t[200]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[202] ? t[187] : t[125];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = ~(t[31] | t[32]);
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[33] ^ t[34]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = x[4] ? t[36] : t[35];
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = x[4] ? t[38] : t[37];
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[8];
  assign t[244] = t[285] ^ x[11];
  assign t[245] = t[286] ^ x[14];
  assign t[246] = t[287] ^ x[17];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = ~(t[39] | t[40]);
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[34];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = ~(t[24] ^ t[41]);
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[68];
  assign t[262] = t[303] ^ x[71];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[79];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[98];
  assign t[26] = x[4] ? t[43] : t[42];
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = ~(t[46]);
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[8];
  assign t[327] = t[409] ^ x[7];
  assign t[328] = t[410] ^ x[11];
  assign t[329] = t[411] ^ x[10];
  assign t[32] = ~(t[206] | t[52]);
  assign t[330] = t[412] ^ x[14];
  assign t[331] = t[413] ^ x[13];
  assign t[332] = t[414] ^ x[17];
  assign t[333] = t[415] ^ x[16];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[34];
  assign t[343] = t[425] ^ x[33];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[68];
  assign t[363] = t[445] ^ x[67];
  assign t[364] = t[446] ^ x[71];
  assign t[365] = t[447] ^ x[70];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[79];
  assign t[369] = t[451] ^ x[78];
  assign t[36] = ~(t[44] ^ t[59]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[98];
  assign t[379] = t[461] ^ x[97];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[35] ^ t[62]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[6]);
  assign t[409] = (x[6]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[9]);
  assign t[411] = (x[9]);
  assign t[412] = (x[12]);
  assign t[413] = (x[12]);
  assign t[414] = (x[15]);
  assign t[415] = (x[15]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[66] ^ t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[32]);
  assign t[425] = (x[32]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[66]);
  assign t[445] = (x[66]);
  assign t[446] = (x[69]);
  assign t[447] = (x[69]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[77]);
  assign t[451] = (x[77]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = (x[96]);
  assign t[461] = (x[96]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[204]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[78] & t[79]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[208]);
  assign t[51] = ~(t[209]);
  assign t[52] = ~(t[82] | t[83]);
  assign t[53] = ~(t[84] | t[85]);
  assign t[54] = ~(t[210] | t[86]);
  assign t[55] = t[87] ? x[36] : x[35];
  assign t[56] = ~(t[88] & t[89]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[58] = ~(t[211] | t[92]);
  assign t[59] = ~(t[93] ^ t[94]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[212] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[213]);
  assign t[64] = ~(t[214]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = t[204] ? x[50] : x[49];
  assign t[67] = t[47] | t[102];
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[215] | t[105]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[108] ^ t[109]);
  assign t[72] = ~(t[110] | t[111]);
  assign t[73] = ~(t[216] | t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117] & t[118]);
  assign t[77] = ~(t[119] & t[120]);
  assign t[78] = ~(t[121]);
  assign t[79] = t[122] | t[123];
  assign t[7] = ~(t[202] & t[203]);
  assign t[80] = ~(t[122]);
  assign t[81] = t[202] ? t[125] : t[124];
  assign t[82] = ~(t[217]);
  assign t[83] = ~(t[208] | t[209]);
  assign t[84] = ~(t[218]);
  assign t[85] = ~(t[219]);
  assign t[86] = ~(t[126] | t[127]);
  assign t[87] = ~(t[46]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = ~(t[204] & t[205]);
  assign t[90] = ~(t[220]);
  assign t[91] = ~(t[221]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = t[87] ? x[73] : x[72];
  assign t[94] = ~(t[134] & t[135]);
  assign t[95] = ~(t[222]);
  assign t[96] = ~(t[223]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[87] ? x[81] : x[80];
  assign t[99] = ~(t[138] & t[139]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind166(x, y);
 input [112:0] x;
 output y;

 wire [315:0] t;
  assign t[0] = t[1] ? t[2] : t[92];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = t[156] ^ x[2];
  assign t[125] = t[157] ^ x[8];
  assign t[126] = t[158] ^ x[11];
  assign t[127] = t[159] ^ x[14];
  assign t[128] = t[160] ^ x[17];
  assign t[129] = t[161] ^ x[22];
  assign t[12] = t[95] ? x[18] : x[19];
  assign t[130] = t[162] ^ x[25];
  assign t[131] = t[163] ^ x[30];
  assign t[132] = t[164] ^ x[33];
  assign t[133] = t[165] ^ x[38];
  assign t[134] = t[166] ^ x[41];
  assign t[135] = t[167] ^ x[44];
  assign t[136] = t[168] ^ x[47];
  assign t[137] = t[169] ^ x[50];
  assign t[138] = t[170] ^ x[55];
  assign t[139] = t[171] ^ x[58];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[63];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[69];
  assign t[143] = t[175] ^ x[74];
  assign t[144] = t[176] ^ x[77];
  assign t[145] = t[177] ^ x[82];
  assign t[146] = t[178] ^ x[85];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = t[180] ^ x[91];
  assign t[149] = t[181] ^ x[94];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[97];
  assign t[151] = t[183] ^ x[100];
  assign t[152] = t[184] ^ x[103];
  assign t[153] = t[185] ^ x[106];
  assign t[154] = t[186] ^ x[109];
  assign t[155] = t[187] ^ x[112];
  assign t[156] = (t[188] & ~t[189]);
  assign t[157] = (t[190] & ~t[191]);
  assign t[158] = (t[192] & ~t[193]);
  assign t[159] = (t[194] & ~t[195]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (t[196] & ~t[197]);
  assign t[161] = (t[198] & ~t[199]);
  assign t[162] = (t[200] & ~t[201]);
  assign t[163] = (t[202] & ~t[203]);
  assign t[164] = (t[204] & ~t[205]);
  assign t[165] = (t[206] & ~t[207]);
  assign t[166] = (t[208] & ~t[209]);
  assign t[167] = (t[210] & ~t[211]);
  assign t[168] = (t[212] & ~t[213]);
  assign t[169] = (t[214] & ~t[215]);
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = (t[216] & ~t[217]);
  assign t[171] = (t[218] & ~t[219]);
  assign t[172] = (t[220] & ~t[221]);
  assign t[173] = (t[222] & ~t[223]);
  assign t[174] = (t[224] & ~t[225]);
  assign t[175] = (t[226] & ~t[227]);
  assign t[176] = (t[228] & ~t[229]);
  assign t[177] = (t[230] & ~t[231]);
  assign t[178] = (t[232] & ~t[233]);
  assign t[179] = (t[234] & ~t[235]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (t[236] & ~t[237]);
  assign t[181] = (t[238] & ~t[239]);
  assign t[182] = (t[240] & ~t[241]);
  assign t[183] = (t[242] & ~t[243]);
  assign t[184] = (t[244] & ~t[245]);
  assign t[185] = (t[246] & ~t[247]);
  assign t[186] = (t[248] & ~t[249]);
  assign t[187] = (t[250] & ~t[251]);
  assign t[188] = t[252] ^ x[2];
  assign t[189] = t[253] ^ x[1];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[254] ^ x[8];
  assign t[191] = t[255] ^ x[7];
  assign t[192] = t[256] ^ x[11];
  assign t[193] = t[257] ^ x[10];
  assign t[194] = t[258] ^ x[14];
  assign t[195] = t[259] ^ x[13];
  assign t[196] = t[260] ^ x[17];
  assign t[197] = t[261] ^ x[16];
  assign t[198] = t[262] ^ x[22];
  assign t[199] = t[263] ^ x[21];
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[264] ^ x[25];
  assign t[201] = t[265] ^ x[24];
  assign t[202] = t[266] ^ x[30];
  assign t[203] = t[267] ^ x[29];
  assign t[204] = t[268] ^ x[33];
  assign t[205] = t[269] ^ x[32];
  assign t[206] = t[270] ^ x[38];
  assign t[207] = t[271] ^ x[37];
  assign t[208] = t[272] ^ x[41];
  assign t[209] = t[273] ^ x[40];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = t[274] ^ x[44];
  assign t[211] = t[275] ^ x[43];
  assign t[212] = t[276] ^ x[47];
  assign t[213] = t[277] ^ x[46];
  assign t[214] = t[278] ^ x[50];
  assign t[215] = t[279] ^ x[49];
  assign t[216] = t[280] ^ x[55];
  assign t[217] = t[281] ^ x[54];
  assign t[218] = t[282] ^ x[58];
  assign t[219] = t[283] ^ x[57];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[284] ^ x[63];
  assign t[221] = t[285] ^ x[62];
  assign t[222] = t[286] ^ x[66];
  assign t[223] = t[287] ^ x[65];
  assign t[224] = t[288] ^ x[69];
  assign t[225] = t[289] ^ x[68];
  assign t[226] = t[290] ^ x[74];
  assign t[227] = t[291] ^ x[73];
  assign t[228] = t[292] ^ x[77];
  assign t[229] = t[293] ^ x[76];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[294] ^ x[82];
  assign t[231] = t[295] ^ x[81];
  assign t[232] = t[296] ^ x[85];
  assign t[233] = t[297] ^ x[84];
  assign t[234] = t[298] ^ x[88];
  assign t[235] = t[299] ^ x[87];
  assign t[236] = t[300] ^ x[91];
  assign t[237] = t[301] ^ x[90];
  assign t[238] = t[302] ^ x[94];
  assign t[239] = t[303] ^ x[93];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[304] ^ x[97];
  assign t[241] = t[305] ^ x[96];
  assign t[242] = t[306] ^ x[100];
  assign t[243] = t[307] ^ x[99];
  assign t[244] = t[308] ^ x[103];
  assign t[245] = t[309] ^ x[102];
  assign t[246] = t[310] ^ x[106];
  assign t[247] = t[311] ^ x[105];
  assign t[248] = t[312] ^ x[109];
  assign t[249] = t[313] ^ x[108];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[314] ^ x[112];
  assign t[251] = t[315] ^ x[111];
  assign t[252] = (x[0]);
  assign t[253] = (x[0]);
  assign t[254] = (x[6]);
  assign t[255] = (x[6]);
  assign t[256] = (x[9]);
  assign t[257] = (x[9]);
  assign t[258] = (x[12]);
  assign t[259] = (x[12]);
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = (x[15]);
  assign t[261] = (x[15]);
  assign t[262] = (x[20]);
  assign t[263] = (x[20]);
  assign t[264] = (x[23]);
  assign t[265] = (x[23]);
  assign t[266] = (x[28]);
  assign t[267] = (x[28]);
  assign t[268] = (x[31]);
  assign t[269] = (x[31]);
  assign t[26] = ~(t[97] & t[41]);
  assign t[270] = (x[36]);
  assign t[271] = (x[36]);
  assign t[272] = (x[39]);
  assign t[273] = (x[39]);
  assign t[274] = (x[42]);
  assign t[275] = (x[42]);
  assign t[276] = (x[45]);
  assign t[277] = (x[45]);
  assign t[278] = (x[48]);
  assign t[279] = (x[48]);
  assign t[27] = ~(t[98] & t[42]);
  assign t[280] = (x[53]);
  assign t[281] = (x[53]);
  assign t[282] = (x[56]);
  assign t[283] = (x[56]);
  assign t[284] = (x[61]);
  assign t[285] = (x[61]);
  assign t[286] = (x[64]);
  assign t[287] = (x[64]);
  assign t[288] = (x[67]);
  assign t[289] = (x[67]);
  assign t[28] = t[43] ? x[27] : x[26];
  assign t[290] = (x[72]);
  assign t[291] = (x[72]);
  assign t[292] = (x[75]);
  assign t[293] = (x[75]);
  assign t[294] = (x[80]);
  assign t[295] = (x[80]);
  assign t[296] = (x[83]);
  assign t[297] = (x[83]);
  assign t[298] = (x[86]);
  assign t[299] = (x[86]);
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[89]);
  assign t[301] = (x[89]);
  assign t[302] = (x[92]);
  assign t[303] = (x[92]);
  assign t[304] = (x[95]);
  assign t[305] = (x[95]);
  assign t[306] = (x[98]);
  assign t[307] = (x[98]);
  assign t[308] = (x[101]);
  assign t[309] = (x[101]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[104]);
  assign t[311] = (x[104]);
  assign t[312] = (x[107]);
  assign t[313] = (x[107]);
  assign t[314] = (x[110]);
  assign t[315] = (x[110]);
  assign t[31] = t[48] ^ t[32];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[37];
  assign t[34] = ~(t[99] & t[52]);
  assign t[35] = ~(t[100] & t[53]);
  assign t[36] = t[95] ? x[35] : x[34];
  assign t[37] = ~(t[54] & t[55]);
  assign t[38] = t[56] ^ t[57];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[101]);
  assign t[42] = ~(t[101] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[102] & t[64]);
  assign t[45] = ~(t[103] & t[65]);
  assign t[46] = ~(t[104] & t[66]);
  assign t[47] = ~(t[105] & t[67]);
  assign t[48] = t[68] ? x[52] : x[51];
  assign t[49] = ~(t[106] & t[69]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[107] & t[70]);
  assign t[51] = t[71] ? x[60] : x[59];
  assign t[52] = ~(t[108]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = ~(t[110] & t[74]);
  assign t[56] = t[95] ? x[71] : x[70];
  assign t[57] = ~(t[75] & t[76]);
  assign t[58] = ~(t[111] & t[77]);
  assign t[59] = ~(t[112] & t[78]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[43] ? x[79] : x[78];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[97]);
  assign t[63] = ~(t[95]);
  assign t[64] = ~(t[113]);
  assign t[65] = ~(t[113] & t[81]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[63]);
  assign t[69] = ~(t[115]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[63]);
  assign t[72] = ~(t[99]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[93] & t[94]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[102]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[106]);
  assign t[84] = ~(t[109]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[122] & t[90]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[123]);
  assign t[89] = ~(t[123] & t[91]);
  assign t[8] = ~(t[95] & t[96]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[120]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [112:0] x;
 output y;

 wire [315:0] t;
  assign t[0] = t[1] ? t[2] : t[92];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = t[156] ^ x[2];
  assign t[125] = t[157] ^ x[8];
  assign t[126] = t[158] ^ x[11];
  assign t[127] = t[159] ^ x[14];
  assign t[128] = t[160] ^ x[17];
  assign t[129] = t[161] ^ x[22];
  assign t[12] = t[95] ? x[18] : x[19];
  assign t[130] = t[162] ^ x[25];
  assign t[131] = t[163] ^ x[30];
  assign t[132] = t[164] ^ x[33];
  assign t[133] = t[165] ^ x[38];
  assign t[134] = t[166] ^ x[41];
  assign t[135] = t[167] ^ x[44];
  assign t[136] = t[168] ^ x[47];
  assign t[137] = t[169] ^ x[50];
  assign t[138] = t[170] ^ x[55];
  assign t[139] = t[171] ^ x[58];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[63];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[69];
  assign t[143] = t[175] ^ x[74];
  assign t[144] = t[176] ^ x[77];
  assign t[145] = t[177] ^ x[82];
  assign t[146] = t[178] ^ x[85];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = t[180] ^ x[91];
  assign t[149] = t[181] ^ x[94];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[97];
  assign t[151] = t[183] ^ x[100];
  assign t[152] = t[184] ^ x[103];
  assign t[153] = t[185] ^ x[106];
  assign t[154] = t[186] ^ x[109];
  assign t[155] = t[187] ^ x[112];
  assign t[156] = (t[188] & ~t[189]);
  assign t[157] = (t[190] & ~t[191]);
  assign t[158] = (t[192] & ~t[193]);
  assign t[159] = (t[194] & ~t[195]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (t[196] & ~t[197]);
  assign t[161] = (t[198] & ~t[199]);
  assign t[162] = (t[200] & ~t[201]);
  assign t[163] = (t[202] & ~t[203]);
  assign t[164] = (t[204] & ~t[205]);
  assign t[165] = (t[206] & ~t[207]);
  assign t[166] = (t[208] & ~t[209]);
  assign t[167] = (t[210] & ~t[211]);
  assign t[168] = (t[212] & ~t[213]);
  assign t[169] = (t[214] & ~t[215]);
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = (t[216] & ~t[217]);
  assign t[171] = (t[218] & ~t[219]);
  assign t[172] = (t[220] & ~t[221]);
  assign t[173] = (t[222] & ~t[223]);
  assign t[174] = (t[224] & ~t[225]);
  assign t[175] = (t[226] & ~t[227]);
  assign t[176] = (t[228] & ~t[229]);
  assign t[177] = (t[230] & ~t[231]);
  assign t[178] = (t[232] & ~t[233]);
  assign t[179] = (t[234] & ~t[235]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (t[236] & ~t[237]);
  assign t[181] = (t[238] & ~t[239]);
  assign t[182] = (t[240] & ~t[241]);
  assign t[183] = (t[242] & ~t[243]);
  assign t[184] = (t[244] & ~t[245]);
  assign t[185] = (t[246] & ~t[247]);
  assign t[186] = (t[248] & ~t[249]);
  assign t[187] = (t[250] & ~t[251]);
  assign t[188] = t[252] ^ x[2];
  assign t[189] = t[253] ^ x[1];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[254] ^ x[8];
  assign t[191] = t[255] ^ x[7];
  assign t[192] = t[256] ^ x[11];
  assign t[193] = t[257] ^ x[10];
  assign t[194] = t[258] ^ x[14];
  assign t[195] = t[259] ^ x[13];
  assign t[196] = t[260] ^ x[17];
  assign t[197] = t[261] ^ x[16];
  assign t[198] = t[262] ^ x[22];
  assign t[199] = t[263] ^ x[21];
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[264] ^ x[25];
  assign t[201] = t[265] ^ x[24];
  assign t[202] = t[266] ^ x[30];
  assign t[203] = t[267] ^ x[29];
  assign t[204] = t[268] ^ x[33];
  assign t[205] = t[269] ^ x[32];
  assign t[206] = t[270] ^ x[38];
  assign t[207] = t[271] ^ x[37];
  assign t[208] = t[272] ^ x[41];
  assign t[209] = t[273] ^ x[40];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = t[274] ^ x[44];
  assign t[211] = t[275] ^ x[43];
  assign t[212] = t[276] ^ x[47];
  assign t[213] = t[277] ^ x[46];
  assign t[214] = t[278] ^ x[50];
  assign t[215] = t[279] ^ x[49];
  assign t[216] = t[280] ^ x[55];
  assign t[217] = t[281] ^ x[54];
  assign t[218] = t[282] ^ x[58];
  assign t[219] = t[283] ^ x[57];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[284] ^ x[63];
  assign t[221] = t[285] ^ x[62];
  assign t[222] = t[286] ^ x[66];
  assign t[223] = t[287] ^ x[65];
  assign t[224] = t[288] ^ x[69];
  assign t[225] = t[289] ^ x[68];
  assign t[226] = t[290] ^ x[74];
  assign t[227] = t[291] ^ x[73];
  assign t[228] = t[292] ^ x[77];
  assign t[229] = t[293] ^ x[76];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[294] ^ x[82];
  assign t[231] = t[295] ^ x[81];
  assign t[232] = t[296] ^ x[85];
  assign t[233] = t[297] ^ x[84];
  assign t[234] = t[298] ^ x[88];
  assign t[235] = t[299] ^ x[87];
  assign t[236] = t[300] ^ x[91];
  assign t[237] = t[301] ^ x[90];
  assign t[238] = t[302] ^ x[94];
  assign t[239] = t[303] ^ x[93];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[304] ^ x[97];
  assign t[241] = t[305] ^ x[96];
  assign t[242] = t[306] ^ x[100];
  assign t[243] = t[307] ^ x[99];
  assign t[244] = t[308] ^ x[103];
  assign t[245] = t[309] ^ x[102];
  assign t[246] = t[310] ^ x[106];
  assign t[247] = t[311] ^ x[105];
  assign t[248] = t[312] ^ x[109];
  assign t[249] = t[313] ^ x[108];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[314] ^ x[112];
  assign t[251] = t[315] ^ x[111];
  assign t[252] = (x[0]);
  assign t[253] = (x[0]);
  assign t[254] = (x[6]);
  assign t[255] = (x[6]);
  assign t[256] = (x[9]);
  assign t[257] = (x[9]);
  assign t[258] = (x[12]);
  assign t[259] = (x[12]);
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = (x[15]);
  assign t[261] = (x[15]);
  assign t[262] = (x[20]);
  assign t[263] = (x[20]);
  assign t[264] = (x[23]);
  assign t[265] = (x[23]);
  assign t[266] = (x[28]);
  assign t[267] = (x[28]);
  assign t[268] = (x[31]);
  assign t[269] = (x[31]);
  assign t[26] = ~(t[97] & t[41]);
  assign t[270] = (x[36]);
  assign t[271] = (x[36]);
  assign t[272] = (x[39]);
  assign t[273] = (x[39]);
  assign t[274] = (x[42]);
  assign t[275] = (x[42]);
  assign t[276] = (x[45]);
  assign t[277] = (x[45]);
  assign t[278] = (x[48]);
  assign t[279] = (x[48]);
  assign t[27] = ~(t[98] & t[42]);
  assign t[280] = (x[53]);
  assign t[281] = (x[53]);
  assign t[282] = (x[56]);
  assign t[283] = (x[56]);
  assign t[284] = (x[61]);
  assign t[285] = (x[61]);
  assign t[286] = (x[64]);
  assign t[287] = (x[64]);
  assign t[288] = (x[67]);
  assign t[289] = (x[67]);
  assign t[28] = t[43] ? x[27] : x[26];
  assign t[290] = (x[72]);
  assign t[291] = (x[72]);
  assign t[292] = (x[75]);
  assign t[293] = (x[75]);
  assign t[294] = (x[80]);
  assign t[295] = (x[80]);
  assign t[296] = (x[83]);
  assign t[297] = (x[83]);
  assign t[298] = (x[86]);
  assign t[299] = (x[86]);
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[89]);
  assign t[301] = (x[89]);
  assign t[302] = (x[92]);
  assign t[303] = (x[92]);
  assign t[304] = (x[95]);
  assign t[305] = (x[95]);
  assign t[306] = (x[98]);
  assign t[307] = (x[98]);
  assign t[308] = (x[101]);
  assign t[309] = (x[101]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[104]);
  assign t[311] = (x[104]);
  assign t[312] = (x[107]);
  assign t[313] = (x[107]);
  assign t[314] = (x[110]);
  assign t[315] = (x[110]);
  assign t[31] = t[48] ^ t[32];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[37];
  assign t[34] = ~(t[99] & t[52]);
  assign t[35] = ~(t[100] & t[53]);
  assign t[36] = t[95] ? x[35] : x[34];
  assign t[37] = ~(t[54] & t[55]);
  assign t[38] = t[56] ^ t[57];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[101]);
  assign t[42] = ~(t[101] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[102] & t[64]);
  assign t[45] = ~(t[103] & t[65]);
  assign t[46] = ~(t[104] & t[66]);
  assign t[47] = ~(t[105] & t[67]);
  assign t[48] = t[68] ? x[52] : x[51];
  assign t[49] = ~(t[106] & t[69]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[107] & t[70]);
  assign t[51] = t[71] ? x[60] : x[59];
  assign t[52] = ~(t[108]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = ~(t[110] & t[74]);
  assign t[56] = t[95] ? x[71] : x[70];
  assign t[57] = ~(t[75] & t[76]);
  assign t[58] = ~(t[111] & t[77]);
  assign t[59] = ~(t[112] & t[78]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[43] ? x[79] : x[78];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[97]);
  assign t[63] = ~(t[95]);
  assign t[64] = ~(t[113]);
  assign t[65] = ~(t[113] & t[81]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[63]);
  assign t[69] = ~(t[115]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[63]);
  assign t[72] = ~(t[99]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[93] & t[94]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[102]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[106]);
  assign t[84] = ~(t[109]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[122] & t[90]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[123]);
  assign t[89] = ~(t[123] & t[91]);
  assign t[8] = ~(t[95] & t[96]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[120]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [139:0] x;
 output y;

 wire [394:0] t;
  assign t[0] = t[1] ? t[2] : t[108];
  assign t[100] = ~(t[144]);
  assign t[101] = ~(t[145]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[106] & t[107]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[147]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[111] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = t[190] ^ x[2];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[8];
  assign t[151] = t[192] ^ x[11];
  assign t[152] = t[193] ^ x[14];
  assign t[153] = t[194] ^ x[17];
  assign t[154] = t[195] ^ x[22];
  assign t[155] = t[196] ^ x[27];
  assign t[156] = t[197] ^ x[32];
  assign t[157] = t[198] ^ x[35];
  assign t[158] = t[199] ^ x[38];
  assign t[159] = t[200] ^ x[41];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[46];
  assign t[161] = t[202] ^ x[51];
  assign t[162] = t[203] ^ x[54];
  assign t[163] = t[204] ^ x[57];
  assign t[164] = t[205] ^ x[62];
  assign t[165] = t[206] ^ x[67];
  assign t[166] = t[207] ^ x[70];
  assign t[167] = t[208] ^ x[73];
  assign t[168] = t[209] ^ x[76];
  assign t[169] = t[210] ^ x[79];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[82];
  assign t[171] = t[212] ^ x[85];
  assign t[172] = t[213] ^ x[88];
  assign t[173] = t[214] ^ x[91];
  assign t[174] = t[215] ^ x[94];
  assign t[175] = t[216] ^ x[97];
  assign t[176] = t[217] ^ x[100];
  assign t[177] = t[218] ^ x[103];
  assign t[178] = t[219] ^ x[106];
  assign t[179] = t[220] ^ x[109];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[112];
  assign t[181] = t[222] ^ x[115];
  assign t[182] = t[223] ^ x[118];
  assign t[183] = t[224] ^ x[121];
  assign t[184] = t[225] ^ x[124];
  assign t[185] = t[226] ^ x[127];
  assign t[186] = t[227] ^ x[130];
  assign t[187] = t[228] ^ x[133];
  assign t[188] = t[229] ^ x[136];
  assign t[189] = t[230] ^ x[139];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[231] & ~t[232]);
  assign t[191] = (t[233] & ~t[234]);
  assign t[192] = (t[235] & ~t[236]);
  assign t[193] = (t[237] & ~t[238]);
  assign t[194] = (t[239] & ~t[240]);
  assign t[195] = (t[241] & ~t[242]);
  assign t[196] = (t[243] & ~t[244]);
  assign t[197] = (t[245] & ~t[246]);
  assign t[198] = (t[247] & ~t[248]);
  assign t[199] = (t[249] & ~t[250]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[251] & ~t[252]);
  assign t[201] = (t[253] & ~t[254]);
  assign t[202] = (t[255] & ~t[256]);
  assign t[203] = (t[257] & ~t[258]);
  assign t[204] = (t[259] & ~t[260]);
  assign t[205] = (t[261] & ~t[262]);
  assign t[206] = (t[263] & ~t[264]);
  assign t[207] = (t[265] & ~t[266]);
  assign t[208] = (t[267] & ~t[268]);
  assign t[209] = (t[269] & ~t[270]);
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = (t[271] & ~t[272]);
  assign t[211] = (t[273] & ~t[274]);
  assign t[212] = (t[275] & ~t[276]);
  assign t[213] = (t[277] & ~t[278]);
  assign t[214] = (t[279] & ~t[280]);
  assign t[215] = (t[281] & ~t[282]);
  assign t[216] = (t[283] & ~t[284]);
  assign t[217] = (t[285] & ~t[286]);
  assign t[218] = (t[287] & ~t[288]);
  assign t[219] = (t[289] & ~t[290]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[291] & ~t[292]);
  assign t[221] = (t[293] & ~t[294]);
  assign t[222] = (t[295] & ~t[296]);
  assign t[223] = (t[297] & ~t[298]);
  assign t[224] = (t[299] & ~t[300]);
  assign t[225] = (t[301] & ~t[302]);
  assign t[226] = (t[303] & ~t[304]);
  assign t[227] = (t[305] & ~t[306]);
  assign t[228] = (t[307] & ~t[308]);
  assign t[229] = (t[309] & ~t[310]);
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = (t[311] & ~t[312]);
  assign t[231] = t[313] ^ x[2];
  assign t[232] = t[314] ^ x[1];
  assign t[233] = t[315] ^ x[8];
  assign t[234] = t[316] ^ x[7];
  assign t[235] = t[317] ^ x[11];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[14];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[17];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[22];
  assign t[242] = t[324] ^ x[21];
  assign t[243] = t[325] ^ x[27];
  assign t[244] = t[326] ^ x[26];
  assign t[245] = t[327] ^ x[32];
  assign t[246] = t[328] ^ x[31];
  assign t[247] = t[329] ^ x[35];
  assign t[248] = t[330] ^ x[34];
  assign t[249] = t[331] ^ x[38];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[37];
  assign t[251] = t[333] ^ x[41];
  assign t[252] = t[334] ^ x[40];
  assign t[253] = t[335] ^ x[46];
  assign t[254] = t[336] ^ x[45];
  assign t[255] = t[337] ^ x[51];
  assign t[256] = t[338] ^ x[50];
  assign t[257] = t[339] ^ x[54];
  assign t[258] = t[340] ^ x[53];
  assign t[259] = t[341] ^ x[57];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[56];
  assign t[261] = t[343] ^ x[62];
  assign t[262] = t[344] ^ x[61];
  assign t[263] = t[345] ^ x[67];
  assign t[264] = t[346] ^ x[66];
  assign t[265] = t[347] ^ x[70];
  assign t[266] = t[348] ^ x[69];
  assign t[267] = t[349] ^ x[73];
  assign t[268] = t[350] ^ x[72];
  assign t[269] = t[351] ^ x[76];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[75];
  assign t[271] = t[353] ^ x[79];
  assign t[272] = t[354] ^ x[78];
  assign t[273] = t[355] ^ x[82];
  assign t[274] = t[356] ^ x[81];
  assign t[275] = t[357] ^ x[85];
  assign t[276] = t[358] ^ x[84];
  assign t[277] = t[359] ^ x[88];
  assign t[278] = t[360] ^ x[87];
  assign t[279] = t[361] ^ x[91];
  assign t[27] = ~(t[43] & t[113]);
  assign t[280] = t[362] ^ x[90];
  assign t[281] = t[363] ^ x[94];
  assign t[282] = t[364] ^ x[93];
  assign t[283] = t[365] ^ x[97];
  assign t[284] = t[366] ^ x[96];
  assign t[285] = t[367] ^ x[100];
  assign t[286] = t[368] ^ x[99];
  assign t[287] = t[369] ^ x[103];
  assign t[288] = t[370] ^ x[102];
  assign t[289] = t[371] ^ x[106];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[105];
  assign t[291] = t[373] ^ x[109];
  assign t[292] = t[374] ^ x[108];
  assign t[293] = t[375] ^ x[112];
  assign t[294] = t[376] ^ x[111];
  assign t[295] = t[377] ^ x[115];
  assign t[296] = t[378] ^ x[114];
  assign t[297] = t[379] ^ x[118];
  assign t[298] = t[380] ^ x[117];
  assign t[299] = t[381] ^ x[121];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[120];
  assign t[301] = t[383] ^ x[124];
  assign t[302] = t[384] ^ x[123];
  assign t[303] = t[385] ^ x[127];
  assign t[304] = t[386] ^ x[126];
  assign t[305] = t[387] ^ x[130];
  assign t[306] = t[388] ^ x[129];
  assign t[307] = t[389] ^ x[133];
  assign t[308] = t[390] ^ x[132];
  assign t[309] = t[391] ^ x[136];
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = t[392] ^ x[135];
  assign t[311] = t[393] ^ x[139];
  assign t[312] = t[394] ^ x[138];
  assign t[313] = (x[0]);
  assign t[314] = (x[0]);
  assign t[315] = (x[6]);
  assign t[316] = (x[6]);
  assign t[317] = (x[9]);
  assign t[318] = (x[9]);
  assign t[319] = (x[12]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[12]);
  assign t[321] = (x[15]);
  assign t[322] = (x[15]);
  assign t[323] = (x[20]);
  assign t[324] = (x[20]);
  assign t[325] = (x[25]);
  assign t[326] = (x[25]);
  assign t[327] = (x[30]);
  assign t[328] = (x[30]);
  assign t[329] = (x[33]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[33]);
  assign t[331] = (x[36]);
  assign t[332] = (x[36]);
  assign t[333] = (x[39]);
  assign t[334] = (x[39]);
  assign t[335] = (x[44]);
  assign t[336] = (x[44]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = t[52] ^ t[30];
  assign t[340] = (x[52]);
  assign t[341] = (x[55]);
  assign t[342] = (x[55]);
  assign t[343] = (x[60]);
  assign t[344] = (x[60]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[71]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[71]);
  assign t[351] = (x[74]);
  assign t[352] = (x[74]);
  assign t[353] = (x[77]);
  assign t[354] = (x[77]);
  assign t[355] = (x[80]);
  assign t[356] = (x[80]);
  assign t[357] = (x[83]);
  assign t[358] = (x[83]);
  assign t[359] = (x[86]);
  assign t[35] = ~(t[55] & t[114]);
  assign t[360] = (x[86]);
  assign t[361] = (x[89]);
  assign t[362] = (x[89]);
  assign t[363] = (x[92]);
  assign t[364] = (x[92]);
  assign t[365] = (x[95]);
  assign t[366] = (x[95]);
  assign t[367] = (x[98]);
  assign t[368] = (x[98]);
  assign t[369] = (x[101]);
  assign t[36] = t[111] ? x[29] : x[28];
  assign t[370] = (x[101]);
  assign t[371] = (x[104]);
  assign t[372] = (x[104]);
  assign t[373] = (x[107]);
  assign t[374] = (x[107]);
  assign t[375] = (x[110]);
  assign t[376] = (x[110]);
  assign t[377] = (x[113]);
  assign t[378] = (x[113]);
  assign t[379] = (x[116]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[116]);
  assign t[381] = (x[119]);
  assign t[382] = (x[119]);
  assign t[383] = (x[122]);
  assign t[384] = (x[122]);
  assign t[385] = (x[125]);
  assign t[386] = (x[125]);
  assign t[387] = (x[128]);
  assign t[388] = (x[128]);
  assign t[389] = (x[131]);
  assign t[38] = t[58] ^ t[59];
  assign t[390] = (x[131]);
  assign t[391] = (x[134]);
  assign t[392] = (x[134]);
  assign t[393] = (x[137]);
  assign t[394] = (x[137]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[115]);
  assign t[42] = ~(t[116]);
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69] & t[117]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[118]);
  assign t[49] = t[44] ? x[43] : x[42];
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[119]);
  assign t[52] = t[111] ? x[48] : x[47];
  assign t[53] = ~(t[120]);
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[76] & t[77]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[80] & t[122]);
  assign t[58] = t[111] ? x[59] : x[58];
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[123]);
  assign t[62] = t[44] ? x[64] : x[63];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[116] & t[115]);
  assign t[65] = ~(t[124]);
  assign t[66] = ~(t[111]);
  assign t[67] = ~(t[125]);
  assign t[68] = ~(t[126]);
  assign t[69] = ~(t[88] & t[89]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[92] & t[93]);
  assign t[76] = ~(t[121] & t[120]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[109] & t[110]);
  assign t[80] = ~(t[94] & t[95]);
  assign t[81] = ~(t[96] & t[97]);
  assign t[82] = ~(t[98] & t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[99] & t[100]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[137]);
  assign t[88] = ~(t[126] & t[125]);
  assign t[89] = ~(t[138]);
  assign t[8] = ~(t[111] & t[112]);
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[133] & t[132]);
  assign t[95] = ~(t[141]);
  assign t[96] = ~(t[142]);
  assign t[97] = ~(t[143]);
  assign t[98] = ~(t[104] & t[105]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [139:0] x;
 output y;

 wire [394:0] t;
  assign t[0] = t[1] ? t[2] : t[108];
  assign t[100] = ~(t[144]);
  assign t[101] = ~(t[145]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[106] & t[107]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[147]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[111] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = t[190] ^ x[2];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[8];
  assign t[151] = t[192] ^ x[11];
  assign t[152] = t[193] ^ x[14];
  assign t[153] = t[194] ^ x[17];
  assign t[154] = t[195] ^ x[22];
  assign t[155] = t[196] ^ x[27];
  assign t[156] = t[197] ^ x[32];
  assign t[157] = t[198] ^ x[35];
  assign t[158] = t[199] ^ x[38];
  assign t[159] = t[200] ^ x[41];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[46];
  assign t[161] = t[202] ^ x[51];
  assign t[162] = t[203] ^ x[54];
  assign t[163] = t[204] ^ x[57];
  assign t[164] = t[205] ^ x[62];
  assign t[165] = t[206] ^ x[67];
  assign t[166] = t[207] ^ x[70];
  assign t[167] = t[208] ^ x[73];
  assign t[168] = t[209] ^ x[76];
  assign t[169] = t[210] ^ x[79];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[82];
  assign t[171] = t[212] ^ x[85];
  assign t[172] = t[213] ^ x[88];
  assign t[173] = t[214] ^ x[91];
  assign t[174] = t[215] ^ x[94];
  assign t[175] = t[216] ^ x[97];
  assign t[176] = t[217] ^ x[100];
  assign t[177] = t[218] ^ x[103];
  assign t[178] = t[219] ^ x[106];
  assign t[179] = t[220] ^ x[109];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[112];
  assign t[181] = t[222] ^ x[115];
  assign t[182] = t[223] ^ x[118];
  assign t[183] = t[224] ^ x[121];
  assign t[184] = t[225] ^ x[124];
  assign t[185] = t[226] ^ x[127];
  assign t[186] = t[227] ^ x[130];
  assign t[187] = t[228] ^ x[133];
  assign t[188] = t[229] ^ x[136];
  assign t[189] = t[230] ^ x[139];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[231] & ~t[232]);
  assign t[191] = (t[233] & ~t[234]);
  assign t[192] = (t[235] & ~t[236]);
  assign t[193] = (t[237] & ~t[238]);
  assign t[194] = (t[239] & ~t[240]);
  assign t[195] = (t[241] & ~t[242]);
  assign t[196] = (t[243] & ~t[244]);
  assign t[197] = (t[245] & ~t[246]);
  assign t[198] = (t[247] & ~t[248]);
  assign t[199] = (t[249] & ~t[250]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[251] & ~t[252]);
  assign t[201] = (t[253] & ~t[254]);
  assign t[202] = (t[255] & ~t[256]);
  assign t[203] = (t[257] & ~t[258]);
  assign t[204] = (t[259] & ~t[260]);
  assign t[205] = (t[261] & ~t[262]);
  assign t[206] = (t[263] & ~t[264]);
  assign t[207] = (t[265] & ~t[266]);
  assign t[208] = (t[267] & ~t[268]);
  assign t[209] = (t[269] & ~t[270]);
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = (t[271] & ~t[272]);
  assign t[211] = (t[273] & ~t[274]);
  assign t[212] = (t[275] & ~t[276]);
  assign t[213] = (t[277] & ~t[278]);
  assign t[214] = (t[279] & ~t[280]);
  assign t[215] = (t[281] & ~t[282]);
  assign t[216] = (t[283] & ~t[284]);
  assign t[217] = (t[285] & ~t[286]);
  assign t[218] = (t[287] & ~t[288]);
  assign t[219] = (t[289] & ~t[290]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[291] & ~t[292]);
  assign t[221] = (t[293] & ~t[294]);
  assign t[222] = (t[295] & ~t[296]);
  assign t[223] = (t[297] & ~t[298]);
  assign t[224] = (t[299] & ~t[300]);
  assign t[225] = (t[301] & ~t[302]);
  assign t[226] = (t[303] & ~t[304]);
  assign t[227] = (t[305] & ~t[306]);
  assign t[228] = (t[307] & ~t[308]);
  assign t[229] = (t[309] & ~t[310]);
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = (t[311] & ~t[312]);
  assign t[231] = t[313] ^ x[2];
  assign t[232] = t[314] ^ x[1];
  assign t[233] = t[315] ^ x[8];
  assign t[234] = t[316] ^ x[7];
  assign t[235] = t[317] ^ x[11];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[14];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[17];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[22];
  assign t[242] = t[324] ^ x[21];
  assign t[243] = t[325] ^ x[27];
  assign t[244] = t[326] ^ x[26];
  assign t[245] = t[327] ^ x[32];
  assign t[246] = t[328] ^ x[31];
  assign t[247] = t[329] ^ x[35];
  assign t[248] = t[330] ^ x[34];
  assign t[249] = t[331] ^ x[38];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[37];
  assign t[251] = t[333] ^ x[41];
  assign t[252] = t[334] ^ x[40];
  assign t[253] = t[335] ^ x[46];
  assign t[254] = t[336] ^ x[45];
  assign t[255] = t[337] ^ x[51];
  assign t[256] = t[338] ^ x[50];
  assign t[257] = t[339] ^ x[54];
  assign t[258] = t[340] ^ x[53];
  assign t[259] = t[341] ^ x[57];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[56];
  assign t[261] = t[343] ^ x[62];
  assign t[262] = t[344] ^ x[61];
  assign t[263] = t[345] ^ x[67];
  assign t[264] = t[346] ^ x[66];
  assign t[265] = t[347] ^ x[70];
  assign t[266] = t[348] ^ x[69];
  assign t[267] = t[349] ^ x[73];
  assign t[268] = t[350] ^ x[72];
  assign t[269] = t[351] ^ x[76];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[75];
  assign t[271] = t[353] ^ x[79];
  assign t[272] = t[354] ^ x[78];
  assign t[273] = t[355] ^ x[82];
  assign t[274] = t[356] ^ x[81];
  assign t[275] = t[357] ^ x[85];
  assign t[276] = t[358] ^ x[84];
  assign t[277] = t[359] ^ x[88];
  assign t[278] = t[360] ^ x[87];
  assign t[279] = t[361] ^ x[91];
  assign t[27] = ~(t[43] & t[113]);
  assign t[280] = t[362] ^ x[90];
  assign t[281] = t[363] ^ x[94];
  assign t[282] = t[364] ^ x[93];
  assign t[283] = t[365] ^ x[97];
  assign t[284] = t[366] ^ x[96];
  assign t[285] = t[367] ^ x[100];
  assign t[286] = t[368] ^ x[99];
  assign t[287] = t[369] ^ x[103];
  assign t[288] = t[370] ^ x[102];
  assign t[289] = t[371] ^ x[106];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[105];
  assign t[291] = t[373] ^ x[109];
  assign t[292] = t[374] ^ x[108];
  assign t[293] = t[375] ^ x[112];
  assign t[294] = t[376] ^ x[111];
  assign t[295] = t[377] ^ x[115];
  assign t[296] = t[378] ^ x[114];
  assign t[297] = t[379] ^ x[118];
  assign t[298] = t[380] ^ x[117];
  assign t[299] = t[381] ^ x[121];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[120];
  assign t[301] = t[383] ^ x[124];
  assign t[302] = t[384] ^ x[123];
  assign t[303] = t[385] ^ x[127];
  assign t[304] = t[386] ^ x[126];
  assign t[305] = t[387] ^ x[130];
  assign t[306] = t[388] ^ x[129];
  assign t[307] = t[389] ^ x[133];
  assign t[308] = t[390] ^ x[132];
  assign t[309] = t[391] ^ x[136];
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = t[392] ^ x[135];
  assign t[311] = t[393] ^ x[139];
  assign t[312] = t[394] ^ x[138];
  assign t[313] = (x[0]);
  assign t[314] = (x[0]);
  assign t[315] = (x[6]);
  assign t[316] = (x[6]);
  assign t[317] = (x[9]);
  assign t[318] = (x[9]);
  assign t[319] = (x[12]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[12]);
  assign t[321] = (x[15]);
  assign t[322] = (x[15]);
  assign t[323] = (x[20]);
  assign t[324] = (x[20]);
  assign t[325] = (x[25]);
  assign t[326] = (x[25]);
  assign t[327] = (x[30]);
  assign t[328] = (x[30]);
  assign t[329] = (x[33]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[33]);
  assign t[331] = (x[36]);
  assign t[332] = (x[36]);
  assign t[333] = (x[39]);
  assign t[334] = (x[39]);
  assign t[335] = (x[44]);
  assign t[336] = (x[44]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = t[52] ^ t[30];
  assign t[340] = (x[52]);
  assign t[341] = (x[55]);
  assign t[342] = (x[55]);
  assign t[343] = (x[60]);
  assign t[344] = (x[60]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[71]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[71]);
  assign t[351] = (x[74]);
  assign t[352] = (x[74]);
  assign t[353] = (x[77]);
  assign t[354] = (x[77]);
  assign t[355] = (x[80]);
  assign t[356] = (x[80]);
  assign t[357] = (x[83]);
  assign t[358] = (x[83]);
  assign t[359] = (x[86]);
  assign t[35] = ~(t[55] & t[114]);
  assign t[360] = (x[86]);
  assign t[361] = (x[89]);
  assign t[362] = (x[89]);
  assign t[363] = (x[92]);
  assign t[364] = (x[92]);
  assign t[365] = (x[95]);
  assign t[366] = (x[95]);
  assign t[367] = (x[98]);
  assign t[368] = (x[98]);
  assign t[369] = (x[101]);
  assign t[36] = t[111] ? x[29] : x[28];
  assign t[370] = (x[101]);
  assign t[371] = (x[104]);
  assign t[372] = (x[104]);
  assign t[373] = (x[107]);
  assign t[374] = (x[107]);
  assign t[375] = (x[110]);
  assign t[376] = (x[110]);
  assign t[377] = (x[113]);
  assign t[378] = (x[113]);
  assign t[379] = (x[116]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[116]);
  assign t[381] = (x[119]);
  assign t[382] = (x[119]);
  assign t[383] = (x[122]);
  assign t[384] = (x[122]);
  assign t[385] = (x[125]);
  assign t[386] = (x[125]);
  assign t[387] = (x[128]);
  assign t[388] = (x[128]);
  assign t[389] = (x[131]);
  assign t[38] = t[58] ^ t[59];
  assign t[390] = (x[131]);
  assign t[391] = (x[134]);
  assign t[392] = (x[134]);
  assign t[393] = (x[137]);
  assign t[394] = (x[137]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[115]);
  assign t[42] = ~(t[116]);
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69] & t[117]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[118]);
  assign t[49] = t[44] ? x[43] : x[42];
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[119]);
  assign t[52] = t[111] ? x[48] : x[47];
  assign t[53] = ~(t[120]);
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[76] & t[77]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[80] & t[122]);
  assign t[58] = t[111] ? x[59] : x[58];
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[123]);
  assign t[62] = t[44] ? x[64] : x[63];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[116] & t[115]);
  assign t[65] = ~(t[124]);
  assign t[66] = ~(t[111]);
  assign t[67] = ~(t[125]);
  assign t[68] = ~(t[126]);
  assign t[69] = ~(t[88] & t[89]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[92] & t[93]);
  assign t[76] = ~(t[121] & t[120]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[109] & t[110]);
  assign t[80] = ~(t[94] & t[95]);
  assign t[81] = ~(t[96] & t[97]);
  assign t[82] = ~(t[98] & t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[99] & t[100]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[137]);
  assign t[88] = ~(t[126] & t[125]);
  assign t[89] = ~(t[138]);
  assign t[8] = ~(t[111] & t[112]);
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[133] & t[132]);
  assign t[95] = ~(t[141]);
  assign t[96] = ~(t[142]);
  assign t[97] = ~(t[143]);
  assign t[98] = ~(t[104] & t[105]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [139:0] x;
 output y;

 wire [386:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[2];
  assign t[142] = t[183] ^ x[8];
  assign t[143] = t[184] ^ x[11];
  assign t[144] = t[185] ^ x[14];
  assign t[145] = t[186] ^ x[17];
  assign t[146] = t[187] ^ x[22];
  assign t[147] = t[188] ^ x[27];
  assign t[148] = t[189] ^ x[32];
  assign t[149] = t[190] ^ x[35];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[38];
  assign t[151] = t[192] ^ x[41];
  assign t[152] = t[193] ^ x[46];
  assign t[153] = t[194] ^ x[51];
  assign t[154] = t[195] ^ x[54];
  assign t[155] = t[196] ^ x[57];
  assign t[156] = t[197] ^ x[62];
  assign t[157] = t[198] ^ x[67];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[73];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[76];
  assign t[161] = t[202] ^ x[79];
  assign t[162] = t[203] ^ x[82];
  assign t[163] = t[204] ^ x[85];
  assign t[164] = t[205] ^ x[88];
  assign t[165] = t[206] ^ x[91];
  assign t[166] = t[207] ^ x[94];
  assign t[167] = t[208] ^ x[97];
  assign t[168] = t[209] ^ x[100];
  assign t[169] = t[210] ^ x[103];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[106];
  assign t[171] = t[212] ^ x[109];
  assign t[172] = t[213] ^ x[112];
  assign t[173] = t[214] ^ x[115];
  assign t[174] = t[215] ^ x[118];
  assign t[175] = t[216] ^ x[121];
  assign t[176] = t[217] ^ x[124];
  assign t[177] = t[218] ^ x[127];
  assign t[178] = t[219] ^ x[130];
  assign t[179] = t[220] ^ x[133];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[136];
  assign t[181] = t[222] ^ x[139];
  assign t[182] = (t[223] & ~t[224]);
  assign t[183] = (t[225] & ~t[226]);
  assign t[184] = (t[227] & ~t[228]);
  assign t[185] = (t[229] & ~t[230]);
  assign t[186] = (t[231] & ~t[232]);
  assign t[187] = (t[233] & ~t[234]);
  assign t[188] = (t[235] & ~t[236]);
  assign t[189] = (t[237] & ~t[238]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[239] & ~t[240]);
  assign t[191] = (t[241] & ~t[242]);
  assign t[192] = (t[243] & ~t[244]);
  assign t[193] = (t[245] & ~t[246]);
  assign t[194] = (t[247] & ~t[248]);
  assign t[195] = (t[249] & ~t[250]);
  assign t[196] = (t[251] & ~t[252]);
  assign t[197] = (t[253] & ~t[254]);
  assign t[198] = (t[255] & ~t[256]);
  assign t[199] = (t[257] & ~t[258]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[259] & ~t[260]);
  assign t[201] = (t[261] & ~t[262]);
  assign t[202] = (t[263] & ~t[264]);
  assign t[203] = (t[265] & ~t[266]);
  assign t[204] = (t[267] & ~t[268]);
  assign t[205] = (t[269] & ~t[270]);
  assign t[206] = (t[271] & ~t[272]);
  assign t[207] = (t[273] & ~t[274]);
  assign t[208] = (t[275] & ~t[276]);
  assign t[209] = (t[277] & ~t[278]);
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = (t[279] & ~t[280]);
  assign t[211] = (t[281] & ~t[282]);
  assign t[212] = (t[283] & ~t[284]);
  assign t[213] = (t[285] & ~t[286]);
  assign t[214] = (t[287] & ~t[288]);
  assign t[215] = (t[289] & ~t[290]);
  assign t[216] = (t[291] & ~t[292]);
  assign t[217] = (t[293] & ~t[294]);
  assign t[218] = (t[295] & ~t[296]);
  assign t[219] = (t[297] & ~t[298]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[299] & ~t[300]);
  assign t[221] = (t[301] & ~t[302]);
  assign t[222] = (t[303] & ~t[304]);
  assign t[223] = t[305] ^ x[2];
  assign t[224] = t[306] ^ x[1];
  assign t[225] = t[307] ^ x[8];
  assign t[226] = t[308] ^ x[7];
  assign t[227] = t[309] ^ x[11];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[14];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[17];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[22];
  assign t[234] = t[316] ^ x[21];
  assign t[235] = t[317] ^ x[27];
  assign t[236] = t[318] ^ x[26];
  assign t[237] = t[319] ^ x[32];
  assign t[238] = t[320] ^ x[31];
  assign t[239] = t[321] ^ x[35];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[322] ^ x[34];
  assign t[241] = t[323] ^ x[38];
  assign t[242] = t[324] ^ x[37];
  assign t[243] = t[325] ^ x[41];
  assign t[244] = t[326] ^ x[40];
  assign t[245] = t[327] ^ x[46];
  assign t[246] = t[328] ^ x[45];
  assign t[247] = t[329] ^ x[51];
  assign t[248] = t[330] ^ x[50];
  assign t[249] = t[331] ^ x[54];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[53];
  assign t[251] = t[333] ^ x[57];
  assign t[252] = t[334] ^ x[56];
  assign t[253] = t[335] ^ x[62];
  assign t[254] = t[336] ^ x[61];
  assign t[255] = t[337] ^ x[67];
  assign t[256] = t[338] ^ x[66];
  assign t[257] = t[339] ^ x[70];
  assign t[258] = t[340] ^ x[69];
  assign t[259] = t[341] ^ x[73];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[72];
  assign t[261] = t[343] ^ x[76];
  assign t[262] = t[344] ^ x[75];
  assign t[263] = t[345] ^ x[79];
  assign t[264] = t[346] ^ x[78];
  assign t[265] = t[347] ^ x[82];
  assign t[266] = t[348] ^ x[81];
  assign t[267] = t[349] ^ x[85];
  assign t[268] = t[350] ^ x[84];
  assign t[269] = t[351] ^ x[88];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[87];
  assign t[271] = t[353] ^ x[91];
  assign t[272] = t[354] ^ x[90];
  assign t[273] = t[355] ^ x[94];
  assign t[274] = t[356] ^ x[93];
  assign t[275] = t[357] ^ x[97];
  assign t[276] = t[358] ^ x[96];
  assign t[277] = t[359] ^ x[100];
  assign t[278] = t[360] ^ x[99];
  assign t[279] = t[361] ^ x[103];
  assign t[27] = t[43] | t[105];
  assign t[280] = t[362] ^ x[102];
  assign t[281] = t[363] ^ x[106];
  assign t[282] = t[364] ^ x[105];
  assign t[283] = t[365] ^ x[109];
  assign t[284] = t[366] ^ x[108];
  assign t[285] = t[367] ^ x[112];
  assign t[286] = t[368] ^ x[111];
  assign t[287] = t[369] ^ x[115];
  assign t[288] = t[370] ^ x[114];
  assign t[289] = t[371] ^ x[118];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[117];
  assign t[291] = t[373] ^ x[121];
  assign t[292] = t[374] ^ x[120];
  assign t[293] = t[375] ^ x[124];
  assign t[294] = t[376] ^ x[123];
  assign t[295] = t[377] ^ x[127];
  assign t[296] = t[378] ^ x[126];
  assign t[297] = t[379] ^ x[130];
  assign t[298] = t[380] ^ x[129];
  assign t[299] = t[381] ^ x[133];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[132];
  assign t[301] = t[383] ^ x[136];
  assign t[302] = t[384] ^ x[135];
  assign t[303] = t[385] ^ x[139];
  assign t[304] = t[386] ^ x[138];
  assign t[305] = (x[0]);
  assign t[306] = (x[0]);
  assign t[307] = (x[6]);
  assign t[308] = (x[6]);
  assign t[309] = (x[9]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = (x[9]);
  assign t[311] = (x[12]);
  assign t[312] = (x[12]);
  assign t[313] = (x[15]);
  assign t[314] = (x[15]);
  assign t[315] = (x[20]);
  assign t[316] = (x[20]);
  assign t[317] = (x[25]);
  assign t[318] = (x[25]);
  assign t[319] = (x[30]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[30]);
  assign t[321] = (x[33]);
  assign t[322] = (x[33]);
  assign t[323] = (x[36]);
  assign t[324] = (x[36]);
  assign t[325] = (x[39]);
  assign t[326] = (x[39]);
  assign t[327] = (x[44]);
  assign t[328] = (x[44]);
  assign t[329] = (x[49]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[49]);
  assign t[331] = (x[52]);
  assign t[332] = (x[52]);
  assign t[333] = (x[55]);
  assign t[334] = (x[55]);
  assign t[335] = (x[60]);
  assign t[336] = (x[60]);
  assign t[337] = (x[65]);
  assign t[338] = (x[65]);
  assign t[339] = (x[68]);
  assign t[33] = t[52] ^ t[30];
  assign t[340] = (x[68]);
  assign t[341] = (x[71]);
  assign t[342] = (x[71]);
  assign t[343] = (x[74]);
  assign t[344] = (x[74]);
  assign t[345] = (x[77]);
  assign t[346] = (x[77]);
  assign t[347] = (x[80]);
  assign t[348] = (x[80]);
  assign t[349] = (x[83]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[83]);
  assign t[351] = (x[86]);
  assign t[352] = (x[86]);
  assign t[353] = (x[89]);
  assign t[354] = (x[89]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[98]);
  assign t[35] = t[55] | t[106];
  assign t[360] = (x[98]);
  assign t[361] = (x[101]);
  assign t[362] = (x[101]);
  assign t[363] = (x[104]);
  assign t[364] = (x[104]);
  assign t[365] = (x[107]);
  assign t[366] = (x[107]);
  assign t[367] = (x[110]);
  assign t[368] = (x[110]);
  assign t[369] = (x[113]);
  assign t[36] = t[103] ? x[29] : x[28];
  assign t[370] = (x[113]);
  assign t[371] = (x[116]);
  assign t[372] = (x[116]);
  assign t[373] = (x[119]);
  assign t[374] = (x[119]);
  assign t[375] = (x[122]);
  assign t[376] = (x[122]);
  assign t[377] = (x[125]);
  assign t[378] = (x[125]);
  assign t[379] = (x[128]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[128]);
  assign t[381] = (x[131]);
  assign t[382] = (x[131]);
  assign t[383] = (x[134]);
  assign t[384] = (x[134]);
  assign t[385] = (x[137]);
  assign t[386] = (x[137]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[64] | t[41]);
  assign t[44] = ~(t[65]);
  assign t[45] = ~(t[66] & t[67]);
  assign t[46] = t[68] | t[109];
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[110];
  assign t[49] = t[44] ? x[43] : x[42];
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[111];
  assign t[52] = t[44] ? x[48] : x[47];
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[113]);
  assign t[55] = ~(t[75] | t[53]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[114];
  assign t[58] = t[103] ? x[59] : x[58];
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[115];
  assign t[62] = t[84] ? x[64] : x[63];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[116]);
  assign t[65] = ~(t[103]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[87] | t[66]);
  assign t[69] = ~(t[119]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[88] | t[69]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[89] | t[72]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[90] | t[76]);
  assign t[79] = ~(t[91] & t[92]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = t[93] | t[126];
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[94] | t[81]);
  assign t[84] = ~(t[65]);
  assign t[85] = ~(t[95] & t[96]);
  assign t[86] = t[97] | t[129];
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[98] | t[91]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[99] | t[95]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind171(x, y);
 input [139:0] x;
 output y;

 wire [386:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[18] : x[19];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[2];
  assign t[142] = t[183] ^ x[8];
  assign t[143] = t[184] ^ x[11];
  assign t[144] = t[185] ^ x[14];
  assign t[145] = t[186] ^ x[17];
  assign t[146] = t[187] ^ x[22];
  assign t[147] = t[188] ^ x[27];
  assign t[148] = t[189] ^ x[32];
  assign t[149] = t[190] ^ x[35];
  assign t[14] = x[4] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[38];
  assign t[151] = t[192] ^ x[41];
  assign t[152] = t[193] ^ x[46];
  assign t[153] = t[194] ^ x[51];
  assign t[154] = t[195] ^ x[54];
  assign t[155] = t[196] ^ x[57];
  assign t[156] = t[197] ^ x[62];
  assign t[157] = t[198] ^ x[67];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[73];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[76];
  assign t[161] = t[202] ^ x[79];
  assign t[162] = t[203] ^ x[82];
  assign t[163] = t[204] ^ x[85];
  assign t[164] = t[205] ^ x[88];
  assign t[165] = t[206] ^ x[91];
  assign t[166] = t[207] ^ x[94];
  assign t[167] = t[208] ^ x[97];
  assign t[168] = t[209] ^ x[100];
  assign t[169] = t[210] ^ x[103];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[106];
  assign t[171] = t[212] ^ x[109];
  assign t[172] = t[213] ^ x[112];
  assign t[173] = t[214] ^ x[115];
  assign t[174] = t[215] ^ x[118];
  assign t[175] = t[216] ^ x[121];
  assign t[176] = t[217] ^ x[124];
  assign t[177] = t[218] ^ x[127];
  assign t[178] = t[219] ^ x[130];
  assign t[179] = t[220] ^ x[133];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[136];
  assign t[181] = t[222] ^ x[139];
  assign t[182] = (t[223] & ~t[224]);
  assign t[183] = (t[225] & ~t[226]);
  assign t[184] = (t[227] & ~t[228]);
  assign t[185] = (t[229] & ~t[230]);
  assign t[186] = (t[231] & ~t[232]);
  assign t[187] = (t[233] & ~t[234]);
  assign t[188] = (t[235] & ~t[236]);
  assign t[189] = (t[237] & ~t[238]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (t[239] & ~t[240]);
  assign t[191] = (t[241] & ~t[242]);
  assign t[192] = (t[243] & ~t[244]);
  assign t[193] = (t[245] & ~t[246]);
  assign t[194] = (t[247] & ~t[248]);
  assign t[195] = (t[249] & ~t[250]);
  assign t[196] = (t[251] & ~t[252]);
  assign t[197] = (t[253] & ~t[254]);
  assign t[198] = (t[255] & ~t[256]);
  assign t[199] = (t[257] & ~t[258]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[259] & ~t[260]);
  assign t[201] = (t[261] & ~t[262]);
  assign t[202] = (t[263] & ~t[264]);
  assign t[203] = (t[265] & ~t[266]);
  assign t[204] = (t[267] & ~t[268]);
  assign t[205] = (t[269] & ~t[270]);
  assign t[206] = (t[271] & ~t[272]);
  assign t[207] = (t[273] & ~t[274]);
  assign t[208] = (t[275] & ~t[276]);
  assign t[209] = (t[277] & ~t[278]);
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[210] = (t[279] & ~t[280]);
  assign t[211] = (t[281] & ~t[282]);
  assign t[212] = (t[283] & ~t[284]);
  assign t[213] = (t[285] & ~t[286]);
  assign t[214] = (t[287] & ~t[288]);
  assign t[215] = (t[289] & ~t[290]);
  assign t[216] = (t[291] & ~t[292]);
  assign t[217] = (t[293] & ~t[294]);
  assign t[218] = (t[295] & ~t[296]);
  assign t[219] = (t[297] & ~t[298]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[299] & ~t[300]);
  assign t[221] = (t[301] & ~t[302]);
  assign t[222] = (t[303] & ~t[304]);
  assign t[223] = t[305] ^ x[2];
  assign t[224] = t[306] ^ x[1];
  assign t[225] = t[307] ^ x[8];
  assign t[226] = t[308] ^ x[7];
  assign t[227] = t[309] ^ x[11];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[14];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[17];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[22];
  assign t[234] = t[316] ^ x[21];
  assign t[235] = t[317] ^ x[27];
  assign t[236] = t[318] ^ x[26];
  assign t[237] = t[319] ^ x[32];
  assign t[238] = t[320] ^ x[31];
  assign t[239] = t[321] ^ x[35];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[322] ^ x[34];
  assign t[241] = t[323] ^ x[38];
  assign t[242] = t[324] ^ x[37];
  assign t[243] = t[325] ^ x[41];
  assign t[244] = t[326] ^ x[40];
  assign t[245] = t[327] ^ x[46];
  assign t[246] = t[328] ^ x[45];
  assign t[247] = t[329] ^ x[51];
  assign t[248] = t[330] ^ x[50];
  assign t[249] = t[331] ^ x[54];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[332] ^ x[53];
  assign t[251] = t[333] ^ x[57];
  assign t[252] = t[334] ^ x[56];
  assign t[253] = t[335] ^ x[62];
  assign t[254] = t[336] ^ x[61];
  assign t[255] = t[337] ^ x[67];
  assign t[256] = t[338] ^ x[66];
  assign t[257] = t[339] ^ x[70];
  assign t[258] = t[340] ^ x[69];
  assign t[259] = t[341] ^ x[73];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[342] ^ x[72];
  assign t[261] = t[343] ^ x[76];
  assign t[262] = t[344] ^ x[75];
  assign t[263] = t[345] ^ x[79];
  assign t[264] = t[346] ^ x[78];
  assign t[265] = t[347] ^ x[82];
  assign t[266] = t[348] ^ x[81];
  assign t[267] = t[349] ^ x[85];
  assign t[268] = t[350] ^ x[84];
  assign t[269] = t[351] ^ x[88];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[352] ^ x[87];
  assign t[271] = t[353] ^ x[91];
  assign t[272] = t[354] ^ x[90];
  assign t[273] = t[355] ^ x[94];
  assign t[274] = t[356] ^ x[93];
  assign t[275] = t[357] ^ x[97];
  assign t[276] = t[358] ^ x[96];
  assign t[277] = t[359] ^ x[100];
  assign t[278] = t[360] ^ x[99];
  assign t[279] = t[361] ^ x[103];
  assign t[27] = t[43] | t[105];
  assign t[280] = t[362] ^ x[102];
  assign t[281] = t[363] ^ x[106];
  assign t[282] = t[364] ^ x[105];
  assign t[283] = t[365] ^ x[109];
  assign t[284] = t[366] ^ x[108];
  assign t[285] = t[367] ^ x[112];
  assign t[286] = t[368] ^ x[111];
  assign t[287] = t[369] ^ x[115];
  assign t[288] = t[370] ^ x[114];
  assign t[289] = t[371] ^ x[118];
  assign t[28] = t[44] ? x[24] : x[23];
  assign t[290] = t[372] ^ x[117];
  assign t[291] = t[373] ^ x[121];
  assign t[292] = t[374] ^ x[120];
  assign t[293] = t[375] ^ x[124];
  assign t[294] = t[376] ^ x[123];
  assign t[295] = t[377] ^ x[127];
  assign t[296] = t[378] ^ x[126];
  assign t[297] = t[379] ^ x[130];
  assign t[298] = t[380] ^ x[129];
  assign t[299] = t[381] ^ x[133];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[132];
  assign t[301] = t[383] ^ x[136];
  assign t[302] = t[384] ^ x[135];
  assign t[303] = t[385] ^ x[139];
  assign t[304] = t[386] ^ x[138];
  assign t[305] = (x[0]);
  assign t[306] = (x[0]);
  assign t[307] = (x[6]);
  assign t[308] = (x[6]);
  assign t[309] = (x[9]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = (x[9]);
  assign t[311] = (x[12]);
  assign t[312] = (x[12]);
  assign t[313] = (x[15]);
  assign t[314] = (x[15]);
  assign t[315] = (x[20]);
  assign t[316] = (x[20]);
  assign t[317] = (x[25]);
  assign t[318] = (x[25]);
  assign t[319] = (x[30]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[30]);
  assign t[321] = (x[33]);
  assign t[322] = (x[33]);
  assign t[323] = (x[36]);
  assign t[324] = (x[36]);
  assign t[325] = (x[39]);
  assign t[326] = (x[39]);
  assign t[327] = (x[44]);
  assign t[328] = (x[44]);
  assign t[329] = (x[49]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[49]);
  assign t[331] = (x[52]);
  assign t[332] = (x[52]);
  assign t[333] = (x[55]);
  assign t[334] = (x[55]);
  assign t[335] = (x[60]);
  assign t[336] = (x[60]);
  assign t[337] = (x[65]);
  assign t[338] = (x[65]);
  assign t[339] = (x[68]);
  assign t[33] = t[52] ^ t[30];
  assign t[340] = (x[68]);
  assign t[341] = (x[71]);
  assign t[342] = (x[71]);
  assign t[343] = (x[74]);
  assign t[344] = (x[74]);
  assign t[345] = (x[77]);
  assign t[346] = (x[77]);
  assign t[347] = (x[80]);
  assign t[348] = (x[80]);
  assign t[349] = (x[83]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[83]);
  assign t[351] = (x[86]);
  assign t[352] = (x[86]);
  assign t[353] = (x[89]);
  assign t[354] = (x[89]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[98]);
  assign t[35] = t[55] | t[106];
  assign t[360] = (x[98]);
  assign t[361] = (x[101]);
  assign t[362] = (x[101]);
  assign t[363] = (x[104]);
  assign t[364] = (x[104]);
  assign t[365] = (x[107]);
  assign t[366] = (x[107]);
  assign t[367] = (x[110]);
  assign t[368] = (x[110]);
  assign t[369] = (x[113]);
  assign t[36] = t[103] ? x[29] : x[28];
  assign t[370] = (x[113]);
  assign t[371] = (x[116]);
  assign t[372] = (x[116]);
  assign t[373] = (x[119]);
  assign t[374] = (x[119]);
  assign t[375] = (x[122]);
  assign t[376] = (x[122]);
  assign t[377] = (x[125]);
  assign t[378] = (x[125]);
  assign t[379] = (x[128]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[128]);
  assign t[381] = (x[131]);
  assign t[382] = (x[131]);
  assign t[383] = (x[134]);
  assign t[384] = (x[134]);
  assign t[385] = (x[137]);
  assign t[386] = (x[137]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[64] | t[41]);
  assign t[44] = ~(t[65]);
  assign t[45] = ~(t[66] & t[67]);
  assign t[46] = t[68] | t[109];
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[110];
  assign t[49] = t[44] ? x[43] : x[42];
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[111];
  assign t[52] = t[44] ? x[48] : x[47];
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[113]);
  assign t[55] = ~(t[75] | t[53]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[114];
  assign t[58] = t[103] ? x[59] : x[58];
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[115];
  assign t[62] = t[84] ? x[64] : x[63];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[116]);
  assign t[65] = ~(t[103]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[87] | t[66]);
  assign t[69] = ~(t[119]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[88] | t[69]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[89] | t[72]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[90] | t[76]);
  assign t[79] = ~(t[91] & t[92]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = t[93] | t[126];
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[94] | t[81]);
  assign t[84] = ~(t[65]);
  assign t[85] = ~(t[95] & t[96]);
  assign t[86] = t[97] | t[129];
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[98] | t[91]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[99] | t[95]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [151:0] x;
 output y;

 wire [519:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = t[144] | t[145];
  assign t[101] = ~(t[227]);
  assign t[102] = ~(t[228]);
  assign t[103] = ~(t[146] | t[147]);
  assign t[104] = ~(t[148] | t[149]);
  assign t[105] = ~(t[229] | t[150]);
  assign t[106] = t[143] ? x[87] : x[86];
  assign t[107] = ~(t[151] & t[152]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[155] | t[156]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[159] | t[160]);
  assign t[118] = ~(t[235] | t[161]);
  assign t[119] = t[30] ? x[107] : x[106];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[162] & t[163]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[164] | t[165]);
  assign t[124] = t[30] ? x[115] : x[114];
  assign t[125] = ~(t[166] & t[167]);
  assign t[126] = ~(t[128] | t[168]);
  assign t[127] = ~(t[86] | t[169]);
  assign t[128] = ~(t[208]);
  assign t[129] = ~(t[170] & t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[173] | t[174];
  assign t[132] = t[206] ? t[170] : t[175];
  assign t[133] = ~(t[173] & t[176]);
  assign t[134] = ~(t[174] & t[209]);
  assign t[135] = ~(t[173] & t[209]);
  assign t[136] = ~(t[174] & t[176]);
  assign t[137] = ~(t[238]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[207] | t[176]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[86] & t[206];
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[49]);
  assign t[144] = ~(t[177] & t[95]);
  assign t[145] = ~(t[86] | t[178]);
  assign t[146] = ~(t[240]);
  assign t[147] = ~(t[227] | t[228]);
  assign t[148] = ~(t[241]);
  assign t[149] = ~(t[242]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[179] | t[180]);
  assign t[151] = ~(t[52]);
  assign t[152] = ~(t[181] | t[145]);
  assign t[153] = ~(t[243]);
  assign t[154] = ~(t[231] | t[232]);
  assign t[155] = ~(t[86] | t[182]);
  assign t[156] = ~(t[32] & t[85]);
  assign t[157] = ~(t[244]);
  assign t[158] = ~(t[233] | t[234]);
  assign t[159] = ~(t[245]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[246]);
  assign t[161] = ~(t[183] | t[184]);
  assign t[162] = ~(t[52] | t[185]);
  assign t[163] = ~(t[100] | t[186]);
  assign t[164] = ~(t[247]);
  assign t[165] = ~(t[236] | t[237]);
  assign t[166] = ~(t[187] | t[155]);
  assign t[167] = ~(t[126] | t[144]);
  assign t[168] = t[206] ? t[133] : t[136];
  assign t[169] = t[206] ? t[175] : t[188];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(x[4] & t[189]);
  assign t[171] = ~(t[209] & t[190]);
  assign t[172] = ~(t[128] | t[206]);
  assign t[173] = ~(x[4] | t[207]);
  assign t[174] = x[4] & t[207];
  assign t[175] = ~(t[190] & t[176]);
  assign t[176] = ~(t[209]);
  assign t[177] = ~(t[191] | t[192]);
  assign t[178] = t[206] ? t[171] : t[170];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[241] | t[242]);
  assign t[181] = ~(t[193]);
  assign t[182] = t[206] ? t[135] : t[136];
  assign t[183] = ~(t[249]);
  assign t[184] = ~(t[245] | t[246]);
  assign t[185] = ~(t[86] | t[194]);
  assign t[186] = ~(t[195] & t[85]);
  assign t[187] = ~(t[86] | t[196]);
  assign t[188] = ~(x[4] & t[139]);
  assign t[189] = ~(t[207] | t[209]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(x[4] | t[197]);
  assign t[191] = ~(t[128] | t[198]);
  assign t[192] = ~(t[128] | t[199]);
  assign t[193] = ~(t[200] | t[53]);
  assign t[194] = t[206] ? t[170] : t[171];
  assign t[195] = ~(t[201] | t[200]);
  assign t[196] = t[206] ? t[133] : t[134];
  assign t[197] = ~(t[207]);
  assign t[198] = t[206] ? t[136] : t[133];
  assign t[199] = t[206] ? t[175] : t[170];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[86] | t[202]);
  assign t[201] = ~(t[203]);
  assign t[202] = t[206] ? t[188] : t[175];
  assign t[203] = ~(t[172] & t[204]);
  assign t[204] = ~(t[171] & t[188]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[2];
  assign t[251] = t[296] ^ x[10];
  assign t[252] = t[297] ^ x[13];
  assign t[253] = t[298] ^ x[16];
  assign t[254] = t[299] ^ x[19];
  assign t[255] = t[300] ^ x[22];
  assign t[256] = t[301] ^ x[25];
  assign t[257] = t[302] ^ x[28];
  assign t[258] = t[303] ^ x[31];
  assign t[259] = t[304] ^ x[34];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[39];
  assign t[261] = t[306] ^ x[42];
  assign t[262] = t[307] ^ x[45];
  assign t[263] = t[308] ^ x[48];
  assign t[264] = t[309] ^ x[51];
  assign t[265] = t[310] ^ x[56];
  assign t[266] = t[311] ^ x[59];
  assign t[267] = t[312] ^ x[62];
  assign t[268] = t[313] ^ x[65];
  assign t[269] = t[314] ^ x[68];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[71];
  assign t[271] = t[316] ^ x[74];
  assign t[272] = t[317] ^ x[79];
  assign t[273] = t[318] ^ x[82];
  assign t[274] = t[319] ^ x[85];
  assign t[275] = t[320] ^ x[90];
  assign t[276] = t[321] ^ x[93];
  assign t[277] = t[322] ^ x[96];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[102];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[105];
  assign t[281] = t[326] ^ x[110];
  assign t[282] = t[327] ^ x[113];
  assign t[283] = t[328] ^ x[118];
  assign t[284] = t[329] ^ x[121];
  assign t[285] = t[330] ^ x[124];
  assign t[286] = t[331] ^ x[127];
  assign t[287] = t[332] ^ x[130];
  assign t[288] = t[333] ^ x[133];
  assign t[289] = t[334] ^ x[136];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[139];
  assign t[291] = t[336] ^ x[142];
  assign t[292] = t[337] ^ x[145];
  assign t[293] = t[338] ^ x[148];
  assign t[294] = t[339] ^ x[151];
  assign t[295] = (t[340] & ~t[341]);
  assign t[296] = (t[342] & ~t[343]);
  assign t[297] = (t[344] & ~t[345]);
  assign t[298] = (t[346] & ~t[347]);
  assign t[299] = (t[348] & ~t[349]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[350] & ~t[351]);
  assign t[301] = (t[352] & ~t[353]);
  assign t[302] = (t[354] & ~t[355]);
  assign t[303] = (t[356] & ~t[357]);
  assign t[304] = (t[358] & ~t[359]);
  assign t[305] = (t[360] & ~t[361]);
  assign t[306] = (t[362] & ~t[363]);
  assign t[307] = (t[364] & ~t[365]);
  assign t[308] = (t[366] & ~t[367]);
  assign t[309] = (t[368] & ~t[369]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[370] & ~t[371]);
  assign t[311] = (t[372] & ~t[373]);
  assign t[312] = (t[374] & ~t[375]);
  assign t[313] = (t[376] & ~t[377]);
  assign t[314] = (t[378] & ~t[379]);
  assign t[315] = (t[380] & ~t[381]);
  assign t[316] = (t[382] & ~t[383]);
  assign t[317] = (t[384] & ~t[385]);
  assign t[318] = (t[386] & ~t[387]);
  assign t[319] = (t[388] & ~t[389]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[390] & ~t[391]);
  assign t[321] = (t[392] & ~t[393]);
  assign t[322] = (t[394] & ~t[395]);
  assign t[323] = (t[396] & ~t[397]);
  assign t[324] = (t[398] & ~t[399]);
  assign t[325] = (t[400] & ~t[401]);
  assign t[326] = (t[402] & ~t[403]);
  assign t[327] = (t[404] & ~t[405]);
  assign t[328] = (t[406] & ~t[407]);
  assign t[329] = (t[408] & ~t[409]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[410] & ~t[411]);
  assign t[331] = (t[412] & ~t[413]);
  assign t[332] = (t[414] & ~t[415]);
  assign t[333] = (t[416] & ~t[417]);
  assign t[334] = (t[418] & ~t[419]);
  assign t[335] = (t[420] & ~t[421]);
  assign t[336] = (t[422] & ~t[423]);
  assign t[337] = (t[424] & ~t[425]);
  assign t[338] = (t[426] & ~t[427]);
  assign t[339] = (t[428] & ~t[429]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = t[430] ^ x[2];
  assign t[341] = t[431] ^ x[1];
  assign t[342] = t[432] ^ x[10];
  assign t[343] = t[433] ^ x[9];
  assign t[344] = t[434] ^ x[13];
  assign t[345] = t[435] ^ x[12];
  assign t[346] = t[436] ^ x[16];
  assign t[347] = t[437] ^ x[15];
  assign t[348] = t[438] ^ x[19];
  assign t[349] = t[439] ^ x[18];
  assign t[34] = ~(t[210] | t[56]);
  assign t[350] = t[440] ^ x[22];
  assign t[351] = t[441] ^ x[21];
  assign t[352] = t[442] ^ x[25];
  assign t[353] = t[443] ^ x[24];
  assign t[354] = t[444] ^ x[28];
  assign t[355] = t[445] ^ x[27];
  assign t[356] = t[446] ^ x[31];
  assign t[357] = t[447] ^ x[30];
  assign t[358] = t[448] ^ x[34];
  assign t[359] = t[449] ^ x[33];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[39];
  assign t[361] = t[451] ^ x[38];
  assign t[362] = t[452] ^ x[42];
  assign t[363] = t[453] ^ x[41];
  assign t[364] = t[454] ^ x[45];
  assign t[365] = t[455] ^ x[44];
  assign t[366] = t[456] ^ x[48];
  assign t[367] = t[457] ^ x[47];
  assign t[368] = t[458] ^ x[51];
  assign t[369] = t[459] ^ x[50];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[56];
  assign t[371] = t[461] ^ x[55];
  assign t[372] = t[462] ^ x[59];
  assign t[373] = t[463] ^ x[58];
  assign t[374] = t[464] ^ x[62];
  assign t[375] = t[465] ^ x[61];
  assign t[376] = t[466] ^ x[65];
  assign t[377] = t[467] ^ x[64];
  assign t[378] = t[468] ^ x[68];
  assign t[379] = t[469] ^ x[67];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[71];
  assign t[381] = t[471] ^ x[70];
  assign t[382] = t[472] ^ x[74];
  assign t[383] = t[473] ^ x[73];
  assign t[384] = t[474] ^ x[79];
  assign t[385] = t[475] ^ x[78];
  assign t[386] = t[476] ^ x[82];
  assign t[387] = t[477] ^ x[81];
  assign t[388] = t[478] ^ x[85];
  assign t[389] = t[479] ^ x[84];
  assign t[38] = ~(t[39] ^ t[63]);
  assign t[390] = t[480] ^ x[90];
  assign t[391] = t[481] ^ x[89];
  assign t[392] = t[482] ^ x[93];
  assign t[393] = t[483] ^ x[92];
  assign t[394] = t[484] ^ x[96];
  assign t[395] = t[485] ^ x[95];
  assign t[396] = t[486] ^ x[99];
  assign t[397] = t[487] ^ x[98];
  assign t[398] = t[488] ^ x[102];
  assign t[399] = t[489] ^ x[101];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[105];
  assign t[401] = t[491] ^ x[104];
  assign t[402] = t[492] ^ x[110];
  assign t[403] = t[493] ^ x[109];
  assign t[404] = t[494] ^ x[113];
  assign t[405] = t[495] ^ x[112];
  assign t[406] = t[496] ^ x[118];
  assign t[407] = t[497] ^ x[117];
  assign t[408] = t[498] ^ x[121];
  assign t[409] = t[499] ^ x[120];
  assign t[40] = ~(t[66] ^ t[67]);
  assign t[410] = t[500] ^ x[124];
  assign t[411] = t[501] ^ x[123];
  assign t[412] = t[502] ^ x[127];
  assign t[413] = t[503] ^ x[126];
  assign t[414] = t[504] ^ x[130];
  assign t[415] = t[505] ^ x[129];
  assign t[416] = t[506] ^ x[133];
  assign t[417] = t[507] ^ x[132];
  assign t[418] = t[508] ^ x[136];
  assign t[419] = t[509] ^ x[135];
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = t[510] ^ x[139];
  assign t[421] = t[511] ^ x[138];
  assign t[422] = t[512] ^ x[142];
  assign t[423] = t[513] ^ x[141];
  assign t[424] = t[514] ^ x[145];
  assign t[425] = t[515] ^ x[144];
  assign t[426] = t[516] ^ x[148];
  assign t[427] = t[517] ^ x[147];
  assign t[428] = t[518] ^ x[151];
  assign t[429] = t[519] ^ x[150];
  assign t[42] = ~(t[211] | t[70]);
  assign t[430] = (x[0]);
  assign t[431] = (x[0]);
  assign t[432] = (x[8]);
  assign t[433] = (x[8]);
  assign t[434] = (x[11]);
  assign t[435] = (x[11]);
  assign t[436] = (x[14]);
  assign t[437] = (x[14]);
  assign t[438] = (x[17]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[20]);
  assign t[441] = (x[20]);
  assign t[442] = (x[23]);
  assign t[443] = (x[23]);
  assign t[444] = (x[26]);
  assign t[445] = (x[26]);
  assign t[446] = (x[29]);
  assign t[447] = (x[29]);
  assign t[448] = (x[32]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[37]);
  assign t[451] = (x[37]);
  assign t[452] = (x[40]);
  assign t[453] = (x[40]);
  assign t[454] = (x[43]);
  assign t[455] = (x[43]);
  assign t[456] = (x[46]);
  assign t[457] = (x[46]);
  assign t[458] = (x[49]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = (x[54]);
  assign t[461] = (x[54]);
  assign t[462] = (x[57]);
  assign t[463] = (x[57]);
  assign t[464] = (x[60]);
  assign t[465] = (x[60]);
  assign t[466] = (x[63]);
  assign t[467] = (x[63]);
  assign t[468] = (x[66]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[77] ^ t[78]);
  assign t[470] = (x[69]);
  assign t[471] = (x[69]);
  assign t[472] = (x[72]);
  assign t[473] = (x[72]);
  assign t[474] = (x[77]);
  assign t[475] = (x[77]);
  assign t[476] = (x[80]);
  assign t[477] = (x[80]);
  assign t[478] = (x[83]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[79] | t[80]);
  assign t[480] = (x[88]);
  assign t[481] = (x[88]);
  assign t[482] = (x[91]);
  assign t[483] = (x[91]);
  assign t[484] = (x[94]);
  assign t[485] = (x[94]);
  assign t[486] = (x[97]);
  assign t[487] = (x[97]);
  assign t[488] = (x[100]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[45] ^ t[81]);
  assign t[490] = (x[103]);
  assign t[491] = (x[103]);
  assign t[492] = (x[108]);
  assign t[493] = (x[108]);
  assign t[494] = (x[111]);
  assign t[495] = (x[111]);
  assign t[496] = (x[116]);
  assign t[497] = (x[116]);
  assign t[498] = (x[119]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[208]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[122]);
  assign t[501] = (x[122]);
  assign t[502] = (x[125]);
  assign t[503] = (x[125]);
  assign t[504] = (x[128]);
  assign t[505] = (x[128]);
  assign t[506] = (x[131]);
  assign t[507] = (x[131]);
  assign t[508] = (x[134]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (x[137]);
  assign t[511] = (x[137]);
  assign t[512] = (x[140]);
  assign t[513] = (x[140]);
  assign t[514] = (x[143]);
  assign t[515] = (x[143]);
  assign t[516] = (x[146]);
  assign t[517] = (x[146]);
  assign t[518] = (x[149]);
  assign t[519] = (x[149]);
  assign t[51] = ~(t[84] & t[85]);
  assign t[52] = ~(t[86] | t[87]);
  assign t[53] = ~(t[86] | t[88]);
  assign t[54] = ~(t[212]);
  assign t[55] = ~(t[213]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[214] | t[93]);
  assign t[59] = t[30] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[215] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[216] | t[103]);
  assign t[66] = ~(t[104] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[217]);
  assign t[69] = ~(t[218]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[219] | t[112]);
  assign t[73] = t[30] ? x[53] : x[52];
  assign t[74] = ~(t[82] & t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[220] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[221] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[126] | t[127]);
  assign t[83] = ~(t[128] & t[129]);
  assign t[84] = ~(t[130] & t[131]);
  assign t[85] = t[128] | t[132];
  assign t[86] = ~(t[128]);
  assign t[87] = t[206] ? t[134] : t[133];
  assign t[88] = t[206] ? t[136] : t[135];
  assign t[89] = ~(t[222]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[212] | t[213]);
  assign t[91] = ~(t[223]);
  assign t[92] = ~(t[224]);
  assign t[93] = ~(t[137] | t[138]);
  assign t[94] = ~(t[52] | t[50]);
  assign t[95] = ~(t[139] & t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = t[143] ? x[76] : x[75];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [151:0] x;
 output y;

 wire [519:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = t[144] | t[145];
  assign t[101] = ~(t[227]);
  assign t[102] = ~(t[228]);
  assign t[103] = ~(t[146] | t[147]);
  assign t[104] = ~(t[148] | t[149]);
  assign t[105] = ~(t[229] | t[150]);
  assign t[106] = t[143] ? x[87] : x[86];
  assign t[107] = ~(t[151] & t[152]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[155] | t[156]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[159] | t[160]);
  assign t[118] = ~(t[235] | t[161]);
  assign t[119] = t[30] ? x[107] : x[106];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[162] & t[163]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[164] | t[165]);
  assign t[124] = t[30] ? x[115] : x[114];
  assign t[125] = ~(t[166] & t[167]);
  assign t[126] = ~(t[128] | t[168]);
  assign t[127] = ~(t[86] | t[169]);
  assign t[128] = ~(t[208]);
  assign t[129] = ~(t[170] & t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[173] | t[174];
  assign t[132] = t[206] ? t[170] : t[175];
  assign t[133] = ~(t[173] & t[176]);
  assign t[134] = ~(t[174] & t[209]);
  assign t[135] = ~(t[173] & t[209]);
  assign t[136] = ~(t[174] & t[176]);
  assign t[137] = ~(t[238]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[207] | t[176]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[86] & t[206];
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[49]);
  assign t[144] = ~(t[177] & t[95]);
  assign t[145] = ~(t[86] | t[178]);
  assign t[146] = ~(t[240]);
  assign t[147] = ~(t[227] | t[228]);
  assign t[148] = ~(t[241]);
  assign t[149] = ~(t[242]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[179] | t[180]);
  assign t[151] = ~(t[52]);
  assign t[152] = ~(t[181] | t[145]);
  assign t[153] = ~(t[243]);
  assign t[154] = ~(t[231] | t[232]);
  assign t[155] = ~(t[86] | t[182]);
  assign t[156] = ~(t[32] & t[85]);
  assign t[157] = ~(t[244]);
  assign t[158] = ~(t[233] | t[234]);
  assign t[159] = ~(t[245]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[246]);
  assign t[161] = ~(t[183] | t[184]);
  assign t[162] = ~(t[52] | t[185]);
  assign t[163] = ~(t[100] | t[186]);
  assign t[164] = ~(t[247]);
  assign t[165] = ~(t[236] | t[237]);
  assign t[166] = ~(t[187] | t[155]);
  assign t[167] = ~(t[126] | t[144]);
  assign t[168] = t[206] ? t[133] : t[136];
  assign t[169] = t[206] ? t[175] : t[188];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(x[4] & t[189]);
  assign t[171] = ~(t[209] & t[190]);
  assign t[172] = ~(t[128] | t[206]);
  assign t[173] = ~(x[4] | t[207]);
  assign t[174] = x[4] & t[207];
  assign t[175] = ~(t[190] & t[176]);
  assign t[176] = ~(t[209]);
  assign t[177] = ~(t[191] | t[192]);
  assign t[178] = t[206] ? t[171] : t[170];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[241] | t[242]);
  assign t[181] = ~(t[193]);
  assign t[182] = t[206] ? t[135] : t[136];
  assign t[183] = ~(t[249]);
  assign t[184] = ~(t[245] | t[246]);
  assign t[185] = ~(t[86] | t[194]);
  assign t[186] = ~(t[195] & t[85]);
  assign t[187] = ~(t[86] | t[196]);
  assign t[188] = ~(x[4] & t[139]);
  assign t[189] = ~(t[207] | t[209]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(x[4] | t[197]);
  assign t[191] = ~(t[128] | t[198]);
  assign t[192] = ~(t[128] | t[199]);
  assign t[193] = ~(t[200] | t[53]);
  assign t[194] = t[206] ? t[170] : t[171];
  assign t[195] = ~(t[201] | t[200]);
  assign t[196] = t[206] ? t[133] : t[134];
  assign t[197] = ~(t[207]);
  assign t[198] = t[206] ? t[136] : t[133];
  assign t[199] = t[206] ? t[175] : t[170];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[86] | t[202]);
  assign t[201] = ~(t[203]);
  assign t[202] = t[206] ? t[188] : t[175];
  assign t[203] = ~(t[172] & t[204]);
  assign t[204] = ~(t[171] & t[188]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[2];
  assign t[251] = t[296] ^ x[10];
  assign t[252] = t[297] ^ x[13];
  assign t[253] = t[298] ^ x[16];
  assign t[254] = t[299] ^ x[19];
  assign t[255] = t[300] ^ x[22];
  assign t[256] = t[301] ^ x[25];
  assign t[257] = t[302] ^ x[28];
  assign t[258] = t[303] ^ x[31];
  assign t[259] = t[304] ^ x[34];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[39];
  assign t[261] = t[306] ^ x[42];
  assign t[262] = t[307] ^ x[45];
  assign t[263] = t[308] ^ x[48];
  assign t[264] = t[309] ^ x[51];
  assign t[265] = t[310] ^ x[56];
  assign t[266] = t[311] ^ x[59];
  assign t[267] = t[312] ^ x[62];
  assign t[268] = t[313] ^ x[65];
  assign t[269] = t[314] ^ x[68];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[71];
  assign t[271] = t[316] ^ x[74];
  assign t[272] = t[317] ^ x[79];
  assign t[273] = t[318] ^ x[82];
  assign t[274] = t[319] ^ x[85];
  assign t[275] = t[320] ^ x[90];
  assign t[276] = t[321] ^ x[93];
  assign t[277] = t[322] ^ x[96];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[102];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[105];
  assign t[281] = t[326] ^ x[110];
  assign t[282] = t[327] ^ x[113];
  assign t[283] = t[328] ^ x[118];
  assign t[284] = t[329] ^ x[121];
  assign t[285] = t[330] ^ x[124];
  assign t[286] = t[331] ^ x[127];
  assign t[287] = t[332] ^ x[130];
  assign t[288] = t[333] ^ x[133];
  assign t[289] = t[334] ^ x[136];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[139];
  assign t[291] = t[336] ^ x[142];
  assign t[292] = t[337] ^ x[145];
  assign t[293] = t[338] ^ x[148];
  assign t[294] = t[339] ^ x[151];
  assign t[295] = (t[340] & ~t[341]);
  assign t[296] = (t[342] & ~t[343]);
  assign t[297] = (t[344] & ~t[345]);
  assign t[298] = (t[346] & ~t[347]);
  assign t[299] = (t[348] & ~t[349]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[350] & ~t[351]);
  assign t[301] = (t[352] & ~t[353]);
  assign t[302] = (t[354] & ~t[355]);
  assign t[303] = (t[356] & ~t[357]);
  assign t[304] = (t[358] & ~t[359]);
  assign t[305] = (t[360] & ~t[361]);
  assign t[306] = (t[362] & ~t[363]);
  assign t[307] = (t[364] & ~t[365]);
  assign t[308] = (t[366] & ~t[367]);
  assign t[309] = (t[368] & ~t[369]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[370] & ~t[371]);
  assign t[311] = (t[372] & ~t[373]);
  assign t[312] = (t[374] & ~t[375]);
  assign t[313] = (t[376] & ~t[377]);
  assign t[314] = (t[378] & ~t[379]);
  assign t[315] = (t[380] & ~t[381]);
  assign t[316] = (t[382] & ~t[383]);
  assign t[317] = (t[384] & ~t[385]);
  assign t[318] = (t[386] & ~t[387]);
  assign t[319] = (t[388] & ~t[389]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[390] & ~t[391]);
  assign t[321] = (t[392] & ~t[393]);
  assign t[322] = (t[394] & ~t[395]);
  assign t[323] = (t[396] & ~t[397]);
  assign t[324] = (t[398] & ~t[399]);
  assign t[325] = (t[400] & ~t[401]);
  assign t[326] = (t[402] & ~t[403]);
  assign t[327] = (t[404] & ~t[405]);
  assign t[328] = (t[406] & ~t[407]);
  assign t[329] = (t[408] & ~t[409]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[410] & ~t[411]);
  assign t[331] = (t[412] & ~t[413]);
  assign t[332] = (t[414] & ~t[415]);
  assign t[333] = (t[416] & ~t[417]);
  assign t[334] = (t[418] & ~t[419]);
  assign t[335] = (t[420] & ~t[421]);
  assign t[336] = (t[422] & ~t[423]);
  assign t[337] = (t[424] & ~t[425]);
  assign t[338] = (t[426] & ~t[427]);
  assign t[339] = (t[428] & ~t[429]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = t[430] ^ x[2];
  assign t[341] = t[431] ^ x[1];
  assign t[342] = t[432] ^ x[10];
  assign t[343] = t[433] ^ x[9];
  assign t[344] = t[434] ^ x[13];
  assign t[345] = t[435] ^ x[12];
  assign t[346] = t[436] ^ x[16];
  assign t[347] = t[437] ^ x[15];
  assign t[348] = t[438] ^ x[19];
  assign t[349] = t[439] ^ x[18];
  assign t[34] = ~(t[210] | t[56]);
  assign t[350] = t[440] ^ x[22];
  assign t[351] = t[441] ^ x[21];
  assign t[352] = t[442] ^ x[25];
  assign t[353] = t[443] ^ x[24];
  assign t[354] = t[444] ^ x[28];
  assign t[355] = t[445] ^ x[27];
  assign t[356] = t[446] ^ x[31];
  assign t[357] = t[447] ^ x[30];
  assign t[358] = t[448] ^ x[34];
  assign t[359] = t[449] ^ x[33];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[39];
  assign t[361] = t[451] ^ x[38];
  assign t[362] = t[452] ^ x[42];
  assign t[363] = t[453] ^ x[41];
  assign t[364] = t[454] ^ x[45];
  assign t[365] = t[455] ^ x[44];
  assign t[366] = t[456] ^ x[48];
  assign t[367] = t[457] ^ x[47];
  assign t[368] = t[458] ^ x[51];
  assign t[369] = t[459] ^ x[50];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[56];
  assign t[371] = t[461] ^ x[55];
  assign t[372] = t[462] ^ x[59];
  assign t[373] = t[463] ^ x[58];
  assign t[374] = t[464] ^ x[62];
  assign t[375] = t[465] ^ x[61];
  assign t[376] = t[466] ^ x[65];
  assign t[377] = t[467] ^ x[64];
  assign t[378] = t[468] ^ x[68];
  assign t[379] = t[469] ^ x[67];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[71];
  assign t[381] = t[471] ^ x[70];
  assign t[382] = t[472] ^ x[74];
  assign t[383] = t[473] ^ x[73];
  assign t[384] = t[474] ^ x[79];
  assign t[385] = t[475] ^ x[78];
  assign t[386] = t[476] ^ x[82];
  assign t[387] = t[477] ^ x[81];
  assign t[388] = t[478] ^ x[85];
  assign t[389] = t[479] ^ x[84];
  assign t[38] = ~(t[39] ^ t[63]);
  assign t[390] = t[480] ^ x[90];
  assign t[391] = t[481] ^ x[89];
  assign t[392] = t[482] ^ x[93];
  assign t[393] = t[483] ^ x[92];
  assign t[394] = t[484] ^ x[96];
  assign t[395] = t[485] ^ x[95];
  assign t[396] = t[486] ^ x[99];
  assign t[397] = t[487] ^ x[98];
  assign t[398] = t[488] ^ x[102];
  assign t[399] = t[489] ^ x[101];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[105];
  assign t[401] = t[491] ^ x[104];
  assign t[402] = t[492] ^ x[110];
  assign t[403] = t[493] ^ x[109];
  assign t[404] = t[494] ^ x[113];
  assign t[405] = t[495] ^ x[112];
  assign t[406] = t[496] ^ x[118];
  assign t[407] = t[497] ^ x[117];
  assign t[408] = t[498] ^ x[121];
  assign t[409] = t[499] ^ x[120];
  assign t[40] = ~(t[66] ^ t[67]);
  assign t[410] = t[500] ^ x[124];
  assign t[411] = t[501] ^ x[123];
  assign t[412] = t[502] ^ x[127];
  assign t[413] = t[503] ^ x[126];
  assign t[414] = t[504] ^ x[130];
  assign t[415] = t[505] ^ x[129];
  assign t[416] = t[506] ^ x[133];
  assign t[417] = t[507] ^ x[132];
  assign t[418] = t[508] ^ x[136];
  assign t[419] = t[509] ^ x[135];
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = t[510] ^ x[139];
  assign t[421] = t[511] ^ x[138];
  assign t[422] = t[512] ^ x[142];
  assign t[423] = t[513] ^ x[141];
  assign t[424] = t[514] ^ x[145];
  assign t[425] = t[515] ^ x[144];
  assign t[426] = t[516] ^ x[148];
  assign t[427] = t[517] ^ x[147];
  assign t[428] = t[518] ^ x[151];
  assign t[429] = t[519] ^ x[150];
  assign t[42] = ~(t[211] | t[70]);
  assign t[430] = (x[0]);
  assign t[431] = (x[0]);
  assign t[432] = (x[8]);
  assign t[433] = (x[8]);
  assign t[434] = (x[11]);
  assign t[435] = (x[11]);
  assign t[436] = (x[14]);
  assign t[437] = (x[14]);
  assign t[438] = (x[17]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[20]);
  assign t[441] = (x[20]);
  assign t[442] = (x[23]);
  assign t[443] = (x[23]);
  assign t[444] = (x[26]);
  assign t[445] = (x[26]);
  assign t[446] = (x[29]);
  assign t[447] = (x[29]);
  assign t[448] = (x[32]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[37]);
  assign t[451] = (x[37]);
  assign t[452] = (x[40]);
  assign t[453] = (x[40]);
  assign t[454] = (x[43]);
  assign t[455] = (x[43]);
  assign t[456] = (x[46]);
  assign t[457] = (x[46]);
  assign t[458] = (x[49]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = (x[54]);
  assign t[461] = (x[54]);
  assign t[462] = (x[57]);
  assign t[463] = (x[57]);
  assign t[464] = (x[60]);
  assign t[465] = (x[60]);
  assign t[466] = (x[63]);
  assign t[467] = (x[63]);
  assign t[468] = (x[66]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[77] ^ t[78]);
  assign t[470] = (x[69]);
  assign t[471] = (x[69]);
  assign t[472] = (x[72]);
  assign t[473] = (x[72]);
  assign t[474] = (x[77]);
  assign t[475] = (x[77]);
  assign t[476] = (x[80]);
  assign t[477] = (x[80]);
  assign t[478] = (x[83]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[79] | t[80]);
  assign t[480] = (x[88]);
  assign t[481] = (x[88]);
  assign t[482] = (x[91]);
  assign t[483] = (x[91]);
  assign t[484] = (x[94]);
  assign t[485] = (x[94]);
  assign t[486] = (x[97]);
  assign t[487] = (x[97]);
  assign t[488] = (x[100]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[45] ^ t[81]);
  assign t[490] = (x[103]);
  assign t[491] = (x[103]);
  assign t[492] = (x[108]);
  assign t[493] = (x[108]);
  assign t[494] = (x[111]);
  assign t[495] = (x[111]);
  assign t[496] = (x[116]);
  assign t[497] = (x[116]);
  assign t[498] = (x[119]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[208]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[122]);
  assign t[501] = (x[122]);
  assign t[502] = (x[125]);
  assign t[503] = (x[125]);
  assign t[504] = (x[128]);
  assign t[505] = (x[128]);
  assign t[506] = (x[131]);
  assign t[507] = (x[131]);
  assign t[508] = (x[134]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (x[137]);
  assign t[511] = (x[137]);
  assign t[512] = (x[140]);
  assign t[513] = (x[140]);
  assign t[514] = (x[143]);
  assign t[515] = (x[143]);
  assign t[516] = (x[146]);
  assign t[517] = (x[146]);
  assign t[518] = (x[149]);
  assign t[519] = (x[149]);
  assign t[51] = ~(t[84] & t[85]);
  assign t[52] = ~(t[86] | t[87]);
  assign t[53] = ~(t[86] | t[88]);
  assign t[54] = ~(t[212]);
  assign t[55] = ~(t[213]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[214] | t[93]);
  assign t[59] = t[30] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[215] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[216] | t[103]);
  assign t[66] = ~(t[104] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[217]);
  assign t[69] = ~(t[218]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[219] | t[112]);
  assign t[73] = t[30] ? x[53] : x[52];
  assign t[74] = ~(t[82] & t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[220] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[221] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[126] | t[127]);
  assign t[83] = ~(t[128] & t[129]);
  assign t[84] = ~(t[130] & t[131]);
  assign t[85] = t[128] | t[132];
  assign t[86] = ~(t[128]);
  assign t[87] = t[206] ? t[134] : t[133];
  assign t[88] = t[206] ? t[136] : t[135];
  assign t[89] = ~(t[222]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[212] | t[213]);
  assign t[91] = ~(t[223]);
  assign t[92] = ~(t[224]);
  assign t[93] = ~(t[137] | t[138]);
  assign t[94] = ~(t[52] | t[50]);
  assign t[95] = ~(t[139] & t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = t[143] ? x[76] : x[75];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[34];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[48] ? x[35] : x[34];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[44];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[68];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[74] ? x[52] : x[51];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[74] ? x[60] : x[59];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[74] ? x[77] : x[76];
  assign t[65] = ~(t[121] & t[84]);
  assign t[66] = ~(t[122] & t[85]);
  assign t[67] = t[48] ? x[85] : x[84];
  assign t[68] = ~(t[86] & t[87]);
  assign t[69] = ~(t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[123]);
  assign t[71] = ~(t[123] & t[88]);
  assign t[72] = ~(t[124]);
  assign t[73] = ~(t[124] & t[89]);
  assign t[74] = ~(t[25]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[34];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[48] ? x[35] : x[34];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[44];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[68];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[74] ? x[52] : x[51];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[74] ? x[60] : x[59];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[74] ? x[77] : x[76];
  assign t[65] = ~(t[121] & t[84]);
  assign t[66] = ~(t[122] & t[85]);
  assign t[67] = t[48] ? x[85] : x[84];
  assign t[68] = ~(t[86] & t[87]);
  assign t[69] = ~(t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[123]);
  assign t[71] = ~(t[123] & t[88]);
  assign t[72] = ~(t[124]);
  assign t[73] = ~(t[124] & t[89]);
  assign t[74] = ~(t[25]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind176(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[155]);
  assign t[104] = ~(t[156]);
  assign t[105] = ~(t[115] & t[116]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[160]);
  assign t[112] = ~(t[117] & t[118]);
  assign t[113] = ~(t[151] & t[150]);
  assign t[114] = ~(t[161]);
  assign t[115] = ~(t[156] & t[155]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[160] & t[159]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[60] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[61] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[129]);
  assign t[53] = t[61] ? x[43] : x[42];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = ~(t[81] & t[130]);
  assign t[56] = t[61] ? x[48] : x[47];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[18] ? x[62] : x[61];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[95]);
  assign t[69] = ~(t[96] & t[135]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[122] ? x[67] : x[66];
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[141]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[142]);
  assign t[81] = ~(t[101] & t[102]);
  assign t[82] = ~(t[103] & t[104]);
  assign t[83] = ~(t[105] & t[143]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[110] & t[111]);
  assign t[93] = ~(t[112] & t[149]);
  assign t[94] = ~(t[150]);
  assign t[95] = ~(t[151]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[155]);
  assign t[104] = ~(t[156]);
  assign t[105] = ~(t[115] & t[116]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[160]);
  assign t[112] = ~(t[117] & t[118]);
  assign t[113] = ~(t[151] & t[150]);
  assign t[114] = ~(t[161]);
  assign t[115] = ~(t[156] & t[155]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[160] & t[159]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[60] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[61] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[129]);
  assign t[53] = t[61] ? x[43] : x[42];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = ~(t[81] & t[130]);
  assign t[56] = t[61] ? x[48] : x[47];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[18] ? x[62] : x[61];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[95]);
  assign t[69] = ~(t[96] & t[135]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[122] ? x[67] : x[66];
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[141]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[142]);
  assign t[81] = ~(t[101] & t[102]);
  assign t[82] = ~(t[103] & t[104]);
  assign t[83] = ~(t[105] & t[143]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[110] & t[111]);
  assign t[93] = ~(t[112] & t[149]);
  assign t[94] = ~(t[150]);
  assign t[95] = ~(t[151]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[108] | t[99]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[109] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[61] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[74] | t[119];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[120];
  assign t[53] = t[78] ? x[43] : x[42];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = t[81] | t[121];
  assign t[56] = t[78] ? x[48] : x[47];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[84] | t[58]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[124];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = t[90] | t[125];
  assign t[66] = t[18] ? x[62] : x[61];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = t[95] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[18] ? x[67] : x[66];
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[132]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[98] | t[79]);
  assign t[82] = ~(t[99] & t[100]);
  assign t[83] = t[101] | t[134];
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[104] & t[105]);
  assign t[92] = t[106] | t[140];
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[107] | t[93]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[108] | t[99]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[109] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[61] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[74] | t[119];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[120];
  assign t[53] = t[78] ? x[43] : x[42];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = t[81] | t[121];
  assign t[56] = t[78] ? x[48] : x[47];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[84] | t[58]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[124];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = t[90] | t[125];
  assign t[66] = t[18] ? x[62] : x[61];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = t[95] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[18] ? x[67] : x[66];
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[132]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[98] | t[79]);
  assign t[82] = ~(t[99] & t[100]);
  assign t[83] = t[101] | t[134];
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[104] & t[105]);
  assign t[92] = t[106] | t[140];
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[107] | t[93]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [139:0] x;
 output y;

 wire [491:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[139] | t[140]);
  assign t[101] = t[141] ? x[78] : x[77];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = ~(t[227]);
  assign t[104] = ~(t[216] | t[217]);
  assign t[105] = ~(t[228]);
  assign t[106] = ~(t[229]);
  assign t[107] = ~(t[144] | t[145]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[232] | t[152]);
  assign t[114] = t[30] ? x[98] : x[97];
  assign t[115] = ~(t[153] & t[154]);
  assign t[116] = ~(t[233]);
  assign t[117] = ~(t[234]);
  assign t[118] = ~(t[155] | t[156]);
  assign t[119] = t[30] ? x[106] : x[105];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[160]);
  assign t[122] = ~(t[161] & t[160]);
  assign t[123] = ~(x[4] & t[162]);
  assign t[124] = ~(t[163] & t[160]);
  assign t[125] = ~(t[161] & t[209]);
  assign t[126] = ~(t[81] | t[164]);
  assign t[127] = ~(t[81] | t[165]);
  assign t[128] = t[206] ? t[166] : t[124];
  assign t[129] = ~(t[79] | t[167]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[168]);
  assign t[131] = ~(t[81] | t[169]);
  assign t[132] = ~(t[235]);
  assign t[133] = ~(t[222] | t[223]);
  assign t[134] = ~(t[236]);
  assign t[135] = ~(t[237]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[127]);
  assign t[138] = ~(t[173] | t[174]);
  assign t[139] = ~(t[238]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[225] | t[226]);
  assign t[141] = ~(t[48]);
  assign t[142] = ~(t[175] | t[176]);
  assign t[143] = ~(t[177]);
  assign t[144] = ~(t[239]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[31] & t[178]);
  assign t[147] = ~(t[179] & t[85]);
  assign t[148] = ~(t[240]);
  assign t[149] = ~(t[230] | t[231]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[241]);
  assign t[151] = ~(t[242]);
  assign t[152] = ~(t[180] | t[181]);
  assign t[153] = ~(t[126] | t[172]);
  assign t[154] = ~(t[182] | t[183]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[233] | t[234]);
  assign t[157] = ~(t[177] | t[51]);
  assign t[158] = ~(t[49] | t[184]);
  assign t[159] = x[4] & t[207];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[209]);
  assign t[161] = ~(x[4] | t[207]);
  assign t[162] = ~(t[207] | t[160]);
  assign t[163] = ~(x[4] | t[185]);
  assign t[164] = t[206] ? t[186] : t[122];
  assign t[165] = t[206] ? t[121] : t[125];
  assign t[166] = ~(x[4] & t[187]);
  assign t[167] = t[206] ? t[124] : t[166];
  assign t[168] = ~(t[175] | t[127]);
  assign t[169] = t[206] ? t[188] : t[166];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(t[244]);
  assign t[171] = ~(t[236] | t[237]);
  assign t[172] = ~(t[81] | t[189]);
  assign t[173] = t[209] & t[190];
  assign t[174] = ~(t[191]);
  assign t[175] = ~(t[81] | t[192]);
  assign t[176] = ~(t[193] & t[191]);
  assign t[177] = ~(t[81] | t[194]);
  assign t[178] = ~(t[79] & t[195]);
  assign t[179] = ~(t[173] & t[196]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[245]);
  assign t[181] = ~(t[241] | t[242]);
  assign t[182] = t[184] | t[131];
  assign t[183] = ~(t[197] & t[85]);
  assign t[184] = ~(t[191] & t[198]);
  assign t[185] = ~(t[207]);
  assign t[186] = ~(t[159] & t[209]);
  assign t[187] = ~(t[207] | t[209]);
  assign t[188] = ~(t[209] & t[163]);
  assign t[189] = t[206] ? t[166] : t[188];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[206]);
  assign t[191] = ~(t[199] | t[129]);
  assign t[192] = t[206] ? t[123] : t[124];
  assign t[193] = ~(t[126] | t[146]);
  assign t[194] = t[206] ? t[122] : t[186];
  assign t[195] = ~(t[166] & t[188]);
  assign t[196] = t[161] | t[159];
  assign t[197] = ~(t[200] | t[175]);
  assign t[198] = ~(t[162] & t[201]);
  assign t[199] = ~(t[79] | t[202]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[203]);
  assign t[201] = t[81] & t[206];
  assign t[202] = t[206] ? t[121] : t[122];
  assign t[203] = ~(t[190] & t[204]);
  assign t[204] = ~(t[188] & t[123]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = (t[283]);
  assign t[243] = (t[284]);
  assign t[244] = (t[285]);
  assign t[245] = (t[286]);
  assign t[246] = t[287] ^ x[2];
  assign t[247] = t[288] ^ x[10];
  assign t[248] = t[289] ^ x[13];
  assign t[249] = t[290] ^ x[16];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[19];
  assign t[251] = t[292] ^ x[22];
  assign t[252] = t[293] ^ x[25];
  assign t[253] = t[294] ^ x[28];
  assign t[254] = t[295] ^ x[31];
  assign t[255] = t[296] ^ x[36];
  assign t[256] = t[297] ^ x[39];
  assign t[257] = t[298] ^ x[42];
  assign t[258] = t[299] ^ x[45];
  assign t[259] = t[300] ^ x[48];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[53];
  assign t[261] = t[302] ^ x[56];
  assign t[262] = t[303] ^ x[59];
  assign t[263] = t[304] ^ x[62];
  assign t[264] = t[305] ^ x[65];
  assign t[265] = t[306] ^ x[68];
  assign t[266] = t[307] ^ x[73];
  assign t[267] = t[308] ^ x[76];
  assign t[268] = t[309] ^ x[81];
  assign t[269] = t[310] ^ x[84];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[87];
  assign t[271] = t[312] ^ x[90];
  assign t[272] = t[313] ^ x[93];
  assign t[273] = t[314] ^ x[96];
  assign t[274] = t[315] ^ x[101];
  assign t[275] = t[316] ^ x[104];
  assign t[276] = t[317] ^ x[109];
  assign t[277] = t[318] ^ x[112];
  assign t[278] = t[319] ^ x[115];
  assign t[279] = t[320] ^ x[118];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[121];
  assign t[281] = t[322] ^ x[124];
  assign t[282] = t[323] ^ x[127];
  assign t[283] = t[324] ^ x[130];
  assign t[284] = t[325] ^ x[133];
  assign t[285] = t[326] ^ x[136];
  assign t[286] = t[327] ^ x[139];
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[354] & ~t[355]);
  assign t[301] = (t[356] & ~t[357]);
  assign t[302] = (t[358] & ~t[359]);
  assign t[303] = (t[360] & ~t[361]);
  assign t[304] = (t[362] & ~t[363]);
  assign t[305] = (t[364] & ~t[365]);
  assign t[306] = (t[366] & ~t[367]);
  assign t[307] = (t[368] & ~t[369]);
  assign t[308] = (t[370] & ~t[371]);
  assign t[309] = (t[372] & ~t[373]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[374] & ~t[375]);
  assign t[311] = (t[376] & ~t[377]);
  assign t[312] = (t[378] & ~t[379]);
  assign t[313] = (t[380] & ~t[381]);
  assign t[314] = (t[382] & ~t[383]);
  assign t[315] = (t[384] & ~t[385]);
  assign t[316] = (t[386] & ~t[387]);
  assign t[317] = (t[388] & ~t[389]);
  assign t[318] = (t[390] & ~t[391]);
  assign t[319] = (t[392] & ~t[393]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[394] & ~t[395]);
  assign t[321] = (t[396] & ~t[397]);
  assign t[322] = (t[398] & ~t[399]);
  assign t[323] = (t[400] & ~t[401]);
  assign t[324] = (t[402] & ~t[403]);
  assign t[325] = (t[404] & ~t[405]);
  assign t[326] = (t[406] & ~t[407]);
  assign t[327] = (t[408] & ~t[409]);
  assign t[328] = t[410] ^ x[2];
  assign t[329] = t[411] ^ x[1];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[10];
  assign t[331] = t[413] ^ x[9];
  assign t[332] = t[414] ^ x[13];
  assign t[333] = t[415] ^ x[12];
  assign t[334] = t[416] ^ x[16];
  assign t[335] = t[417] ^ x[15];
  assign t[336] = t[418] ^ x[19];
  assign t[337] = t[419] ^ x[18];
  assign t[338] = t[420] ^ x[22];
  assign t[339] = t[421] ^ x[21];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[25];
  assign t[341] = t[423] ^ x[24];
  assign t[342] = t[424] ^ x[28];
  assign t[343] = t[425] ^ x[27];
  assign t[344] = t[426] ^ x[31];
  assign t[345] = t[427] ^ x[30];
  assign t[346] = t[428] ^ x[36];
  assign t[347] = t[429] ^ x[35];
  assign t[348] = t[430] ^ x[39];
  assign t[349] = t[431] ^ x[38];
  assign t[34] = ~(t[210] | t[55]);
  assign t[350] = t[432] ^ x[42];
  assign t[351] = t[433] ^ x[41];
  assign t[352] = t[434] ^ x[45];
  assign t[353] = t[435] ^ x[44];
  assign t[354] = t[436] ^ x[48];
  assign t[355] = t[437] ^ x[47];
  assign t[356] = t[438] ^ x[53];
  assign t[357] = t[439] ^ x[52];
  assign t[358] = t[440] ^ x[56];
  assign t[359] = t[441] ^ x[55];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[59];
  assign t[361] = t[443] ^ x[58];
  assign t[362] = t[444] ^ x[62];
  assign t[363] = t[445] ^ x[61];
  assign t[364] = t[446] ^ x[65];
  assign t[365] = t[447] ^ x[64];
  assign t[366] = t[448] ^ x[68];
  assign t[367] = t[449] ^ x[67];
  assign t[368] = t[450] ^ x[73];
  assign t[369] = t[451] ^ x[72];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[76];
  assign t[371] = t[453] ^ x[75];
  assign t[372] = t[454] ^ x[81];
  assign t[373] = t[455] ^ x[80];
  assign t[374] = t[456] ^ x[84];
  assign t[375] = t[457] ^ x[83];
  assign t[376] = t[458] ^ x[87];
  assign t[377] = t[459] ^ x[86];
  assign t[378] = t[460] ^ x[90];
  assign t[379] = t[461] ^ x[89];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[462] ^ x[93];
  assign t[381] = t[463] ^ x[92];
  assign t[382] = t[464] ^ x[96];
  assign t[383] = t[465] ^ x[95];
  assign t[384] = t[466] ^ x[101];
  assign t[385] = t[467] ^ x[100];
  assign t[386] = t[468] ^ x[104];
  assign t[387] = t[469] ^ x[103];
  assign t[388] = t[470] ^ x[109];
  assign t[389] = t[471] ^ x[108];
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = t[472] ^ x[112];
  assign t[391] = t[473] ^ x[111];
  assign t[392] = t[474] ^ x[115];
  assign t[393] = t[475] ^ x[114];
  assign t[394] = t[476] ^ x[118];
  assign t[395] = t[477] ^ x[117];
  assign t[396] = t[478] ^ x[121];
  assign t[397] = t[479] ^ x[120];
  assign t[398] = t[480] ^ x[124];
  assign t[399] = t[481] ^ x[123];
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[127];
  assign t[401] = t[483] ^ x[126];
  assign t[402] = t[484] ^ x[130];
  assign t[403] = t[485] ^ x[129];
  assign t[404] = t[486] ^ x[133];
  assign t[405] = t[487] ^ x[132];
  assign t[406] = t[488] ^ x[136];
  assign t[407] = t[489] ^ x[135];
  assign t[408] = t[490] ^ x[139];
  assign t[409] = t[491] ^ x[138];
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[0]);
  assign t[411] = (x[0]);
  assign t[412] = (x[8]);
  assign t[413] = (x[8]);
  assign t[414] = (x[11]);
  assign t[415] = (x[11]);
  assign t[416] = (x[14]);
  assign t[417] = (x[14]);
  assign t[418] = (x[17]);
  assign t[419] = (x[17]);
  assign t[41] = ~(t[211] | t[67]);
  assign t[420] = (x[20]);
  assign t[421] = (x[20]);
  assign t[422] = (x[23]);
  assign t[423] = (x[23]);
  assign t[424] = (x[26]);
  assign t[425] = (x[26]);
  assign t[426] = (x[29]);
  assign t[427] = (x[29]);
  assign t[428] = (x[34]);
  assign t[429] = (x[34]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[37]);
  assign t[431] = (x[37]);
  assign t[432] = (x[40]);
  assign t[433] = (x[40]);
  assign t[434] = (x[43]);
  assign t[435] = (x[43]);
  assign t[436] = (x[46]);
  assign t[437] = (x[46]);
  assign t[438] = (x[51]);
  assign t[439] = (x[51]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[54]);
  assign t[441] = (x[54]);
  assign t[442] = (x[57]);
  assign t[443] = (x[57]);
  assign t[444] = (x[60]);
  assign t[445] = (x[60]);
  assign t[446] = (x[63]);
  assign t[447] = (x[63]);
  assign t[448] = (x[66]);
  assign t[449] = (x[66]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[71]);
  assign t[451] = (x[71]);
  assign t[452] = (x[74]);
  assign t[453] = (x[74]);
  assign t[454] = (x[79]);
  assign t[455] = (x[79]);
  assign t[456] = (x[82]);
  assign t[457] = (x[82]);
  assign t[458] = (x[85]);
  assign t[459] = (x[85]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = (x[88]);
  assign t[461] = (x[88]);
  assign t[462] = (x[91]);
  assign t[463] = (x[91]);
  assign t[464] = (x[94]);
  assign t[465] = (x[94]);
  assign t[466] = (x[99]);
  assign t[467] = (x[99]);
  assign t[468] = (x[102]);
  assign t[469] = (x[102]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[470] = (x[107]);
  assign t[471] = (x[107]);
  assign t[472] = (x[110]);
  assign t[473] = (x[110]);
  assign t[474] = (x[113]);
  assign t[475] = (x[113]);
  assign t[476] = (x[116]);
  assign t[477] = (x[116]);
  assign t[478] = (x[119]);
  assign t[479] = (x[119]);
  assign t[47] = ~(t[44] ^ t[78]);
  assign t[480] = (x[122]);
  assign t[481] = (x[122]);
  assign t[482] = (x[125]);
  assign t[483] = (x[125]);
  assign t[484] = (x[128]);
  assign t[485] = (x[128]);
  assign t[486] = (x[131]);
  assign t[487] = (x[131]);
  assign t[488] = (x[134]);
  assign t[489] = (x[134]);
  assign t[48] = ~(t[208]);
  assign t[490] = (x[137]);
  assign t[491] = (x[137]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] | t[82]);
  assign t[51] = ~(t[81] | t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = t[88] ? x[33] : x[32];
  assign t[57] = ~(t[89] & t[90]);
  assign t[58] = ~(t[91] | t[92]);
  assign t[59] = ~(t[214] | t[93]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[215] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[103] | t[104]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[218] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[50] : x[49];
  assign t[71] = ~(t[108] & t[84]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[219] | t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[114] ^ t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[220] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[208]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[206] ? t[122] : t[121];
  assign t[81] = ~(t[79]);
  assign t[82] = t[206] ? t[124] : t[123];
  assign t[83] = t[206] ? t[125] : t[121];
  assign t[84] = ~(t[126] | t[127]);
  assign t[85] = t[79] | t[128];
  assign t[86] = ~(t[221]);
  assign t[87] = ~(t[212] | t[213]);
  assign t[88] = ~(t[48]);
  assign t[89] = ~(t[49] | t[129]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[222]);
  assign t[92] = ~(t[223]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[224] | t[136]);
  assign t[96] = t[88] ? x[70] : x[69];
  assign t[97] = ~(t[137] & t[138]);
  assign t[98] = ~(t[225]);
  assign t[99] = ~(t[226]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind181(x, y);
 input [139:0] x;
 output y;

 wire [491:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[139] | t[140]);
  assign t[101] = t[141] ? x[78] : x[77];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = ~(t[227]);
  assign t[104] = ~(t[216] | t[217]);
  assign t[105] = ~(t[228]);
  assign t[106] = ~(t[229]);
  assign t[107] = ~(t[144] | t[145]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[232] | t[152]);
  assign t[114] = t[30] ? x[98] : x[97];
  assign t[115] = ~(t[153] & t[154]);
  assign t[116] = ~(t[233]);
  assign t[117] = ~(t[234]);
  assign t[118] = ~(t[155] | t[156]);
  assign t[119] = t[30] ? x[106] : x[105];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[160]);
  assign t[122] = ~(t[161] & t[160]);
  assign t[123] = ~(x[4] & t[162]);
  assign t[124] = ~(t[163] & t[160]);
  assign t[125] = ~(t[161] & t[209]);
  assign t[126] = ~(t[81] | t[164]);
  assign t[127] = ~(t[81] | t[165]);
  assign t[128] = t[206] ? t[166] : t[124];
  assign t[129] = ~(t[79] | t[167]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[168]);
  assign t[131] = ~(t[81] | t[169]);
  assign t[132] = ~(t[235]);
  assign t[133] = ~(t[222] | t[223]);
  assign t[134] = ~(t[236]);
  assign t[135] = ~(t[237]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[127]);
  assign t[138] = ~(t[173] | t[174]);
  assign t[139] = ~(t[238]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[225] | t[226]);
  assign t[141] = ~(t[48]);
  assign t[142] = ~(t[175] | t[176]);
  assign t[143] = ~(t[177]);
  assign t[144] = ~(t[239]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[31] & t[178]);
  assign t[147] = ~(t[179] & t[85]);
  assign t[148] = ~(t[240]);
  assign t[149] = ~(t[230] | t[231]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[241]);
  assign t[151] = ~(t[242]);
  assign t[152] = ~(t[180] | t[181]);
  assign t[153] = ~(t[126] | t[172]);
  assign t[154] = ~(t[182] | t[183]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[233] | t[234]);
  assign t[157] = ~(t[177] | t[51]);
  assign t[158] = ~(t[49] | t[184]);
  assign t[159] = x[4] & t[207];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[209]);
  assign t[161] = ~(x[4] | t[207]);
  assign t[162] = ~(t[207] | t[160]);
  assign t[163] = ~(x[4] | t[185]);
  assign t[164] = t[206] ? t[186] : t[122];
  assign t[165] = t[206] ? t[121] : t[125];
  assign t[166] = ~(x[4] & t[187]);
  assign t[167] = t[206] ? t[124] : t[166];
  assign t[168] = ~(t[175] | t[127]);
  assign t[169] = t[206] ? t[188] : t[166];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(t[244]);
  assign t[171] = ~(t[236] | t[237]);
  assign t[172] = ~(t[81] | t[189]);
  assign t[173] = t[209] & t[190];
  assign t[174] = ~(t[191]);
  assign t[175] = ~(t[81] | t[192]);
  assign t[176] = ~(t[193] & t[191]);
  assign t[177] = ~(t[81] | t[194]);
  assign t[178] = ~(t[79] & t[195]);
  assign t[179] = ~(t[173] & t[196]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[245]);
  assign t[181] = ~(t[241] | t[242]);
  assign t[182] = t[184] | t[131];
  assign t[183] = ~(t[197] & t[85]);
  assign t[184] = ~(t[191] & t[198]);
  assign t[185] = ~(t[207]);
  assign t[186] = ~(t[159] & t[209]);
  assign t[187] = ~(t[207] | t[209]);
  assign t[188] = ~(t[209] & t[163]);
  assign t[189] = t[206] ? t[166] : t[188];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[206]);
  assign t[191] = ~(t[199] | t[129]);
  assign t[192] = t[206] ? t[123] : t[124];
  assign t[193] = ~(t[126] | t[146]);
  assign t[194] = t[206] ? t[122] : t[186];
  assign t[195] = ~(t[166] & t[188]);
  assign t[196] = t[161] | t[159];
  assign t[197] = ~(t[200] | t[175]);
  assign t[198] = ~(t[162] & t[201]);
  assign t[199] = ~(t[79] | t[202]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[203]);
  assign t[201] = t[81] & t[206];
  assign t[202] = t[206] ? t[121] : t[122];
  assign t[203] = ~(t[190] & t[204]);
  assign t[204] = ~(t[188] & t[123]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = (t[283]);
  assign t[243] = (t[284]);
  assign t[244] = (t[285]);
  assign t[245] = (t[286]);
  assign t[246] = t[287] ^ x[2];
  assign t[247] = t[288] ^ x[10];
  assign t[248] = t[289] ^ x[13];
  assign t[249] = t[290] ^ x[16];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[19];
  assign t[251] = t[292] ^ x[22];
  assign t[252] = t[293] ^ x[25];
  assign t[253] = t[294] ^ x[28];
  assign t[254] = t[295] ^ x[31];
  assign t[255] = t[296] ^ x[36];
  assign t[256] = t[297] ^ x[39];
  assign t[257] = t[298] ^ x[42];
  assign t[258] = t[299] ^ x[45];
  assign t[259] = t[300] ^ x[48];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[53];
  assign t[261] = t[302] ^ x[56];
  assign t[262] = t[303] ^ x[59];
  assign t[263] = t[304] ^ x[62];
  assign t[264] = t[305] ^ x[65];
  assign t[265] = t[306] ^ x[68];
  assign t[266] = t[307] ^ x[73];
  assign t[267] = t[308] ^ x[76];
  assign t[268] = t[309] ^ x[81];
  assign t[269] = t[310] ^ x[84];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[87];
  assign t[271] = t[312] ^ x[90];
  assign t[272] = t[313] ^ x[93];
  assign t[273] = t[314] ^ x[96];
  assign t[274] = t[315] ^ x[101];
  assign t[275] = t[316] ^ x[104];
  assign t[276] = t[317] ^ x[109];
  assign t[277] = t[318] ^ x[112];
  assign t[278] = t[319] ^ x[115];
  assign t[279] = t[320] ^ x[118];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[121];
  assign t[281] = t[322] ^ x[124];
  assign t[282] = t[323] ^ x[127];
  assign t[283] = t[324] ^ x[130];
  assign t[284] = t[325] ^ x[133];
  assign t[285] = t[326] ^ x[136];
  assign t[286] = t[327] ^ x[139];
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[354] & ~t[355]);
  assign t[301] = (t[356] & ~t[357]);
  assign t[302] = (t[358] & ~t[359]);
  assign t[303] = (t[360] & ~t[361]);
  assign t[304] = (t[362] & ~t[363]);
  assign t[305] = (t[364] & ~t[365]);
  assign t[306] = (t[366] & ~t[367]);
  assign t[307] = (t[368] & ~t[369]);
  assign t[308] = (t[370] & ~t[371]);
  assign t[309] = (t[372] & ~t[373]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[374] & ~t[375]);
  assign t[311] = (t[376] & ~t[377]);
  assign t[312] = (t[378] & ~t[379]);
  assign t[313] = (t[380] & ~t[381]);
  assign t[314] = (t[382] & ~t[383]);
  assign t[315] = (t[384] & ~t[385]);
  assign t[316] = (t[386] & ~t[387]);
  assign t[317] = (t[388] & ~t[389]);
  assign t[318] = (t[390] & ~t[391]);
  assign t[319] = (t[392] & ~t[393]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[394] & ~t[395]);
  assign t[321] = (t[396] & ~t[397]);
  assign t[322] = (t[398] & ~t[399]);
  assign t[323] = (t[400] & ~t[401]);
  assign t[324] = (t[402] & ~t[403]);
  assign t[325] = (t[404] & ~t[405]);
  assign t[326] = (t[406] & ~t[407]);
  assign t[327] = (t[408] & ~t[409]);
  assign t[328] = t[410] ^ x[2];
  assign t[329] = t[411] ^ x[1];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[10];
  assign t[331] = t[413] ^ x[9];
  assign t[332] = t[414] ^ x[13];
  assign t[333] = t[415] ^ x[12];
  assign t[334] = t[416] ^ x[16];
  assign t[335] = t[417] ^ x[15];
  assign t[336] = t[418] ^ x[19];
  assign t[337] = t[419] ^ x[18];
  assign t[338] = t[420] ^ x[22];
  assign t[339] = t[421] ^ x[21];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[25];
  assign t[341] = t[423] ^ x[24];
  assign t[342] = t[424] ^ x[28];
  assign t[343] = t[425] ^ x[27];
  assign t[344] = t[426] ^ x[31];
  assign t[345] = t[427] ^ x[30];
  assign t[346] = t[428] ^ x[36];
  assign t[347] = t[429] ^ x[35];
  assign t[348] = t[430] ^ x[39];
  assign t[349] = t[431] ^ x[38];
  assign t[34] = ~(t[210] | t[55]);
  assign t[350] = t[432] ^ x[42];
  assign t[351] = t[433] ^ x[41];
  assign t[352] = t[434] ^ x[45];
  assign t[353] = t[435] ^ x[44];
  assign t[354] = t[436] ^ x[48];
  assign t[355] = t[437] ^ x[47];
  assign t[356] = t[438] ^ x[53];
  assign t[357] = t[439] ^ x[52];
  assign t[358] = t[440] ^ x[56];
  assign t[359] = t[441] ^ x[55];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[59];
  assign t[361] = t[443] ^ x[58];
  assign t[362] = t[444] ^ x[62];
  assign t[363] = t[445] ^ x[61];
  assign t[364] = t[446] ^ x[65];
  assign t[365] = t[447] ^ x[64];
  assign t[366] = t[448] ^ x[68];
  assign t[367] = t[449] ^ x[67];
  assign t[368] = t[450] ^ x[73];
  assign t[369] = t[451] ^ x[72];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[76];
  assign t[371] = t[453] ^ x[75];
  assign t[372] = t[454] ^ x[81];
  assign t[373] = t[455] ^ x[80];
  assign t[374] = t[456] ^ x[84];
  assign t[375] = t[457] ^ x[83];
  assign t[376] = t[458] ^ x[87];
  assign t[377] = t[459] ^ x[86];
  assign t[378] = t[460] ^ x[90];
  assign t[379] = t[461] ^ x[89];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[462] ^ x[93];
  assign t[381] = t[463] ^ x[92];
  assign t[382] = t[464] ^ x[96];
  assign t[383] = t[465] ^ x[95];
  assign t[384] = t[466] ^ x[101];
  assign t[385] = t[467] ^ x[100];
  assign t[386] = t[468] ^ x[104];
  assign t[387] = t[469] ^ x[103];
  assign t[388] = t[470] ^ x[109];
  assign t[389] = t[471] ^ x[108];
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = t[472] ^ x[112];
  assign t[391] = t[473] ^ x[111];
  assign t[392] = t[474] ^ x[115];
  assign t[393] = t[475] ^ x[114];
  assign t[394] = t[476] ^ x[118];
  assign t[395] = t[477] ^ x[117];
  assign t[396] = t[478] ^ x[121];
  assign t[397] = t[479] ^ x[120];
  assign t[398] = t[480] ^ x[124];
  assign t[399] = t[481] ^ x[123];
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[127];
  assign t[401] = t[483] ^ x[126];
  assign t[402] = t[484] ^ x[130];
  assign t[403] = t[485] ^ x[129];
  assign t[404] = t[486] ^ x[133];
  assign t[405] = t[487] ^ x[132];
  assign t[406] = t[488] ^ x[136];
  assign t[407] = t[489] ^ x[135];
  assign t[408] = t[490] ^ x[139];
  assign t[409] = t[491] ^ x[138];
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[0]);
  assign t[411] = (x[0]);
  assign t[412] = (x[8]);
  assign t[413] = (x[8]);
  assign t[414] = (x[11]);
  assign t[415] = (x[11]);
  assign t[416] = (x[14]);
  assign t[417] = (x[14]);
  assign t[418] = (x[17]);
  assign t[419] = (x[17]);
  assign t[41] = ~(t[211] | t[67]);
  assign t[420] = (x[20]);
  assign t[421] = (x[20]);
  assign t[422] = (x[23]);
  assign t[423] = (x[23]);
  assign t[424] = (x[26]);
  assign t[425] = (x[26]);
  assign t[426] = (x[29]);
  assign t[427] = (x[29]);
  assign t[428] = (x[34]);
  assign t[429] = (x[34]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[37]);
  assign t[431] = (x[37]);
  assign t[432] = (x[40]);
  assign t[433] = (x[40]);
  assign t[434] = (x[43]);
  assign t[435] = (x[43]);
  assign t[436] = (x[46]);
  assign t[437] = (x[46]);
  assign t[438] = (x[51]);
  assign t[439] = (x[51]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[54]);
  assign t[441] = (x[54]);
  assign t[442] = (x[57]);
  assign t[443] = (x[57]);
  assign t[444] = (x[60]);
  assign t[445] = (x[60]);
  assign t[446] = (x[63]);
  assign t[447] = (x[63]);
  assign t[448] = (x[66]);
  assign t[449] = (x[66]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[71]);
  assign t[451] = (x[71]);
  assign t[452] = (x[74]);
  assign t[453] = (x[74]);
  assign t[454] = (x[79]);
  assign t[455] = (x[79]);
  assign t[456] = (x[82]);
  assign t[457] = (x[82]);
  assign t[458] = (x[85]);
  assign t[459] = (x[85]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = (x[88]);
  assign t[461] = (x[88]);
  assign t[462] = (x[91]);
  assign t[463] = (x[91]);
  assign t[464] = (x[94]);
  assign t[465] = (x[94]);
  assign t[466] = (x[99]);
  assign t[467] = (x[99]);
  assign t[468] = (x[102]);
  assign t[469] = (x[102]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[470] = (x[107]);
  assign t[471] = (x[107]);
  assign t[472] = (x[110]);
  assign t[473] = (x[110]);
  assign t[474] = (x[113]);
  assign t[475] = (x[113]);
  assign t[476] = (x[116]);
  assign t[477] = (x[116]);
  assign t[478] = (x[119]);
  assign t[479] = (x[119]);
  assign t[47] = ~(t[44] ^ t[78]);
  assign t[480] = (x[122]);
  assign t[481] = (x[122]);
  assign t[482] = (x[125]);
  assign t[483] = (x[125]);
  assign t[484] = (x[128]);
  assign t[485] = (x[128]);
  assign t[486] = (x[131]);
  assign t[487] = (x[131]);
  assign t[488] = (x[134]);
  assign t[489] = (x[134]);
  assign t[48] = ~(t[208]);
  assign t[490] = (x[137]);
  assign t[491] = (x[137]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] | t[82]);
  assign t[51] = ~(t[81] | t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = t[88] ? x[33] : x[32];
  assign t[57] = ~(t[89] & t[90]);
  assign t[58] = ~(t[91] | t[92]);
  assign t[59] = ~(t[214] | t[93]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[215] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[103] | t[104]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[218] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[50] : x[49];
  assign t[71] = ~(t[108] & t[84]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[219] | t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[114] ^ t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[220] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[208]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[206] ? t[122] : t[121];
  assign t[81] = ~(t[79]);
  assign t[82] = t[206] ? t[124] : t[123];
  assign t[83] = t[206] ? t[125] : t[121];
  assign t[84] = ~(t[126] | t[127]);
  assign t[85] = t[79] | t[128];
  assign t[86] = ~(t[221]);
  assign t[87] = ~(t[212] | t[213]);
  assign t[88] = ~(t[48]);
  assign t[89] = ~(t[49] | t[129]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[222]);
  assign t[92] = ~(t[223]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[224] | t[136]);
  assign t[96] = t[88] ? x[70] : x[69];
  assign t[97] = ~(t[137] & t[138]);
  assign t[98] = ~(t[225]);
  assign t[99] = ~(t[226]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[49];
  assign t[139] = t[171] ^ x[52];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[57];
  assign t[141] = t[173] ^ x[60];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[49];
  assign t[215] = t[279] ^ x[48];
  assign t[216] = t[280] ^ x[52];
  assign t[217] = t[281] ^ x[51];
  assign t[218] = t[282] ^ x[57];
  assign t[219] = t[283] ^ x[56];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[60];
  assign t[221] = t[285] ^ x[59];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[47]);
  assign t[279] = (x[47]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[50]);
  assign t[282] = (x[55]);
  assign t[283] = (x[55]);
  assign t[284] = (x[58]);
  assign t[285] = (x[58]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[27] : x[26];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[41];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[54];
  assign t[37] = ~(t[101] & t[55]);
  assign t[38] = ~(t[102] & t[56]);
  assign t[39] = t[47] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[43];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[69] ? x[46] : x[45];
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[47] ? x[54] : x[53];
  assign t[54] = ~(t[72] & t[73]);
  assign t[55] = ~(t[108]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = ~(t[109] & t[75]);
  assign t[58] = ~(t[110] & t[76]);
  assign t[59] = ~(t[111] & t[77]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[112] & t[78]);
  assign t[61] = t[69] ? x[71] : x[70];
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[79] : x[78];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[25]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[118] & t[86]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[119]);
  assign t[76] = ~(t[119] & t[87]);
  assign t[77] = ~(t[120]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[124]);
  assign t[86] = ~(t[124] & t[92]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[49];
  assign t[139] = t[171] ^ x[52];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[57];
  assign t[141] = t[173] ^ x[60];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[49];
  assign t[215] = t[279] ^ x[48];
  assign t[216] = t[280] ^ x[52];
  assign t[217] = t[281] ^ x[51];
  assign t[218] = t[282] ^ x[57];
  assign t[219] = t[283] ^ x[56];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[60];
  assign t[221] = t[285] ^ x[59];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[47]);
  assign t[279] = (x[47]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[50]);
  assign t[282] = (x[55]);
  assign t[283] = (x[55]);
  assign t[284] = (x[58]);
  assign t[285] = (x[58]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[27] : x[26];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[41];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[54];
  assign t[37] = ~(t[101] & t[55]);
  assign t[38] = ~(t[102] & t[56]);
  assign t[39] = t[47] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[43];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[69] ? x[46] : x[45];
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[47] ? x[54] : x[53];
  assign t[54] = ~(t[72] & t[73]);
  assign t[55] = ~(t[108]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = ~(t[109] & t[75]);
  assign t[58] = ~(t[110] & t[76]);
  assign t[59] = ~(t[111] & t[77]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[112] & t[78]);
  assign t[61] = t[69] ? x[71] : x[70];
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[79] : x[78];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[25]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[118] & t[86]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[119]);
  assign t[76] = ~(t[119] & t[87]);
  assign t[77] = ~(t[120]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[124]);
  assign t[86] = ~(t[124] & t[92]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [139:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[110] & t[111]);
  assign t[106] = ~(t[141] & t[140]);
  assign t[107] = ~(t[150]);
  assign t[108] = ~(t[145] & t[144]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[149] & t[148]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[2];
  assign t[154] = t[195] ^ x[10];
  assign t[155] = t[196] ^ x[13];
  assign t[156] = t[197] ^ x[16];
  assign t[157] = t[198] ^ x[19];
  assign t[158] = t[199] ^ x[22];
  assign t[159] = t[200] ^ x[27];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[32];
  assign t[161] = t[202] ^ x[35];
  assign t[162] = t[203] ^ x[38];
  assign t[163] = t[204] ^ x[43];
  assign t[164] = t[205] ^ x[48];
  assign t[165] = t[206] ^ x[51];
  assign t[166] = t[207] ^ x[54];
  assign t[167] = t[208] ^ x[57];
  assign t[168] = t[209] ^ x[62];
  assign t[169] = t[210] ^ x[67];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[70];
  assign t[171] = t[212] ^ x[73];
  assign t[172] = t[213] ^ x[76];
  assign t[173] = t[214] ^ x[79];
  assign t[174] = t[215] ^ x[82];
  assign t[175] = t[216] ^ x[85];
  assign t[176] = t[217] ^ x[88];
  assign t[177] = t[218] ^ x[91];
  assign t[178] = t[219] ^ x[94];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[100];
  assign t[181] = t[222] ^ x[103];
  assign t[182] = t[223] ^ x[106];
  assign t[183] = t[224] ^ x[109];
  assign t[184] = t[225] ^ x[112];
  assign t[185] = t[226] ^ x[115];
  assign t[186] = t[227] ^ x[118];
  assign t[187] = t[228] ^ x[121];
  assign t[188] = t[229] ^ x[124];
  assign t[189] = t[230] ^ x[127];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[130];
  assign t[191] = t[232] ^ x[133];
  assign t[192] = t[233] ^ x[136];
  assign t[193] = t[234] ^ x[139];
  assign t[194] = (t[235] & ~t[236]);
  assign t[195] = (t[237] & ~t[238]);
  assign t[196] = (t[239] & ~t[240]);
  assign t[197] = (t[241] & ~t[242]);
  assign t[198] = (t[243] & ~t[244]);
  assign t[199] = (t[245] & ~t[246]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[247] & ~t[248]);
  assign t[201] = (t[249] & ~t[250]);
  assign t[202] = (t[251] & ~t[252]);
  assign t[203] = (t[253] & ~t[254]);
  assign t[204] = (t[255] & ~t[256]);
  assign t[205] = (t[257] & ~t[258]);
  assign t[206] = (t[259] & ~t[260]);
  assign t[207] = (t[261] & ~t[262]);
  assign t[208] = (t[263] & ~t[264]);
  assign t[209] = (t[265] & ~t[266]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[267] & ~t[268]);
  assign t[211] = (t[269] & ~t[270]);
  assign t[212] = (t[271] & ~t[272]);
  assign t[213] = (t[273] & ~t[274]);
  assign t[214] = (t[275] & ~t[276]);
  assign t[215] = (t[277] & ~t[278]);
  assign t[216] = (t[279] & ~t[280]);
  assign t[217] = (t[281] & ~t[282]);
  assign t[218] = (t[283] & ~t[284]);
  assign t[219] = (t[285] & ~t[286]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[287] & ~t[288]);
  assign t[221] = (t[289] & ~t[290]);
  assign t[222] = (t[291] & ~t[292]);
  assign t[223] = (t[293] & ~t[294]);
  assign t[224] = (t[295] & ~t[296]);
  assign t[225] = (t[297] & ~t[298]);
  assign t[226] = (t[299] & ~t[300]);
  assign t[227] = (t[301] & ~t[302]);
  assign t[228] = (t[303] & ~t[304]);
  assign t[229] = (t[305] & ~t[306]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (t[307] & ~t[308]);
  assign t[231] = (t[309] & ~t[310]);
  assign t[232] = (t[311] & ~t[312]);
  assign t[233] = (t[313] & ~t[314]);
  assign t[234] = (t[315] & ~t[316]);
  assign t[235] = t[317] ^ x[2];
  assign t[236] = t[318] ^ x[1];
  assign t[237] = t[319] ^ x[10];
  assign t[238] = t[320] ^ x[9];
  assign t[239] = t[321] ^ x[13];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[12];
  assign t[241] = t[323] ^ x[16];
  assign t[242] = t[324] ^ x[15];
  assign t[243] = t[325] ^ x[19];
  assign t[244] = t[326] ^ x[18];
  assign t[245] = t[327] ^ x[22];
  assign t[246] = t[328] ^ x[21];
  assign t[247] = t[329] ^ x[27];
  assign t[248] = t[330] ^ x[26];
  assign t[249] = t[331] ^ x[32];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[31];
  assign t[251] = t[333] ^ x[35];
  assign t[252] = t[334] ^ x[34];
  assign t[253] = t[335] ^ x[38];
  assign t[254] = t[336] ^ x[37];
  assign t[255] = t[337] ^ x[43];
  assign t[256] = t[338] ^ x[42];
  assign t[257] = t[339] ^ x[48];
  assign t[258] = t[340] ^ x[47];
  assign t[259] = t[341] ^ x[51];
  assign t[25] = ~(t[115]);
  assign t[260] = t[342] ^ x[50];
  assign t[261] = t[343] ^ x[54];
  assign t[262] = t[344] ^ x[53];
  assign t[263] = t[345] ^ x[57];
  assign t[264] = t[346] ^ x[56];
  assign t[265] = t[347] ^ x[62];
  assign t[266] = t[348] ^ x[61];
  assign t[267] = t[349] ^ x[67];
  assign t[268] = t[350] ^ x[66];
  assign t[269] = t[351] ^ x[70];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[69];
  assign t[271] = t[353] ^ x[73];
  assign t[272] = t[354] ^ x[72];
  assign t[273] = t[355] ^ x[76];
  assign t[274] = t[356] ^ x[75];
  assign t[275] = t[357] ^ x[79];
  assign t[276] = t[358] ^ x[78];
  assign t[277] = t[359] ^ x[82];
  assign t[278] = t[360] ^ x[81];
  assign t[279] = t[361] ^ x[85];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[84];
  assign t[281] = t[363] ^ x[88];
  assign t[282] = t[364] ^ x[87];
  assign t[283] = t[365] ^ x[91];
  assign t[284] = t[366] ^ x[90];
  assign t[285] = t[367] ^ x[94];
  assign t[286] = t[368] ^ x[93];
  assign t[287] = t[369] ^ x[97];
  assign t[288] = t[370] ^ x[96];
  assign t[289] = t[371] ^ x[100];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[99];
  assign t[291] = t[373] ^ x[103];
  assign t[292] = t[374] ^ x[102];
  assign t[293] = t[375] ^ x[106];
  assign t[294] = t[376] ^ x[105];
  assign t[295] = t[377] ^ x[109];
  assign t[296] = t[378] ^ x[108];
  assign t[297] = t[379] ^ x[112];
  assign t[298] = t[380] ^ x[111];
  assign t[299] = t[381] ^ x[115];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[114];
  assign t[301] = t[383] ^ x[118];
  assign t[302] = t[384] ^ x[117];
  assign t[303] = t[385] ^ x[121];
  assign t[304] = t[386] ^ x[120];
  assign t[305] = t[387] ^ x[124];
  assign t[306] = t[388] ^ x[123];
  assign t[307] = t[389] ^ x[127];
  assign t[308] = t[390] ^ x[126];
  assign t[309] = t[391] ^ x[130];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[129];
  assign t[311] = t[393] ^ x[133];
  assign t[312] = t[394] ^ x[132];
  assign t[313] = t[395] ^ x[136];
  assign t[314] = t[396] ^ x[135];
  assign t[315] = t[397] ^ x[139];
  assign t[316] = t[398] ^ x[138];
  assign t[317] = (x[0]);
  assign t[318] = (x[0]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[8]);
  assign t[321] = (x[11]);
  assign t[322] = (x[11]);
  assign t[323] = (x[14]);
  assign t[324] = (x[14]);
  assign t[325] = (x[17]);
  assign t[326] = (x[17]);
  assign t[327] = (x[20]);
  assign t[328] = (x[20]);
  assign t[329] = (x[25]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[25]);
  assign t[331] = (x[30]);
  assign t[332] = (x[30]);
  assign t[333] = (x[33]);
  assign t[334] = (x[33]);
  assign t[335] = (x[36]);
  assign t[336] = (x[36]);
  assign t[337] = (x[41]);
  assign t[338] = (x[41]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[46]);
  assign t[341] = (x[49]);
  assign t[342] = (x[49]);
  assign t[343] = (x[52]);
  assign t[344] = (x[52]);
  assign t[345] = (x[55]);
  assign t[346] = (x[55]);
  assign t[347] = (x[60]);
  assign t[348] = (x[60]);
  assign t[349] = (x[65]);
  assign t[34] = t[51] ^ t[43];
  assign t[350] = (x[65]);
  assign t[351] = (x[68]);
  assign t[352] = (x[68]);
  assign t[353] = (x[71]);
  assign t[354] = (x[71]);
  assign t[355] = (x[74]);
  assign t[356] = (x[74]);
  assign t[357] = (x[77]);
  assign t[358] = (x[77]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[80]);
  assign t[361] = (x[83]);
  assign t[362] = (x[83]);
  assign t[363] = (x[86]);
  assign t[364] = (x[86]);
  assign t[365] = (x[89]);
  assign t[366] = (x[89]);
  assign t[367] = (x[92]);
  assign t[368] = (x[92]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[55];
  assign t[370] = (x[95]);
  assign t[371] = (x[98]);
  assign t[372] = (x[98]);
  assign t[373] = (x[101]);
  assign t[374] = (x[101]);
  assign t[375] = (x[104]);
  assign t[376] = (x[104]);
  assign t[377] = (x[107]);
  assign t[378] = (x[107]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[110]);
  assign t[381] = (x[113]);
  assign t[382] = (x[113]);
  assign t[383] = (x[116]);
  assign t[384] = (x[116]);
  assign t[385] = (x[119]);
  assign t[386] = (x[119]);
  assign t[387] = (x[122]);
  assign t[388] = (x[122]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[58] & t[118]);
  assign t[390] = (x[125]);
  assign t[391] = (x[128]);
  assign t[392] = (x[128]);
  assign t[393] = (x[131]);
  assign t[394] = (x[131]);
  assign t[395] = (x[134]);
  assign t[396] = (x[134]);
  assign t[397] = (x[137]);
  assign t[398] = (x[137]);
  assign t[39] = t[59] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[41];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[121]);
  assign t[51] = t[18] ? x[40] : x[39];
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[122]);
  assign t[54] = t[48] ? x[45] : x[44];
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = ~(t[83] & t[125]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[86] & t[126]);
  assign t[64] = t[59] ? x[59] : x[58];
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[91] & t[127]);
  assign t[68] = t[115] ? x[64] : x[63];
  assign t[69] = ~(t[120] & t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[130]);
  assign t[73] = ~(t[92] & t[93]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[94] & t[95]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[98] & t[133]);
  assign t[79] = ~(t[124] & t[123]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[99] & t[100]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[138]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[104]);
  assign t[88] = ~(t[105] & t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[141]);
  assign t[91] = ~(t[106] & t[107]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[145]);
  assign t[98] = ~(t[108] & t[109]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [139:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[110] & t[111]);
  assign t[106] = ~(t[141] & t[140]);
  assign t[107] = ~(t[150]);
  assign t[108] = ~(t[145] & t[144]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[149] & t[148]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[2];
  assign t[154] = t[195] ^ x[10];
  assign t[155] = t[196] ^ x[13];
  assign t[156] = t[197] ^ x[16];
  assign t[157] = t[198] ^ x[19];
  assign t[158] = t[199] ^ x[22];
  assign t[159] = t[200] ^ x[27];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[32];
  assign t[161] = t[202] ^ x[35];
  assign t[162] = t[203] ^ x[38];
  assign t[163] = t[204] ^ x[43];
  assign t[164] = t[205] ^ x[48];
  assign t[165] = t[206] ^ x[51];
  assign t[166] = t[207] ^ x[54];
  assign t[167] = t[208] ^ x[57];
  assign t[168] = t[209] ^ x[62];
  assign t[169] = t[210] ^ x[67];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[70];
  assign t[171] = t[212] ^ x[73];
  assign t[172] = t[213] ^ x[76];
  assign t[173] = t[214] ^ x[79];
  assign t[174] = t[215] ^ x[82];
  assign t[175] = t[216] ^ x[85];
  assign t[176] = t[217] ^ x[88];
  assign t[177] = t[218] ^ x[91];
  assign t[178] = t[219] ^ x[94];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[100];
  assign t[181] = t[222] ^ x[103];
  assign t[182] = t[223] ^ x[106];
  assign t[183] = t[224] ^ x[109];
  assign t[184] = t[225] ^ x[112];
  assign t[185] = t[226] ^ x[115];
  assign t[186] = t[227] ^ x[118];
  assign t[187] = t[228] ^ x[121];
  assign t[188] = t[229] ^ x[124];
  assign t[189] = t[230] ^ x[127];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[130];
  assign t[191] = t[232] ^ x[133];
  assign t[192] = t[233] ^ x[136];
  assign t[193] = t[234] ^ x[139];
  assign t[194] = (t[235] & ~t[236]);
  assign t[195] = (t[237] & ~t[238]);
  assign t[196] = (t[239] & ~t[240]);
  assign t[197] = (t[241] & ~t[242]);
  assign t[198] = (t[243] & ~t[244]);
  assign t[199] = (t[245] & ~t[246]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[247] & ~t[248]);
  assign t[201] = (t[249] & ~t[250]);
  assign t[202] = (t[251] & ~t[252]);
  assign t[203] = (t[253] & ~t[254]);
  assign t[204] = (t[255] & ~t[256]);
  assign t[205] = (t[257] & ~t[258]);
  assign t[206] = (t[259] & ~t[260]);
  assign t[207] = (t[261] & ~t[262]);
  assign t[208] = (t[263] & ~t[264]);
  assign t[209] = (t[265] & ~t[266]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[267] & ~t[268]);
  assign t[211] = (t[269] & ~t[270]);
  assign t[212] = (t[271] & ~t[272]);
  assign t[213] = (t[273] & ~t[274]);
  assign t[214] = (t[275] & ~t[276]);
  assign t[215] = (t[277] & ~t[278]);
  assign t[216] = (t[279] & ~t[280]);
  assign t[217] = (t[281] & ~t[282]);
  assign t[218] = (t[283] & ~t[284]);
  assign t[219] = (t[285] & ~t[286]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[287] & ~t[288]);
  assign t[221] = (t[289] & ~t[290]);
  assign t[222] = (t[291] & ~t[292]);
  assign t[223] = (t[293] & ~t[294]);
  assign t[224] = (t[295] & ~t[296]);
  assign t[225] = (t[297] & ~t[298]);
  assign t[226] = (t[299] & ~t[300]);
  assign t[227] = (t[301] & ~t[302]);
  assign t[228] = (t[303] & ~t[304]);
  assign t[229] = (t[305] & ~t[306]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (t[307] & ~t[308]);
  assign t[231] = (t[309] & ~t[310]);
  assign t[232] = (t[311] & ~t[312]);
  assign t[233] = (t[313] & ~t[314]);
  assign t[234] = (t[315] & ~t[316]);
  assign t[235] = t[317] ^ x[2];
  assign t[236] = t[318] ^ x[1];
  assign t[237] = t[319] ^ x[10];
  assign t[238] = t[320] ^ x[9];
  assign t[239] = t[321] ^ x[13];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[12];
  assign t[241] = t[323] ^ x[16];
  assign t[242] = t[324] ^ x[15];
  assign t[243] = t[325] ^ x[19];
  assign t[244] = t[326] ^ x[18];
  assign t[245] = t[327] ^ x[22];
  assign t[246] = t[328] ^ x[21];
  assign t[247] = t[329] ^ x[27];
  assign t[248] = t[330] ^ x[26];
  assign t[249] = t[331] ^ x[32];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[31];
  assign t[251] = t[333] ^ x[35];
  assign t[252] = t[334] ^ x[34];
  assign t[253] = t[335] ^ x[38];
  assign t[254] = t[336] ^ x[37];
  assign t[255] = t[337] ^ x[43];
  assign t[256] = t[338] ^ x[42];
  assign t[257] = t[339] ^ x[48];
  assign t[258] = t[340] ^ x[47];
  assign t[259] = t[341] ^ x[51];
  assign t[25] = ~(t[115]);
  assign t[260] = t[342] ^ x[50];
  assign t[261] = t[343] ^ x[54];
  assign t[262] = t[344] ^ x[53];
  assign t[263] = t[345] ^ x[57];
  assign t[264] = t[346] ^ x[56];
  assign t[265] = t[347] ^ x[62];
  assign t[266] = t[348] ^ x[61];
  assign t[267] = t[349] ^ x[67];
  assign t[268] = t[350] ^ x[66];
  assign t[269] = t[351] ^ x[70];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[69];
  assign t[271] = t[353] ^ x[73];
  assign t[272] = t[354] ^ x[72];
  assign t[273] = t[355] ^ x[76];
  assign t[274] = t[356] ^ x[75];
  assign t[275] = t[357] ^ x[79];
  assign t[276] = t[358] ^ x[78];
  assign t[277] = t[359] ^ x[82];
  assign t[278] = t[360] ^ x[81];
  assign t[279] = t[361] ^ x[85];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[84];
  assign t[281] = t[363] ^ x[88];
  assign t[282] = t[364] ^ x[87];
  assign t[283] = t[365] ^ x[91];
  assign t[284] = t[366] ^ x[90];
  assign t[285] = t[367] ^ x[94];
  assign t[286] = t[368] ^ x[93];
  assign t[287] = t[369] ^ x[97];
  assign t[288] = t[370] ^ x[96];
  assign t[289] = t[371] ^ x[100];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[99];
  assign t[291] = t[373] ^ x[103];
  assign t[292] = t[374] ^ x[102];
  assign t[293] = t[375] ^ x[106];
  assign t[294] = t[376] ^ x[105];
  assign t[295] = t[377] ^ x[109];
  assign t[296] = t[378] ^ x[108];
  assign t[297] = t[379] ^ x[112];
  assign t[298] = t[380] ^ x[111];
  assign t[299] = t[381] ^ x[115];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[114];
  assign t[301] = t[383] ^ x[118];
  assign t[302] = t[384] ^ x[117];
  assign t[303] = t[385] ^ x[121];
  assign t[304] = t[386] ^ x[120];
  assign t[305] = t[387] ^ x[124];
  assign t[306] = t[388] ^ x[123];
  assign t[307] = t[389] ^ x[127];
  assign t[308] = t[390] ^ x[126];
  assign t[309] = t[391] ^ x[130];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[129];
  assign t[311] = t[393] ^ x[133];
  assign t[312] = t[394] ^ x[132];
  assign t[313] = t[395] ^ x[136];
  assign t[314] = t[396] ^ x[135];
  assign t[315] = t[397] ^ x[139];
  assign t[316] = t[398] ^ x[138];
  assign t[317] = (x[0]);
  assign t[318] = (x[0]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[8]);
  assign t[321] = (x[11]);
  assign t[322] = (x[11]);
  assign t[323] = (x[14]);
  assign t[324] = (x[14]);
  assign t[325] = (x[17]);
  assign t[326] = (x[17]);
  assign t[327] = (x[20]);
  assign t[328] = (x[20]);
  assign t[329] = (x[25]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[25]);
  assign t[331] = (x[30]);
  assign t[332] = (x[30]);
  assign t[333] = (x[33]);
  assign t[334] = (x[33]);
  assign t[335] = (x[36]);
  assign t[336] = (x[36]);
  assign t[337] = (x[41]);
  assign t[338] = (x[41]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[46]);
  assign t[341] = (x[49]);
  assign t[342] = (x[49]);
  assign t[343] = (x[52]);
  assign t[344] = (x[52]);
  assign t[345] = (x[55]);
  assign t[346] = (x[55]);
  assign t[347] = (x[60]);
  assign t[348] = (x[60]);
  assign t[349] = (x[65]);
  assign t[34] = t[51] ^ t[43];
  assign t[350] = (x[65]);
  assign t[351] = (x[68]);
  assign t[352] = (x[68]);
  assign t[353] = (x[71]);
  assign t[354] = (x[71]);
  assign t[355] = (x[74]);
  assign t[356] = (x[74]);
  assign t[357] = (x[77]);
  assign t[358] = (x[77]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[80]);
  assign t[361] = (x[83]);
  assign t[362] = (x[83]);
  assign t[363] = (x[86]);
  assign t[364] = (x[86]);
  assign t[365] = (x[89]);
  assign t[366] = (x[89]);
  assign t[367] = (x[92]);
  assign t[368] = (x[92]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[55];
  assign t[370] = (x[95]);
  assign t[371] = (x[98]);
  assign t[372] = (x[98]);
  assign t[373] = (x[101]);
  assign t[374] = (x[101]);
  assign t[375] = (x[104]);
  assign t[376] = (x[104]);
  assign t[377] = (x[107]);
  assign t[378] = (x[107]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[56] & t[57]);
  assign t[380] = (x[110]);
  assign t[381] = (x[113]);
  assign t[382] = (x[113]);
  assign t[383] = (x[116]);
  assign t[384] = (x[116]);
  assign t[385] = (x[119]);
  assign t[386] = (x[119]);
  assign t[387] = (x[122]);
  assign t[388] = (x[122]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[58] & t[118]);
  assign t[390] = (x[125]);
  assign t[391] = (x[128]);
  assign t[392] = (x[128]);
  assign t[393] = (x[131]);
  assign t[394] = (x[131]);
  assign t[395] = (x[134]);
  assign t[396] = (x[134]);
  assign t[397] = (x[137]);
  assign t[398] = (x[137]);
  assign t[39] = t[59] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[41];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[121]);
  assign t[51] = t[18] ? x[40] : x[39];
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[122]);
  assign t[54] = t[48] ? x[45] : x[44];
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = ~(t[83] & t[125]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[86] & t[126]);
  assign t[64] = t[59] ? x[59] : x[58];
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[91] & t[127]);
  assign t[68] = t[115] ? x[64] : x[63];
  assign t[69] = ~(t[120] & t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[130]);
  assign t[73] = ~(t[92] & t[93]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[94] & t[95]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[98] & t[133]);
  assign t[79] = ~(t[124] & t[123]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[99] & t[100]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[138]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[104]);
  assign t[88] = ~(t[105] & t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[141]);
  assign t[91] = ~(t[106] & t[107]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[145]);
  assign t[98] = ~(t[108] & t[109]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind186(x, y);
 input [139:0] x;
 output y;

 wire [389:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[2];
  assign t[145] = t[186] ^ x[10];
  assign t[146] = t[187] ^ x[13];
  assign t[147] = t[188] ^ x[16];
  assign t[148] = t[189] ^ x[19];
  assign t[149] = t[190] ^ x[22];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[27];
  assign t[151] = t[192] ^ x[32];
  assign t[152] = t[193] ^ x[35];
  assign t[153] = t[194] ^ x[38];
  assign t[154] = t[195] ^ x[43];
  assign t[155] = t[196] ^ x[48];
  assign t[156] = t[197] ^ x[51];
  assign t[157] = t[198] ^ x[54];
  assign t[158] = t[199] ^ x[57];
  assign t[159] = t[200] ^ x[62];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[67];
  assign t[161] = t[202] ^ x[70];
  assign t[162] = t[203] ^ x[73];
  assign t[163] = t[204] ^ x[76];
  assign t[164] = t[205] ^ x[79];
  assign t[165] = t[206] ^ x[82];
  assign t[166] = t[207] ^ x[85];
  assign t[167] = t[208] ^ x[88];
  assign t[168] = t[209] ^ x[91];
  assign t[169] = t[210] ^ x[94];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[100];
  assign t[172] = t[213] ^ x[103];
  assign t[173] = t[214] ^ x[106];
  assign t[174] = t[215] ^ x[109];
  assign t[175] = t[216] ^ x[112];
  assign t[176] = t[217] ^ x[115];
  assign t[177] = t[218] ^ x[118];
  assign t[178] = t[219] ^ x[121];
  assign t[179] = t[220] ^ x[124];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[127];
  assign t[181] = t[222] ^ x[130];
  assign t[182] = t[223] ^ x[133];
  assign t[183] = t[224] ^ x[136];
  assign t[184] = t[225] ^ x[139];
  assign t[185] = (t[226] & ~t[227]);
  assign t[186] = (t[228] & ~t[229]);
  assign t[187] = (t[230] & ~t[231]);
  assign t[188] = (t[232] & ~t[233]);
  assign t[189] = (t[234] & ~t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[236] & ~t[237]);
  assign t[191] = (t[238] & ~t[239]);
  assign t[192] = (t[240] & ~t[241]);
  assign t[193] = (t[242] & ~t[243]);
  assign t[194] = (t[244] & ~t[245]);
  assign t[195] = (t[246] & ~t[247]);
  assign t[196] = (t[248] & ~t[249]);
  assign t[197] = (t[250] & ~t[251]);
  assign t[198] = (t[252] & ~t[253]);
  assign t[199] = (t[254] & ~t[255]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[256] & ~t[257]);
  assign t[201] = (t[258] & ~t[259]);
  assign t[202] = (t[260] & ~t[261]);
  assign t[203] = (t[262] & ~t[263]);
  assign t[204] = (t[264] & ~t[265]);
  assign t[205] = (t[266] & ~t[267]);
  assign t[206] = (t[268] & ~t[269]);
  assign t[207] = (t[270] & ~t[271]);
  assign t[208] = (t[272] & ~t[273]);
  assign t[209] = (t[274] & ~t[275]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[276] & ~t[277]);
  assign t[211] = (t[278] & ~t[279]);
  assign t[212] = (t[280] & ~t[281]);
  assign t[213] = (t[282] & ~t[283]);
  assign t[214] = (t[284] & ~t[285]);
  assign t[215] = (t[286] & ~t[287]);
  assign t[216] = (t[288] & ~t[289]);
  assign t[217] = (t[290] & ~t[291]);
  assign t[218] = (t[292] & ~t[293]);
  assign t[219] = (t[294] & ~t[295]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[296] & ~t[297]);
  assign t[221] = (t[298] & ~t[299]);
  assign t[222] = (t[300] & ~t[301]);
  assign t[223] = (t[302] & ~t[303]);
  assign t[224] = (t[304] & ~t[305]);
  assign t[225] = (t[306] & ~t[307]);
  assign t[226] = t[308] ^ x[2];
  assign t[227] = t[309] ^ x[1];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[9];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[12];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[15];
  assign t[234] = t[316] ^ x[19];
  assign t[235] = t[317] ^ x[18];
  assign t[236] = t[318] ^ x[22];
  assign t[237] = t[319] ^ x[21];
  assign t[238] = t[320] ^ x[27];
  assign t[239] = t[321] ^ x[26];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[32];
  assign t[241] = t[323] ^ x[31];
  assign t[242] = t[324] ^ x[35];
  assign t[243] = t[325] ^ x[34];
  assign t[244] = t[326] ^ x[38];
  assign t[245] = t[327] ^ x[37];
  assign t[246] = t[328] ^ x[43];
  assign t[247] = t[329] ^ x[42];
  assign t[248] = t[330] ^ x[48];
  assign t[249] = t[331] ^ x[47];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[51];
  assign t[251] = t[333] ^ x[50];
  assign t[252] = t[334] ^ x[54];
  assign t[253] = t[335] ^ x[53];
  assign t[254] = t[336] ^ x[57];
  assign t[255] = t[337] ^ x[56];
  assign t[256] = t[338] ^ x[62];
  assign t[257] = t[339] ^ x[61];
  assign t[258] = t[340] ^ x[67];
  assign t[259] = t[341] ^ x[66];
  assign t[25] = ~(t[106]);
  assign t[260] = t[342] ^ x[70];
  assign t[261] = t[343] ^ x[69];
  assign t[262] = t[344] ^ x[73];
  assign t[263] = t[345] ^ x[72];
  assign t[264] = t[346] ^ x[76];
  assign t[265] = t[347] ^ x[75];
  assign t[266] = t[348] ^ x[79];
  assign t[267] = t[349] ^ x[78];
  assign t[268] = t[350] ^ x[82];
  assign t[269] = t[351] ^ x[81];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[85];
  assign t[271] = t[353] ^ x[84];
  assign t[272] = t[354] ^ x[88];
  assign t[273] = t[355] ^ x[87];
  assign t[274] = t[356] ^ x[91];
  assign t[275] = t[357] ^ x[90];
  assign t[276] = t[358] ^ x[94];
  assign t[277] = t[359] ^ x[93];
  assign t[278] = t[360] ^ x[97];
  assign t[279] = t[361] ^ x[96];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[100];
  assign t[281] = t[363] ^ x[99];
  assign t[282] = t[364] ^ x[103];
  assign t[283] = t[365] ^ x[102];
  assign t[284] = t[366] ^ x[106];
  assign t[285] = t[367] ^ x[105];
  assign t[286] = t[368] ^ x[109];
  assign t[287] = t[369] ^ x[108];
  assign t[288] = t[370] ^ x[112];
  assign t[289] = t[371] ^ x[111];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[115];
  assign t[291] = t[373] ^ x[114];
  assign t[292] = t[374] ^ x[118];
  assign t[293] = t[375] ^ x[117];
  assign t[294] = t[376] ^ x[121];
  assign t[295] = t[377] ^ x[120];
  assign t[296] = t[378] ^ x[124];
  assign t[297] = t[379] ^ x[123];
  assign t[298] = t[380] ^ x[127];
  assign t[299] = t[381] ^ x[126];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[130];
  assign t[301] = t[383] ^ x[129];
  assign t[302] = t[384] ^ x[133];
  assign t[303] = t[385] ^ x[132];
  assign t[304] = t[386] ^ x[136];
  assign t[305] = t[387] ^ x[135];
  assign t[306] = t[388] ^ x[139];
  assign t[307] = t[389] ^ x[138];
  assign t[308] = (x[0]);
  assign t[309] = (x[0]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[8]);
  assign t[312] = (x[11]);
  assign t[313] = (x[11]);
  assign t[314] = (x[14]);
  assign t[315] = (x[14]);
  assign t[316] = (x[17]);
  assign t[317] = (x[17]);
  assign t[318] = (x[20]);
  assign t[319] = (x[20]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[25]);
  assign t[321] = (x[25]);
  assign t[322] = (x[30]);
  assign t[323] = (x[30]);
  assign t[324] = (x[33]);
  assign t[325] = (x[33]);
  assign t[326] = (x[36]);
  assign t[327] = (x[36]);
  assign t[328] = (x[41]);
  assign t[329] = (x[41]);
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[46]);
  assign t[332] = (x[49]);
  assign t[333] = (x[49]);
  assign t[334] = (x[52]);
  assign t[335] = (x[52]);
  assign t[336] = (x[55]);
  assign t[337] = (x[55]);
  assign t[338] = (x[60]);
  assign t[339] = (x[60]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[65]);
  assign t[342] = (x[68]);
  assign t[343] = (x[68]);
  assign t[344] = (x[71]);
  assign t[345] = (x[71]);
  assign t[346] = (x[74]);
  assign t[347] = (x[74]);
  assign t[348] = (x[77]);
  assign t[349] = (x[77]);
  assign t[34] = t[50] ^ t[43];
  assign t[350] = (x[80]);
  assign t[351] = (x[80]);
  assign t[352] = (x[83]);
  assign t[353] = (x[83]);
  assign t[354] = (x[86]);
  assign t[355] = (x[86]);
  assign t[356] = (x[89]);
  assign t[357] = (x[89]);
  assign t[358] = (x[92]);
  assign t[359] = (x[92]);
  assign t[35] = ~(t[51] & t[52]);
  assign t[360] = (x[95]);
  assign t[361] = (x[95]);
  assign t[362] = (x[98]);
  assign t[363] = (x[98]);
  assign t[364] = (x[101]);
  assign t[365] = (x[101]);
  assign t[366] = (x[104]);
  assign t[367] = (x[104]);
  assign t[368] = (x[107]);
  assign t[369] = (x[107]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[110]);
  assign t[371] = (x[110]);
  assign t[372] = (x[113]);
  assign t[373] = (x[113]);
  assign t[374] = (x[116]);
  assign t[375] = (x[116]);
  assign t[376] = (x[119]);
  assign t[377] = (x[119]);
  assign t[378] = (x[122]);
  assign t[379] = (x[122]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[125]);
  assign t[382] = (x[128]);
  assign t[383] = (x[128]);
  assign t[384] = (x[131]);
  assign t[385] = (x[131]);
  assign t[386] = (x[134]);
  assign t[387] = (x[134]);
  assign t[388] = (x[137]);
  assign t[389] = (x[137]);
  assign t[38] = t[57] | t[109];
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[41];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[112];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[72] ? x[40] : x[39];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = t[75] | t[113];
  assign t[53] = t[18] ? x[45] : x[44];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = ~(t[114]);
  assign t[56] = ~(t[115]);
  assign t[57] = ~(t[78] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[81] | t[116];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[117];
  assign t[63] = t[58] ? x[59] : x[58];
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = t[89] | t[118];
  assign t[67] = t[58] ? x[64] : x[63];
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[91] | t[73]);
  assign t[76] = ~(t[92] & t[93]);
  assign t[77] = t[94] | t[124];
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[95] | t[79]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[96] | t[82]);
  assign t[85] = ~(t[97] & t[98]);
  assign t[86] = t[99] | t[130];
  assign t[87] = ~(t[131]);
  assign t[88] = ~(t[132]);
  assign t[89] = ~(t[100] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[101] | t[92]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[102] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [139:0] x;
 output y;

 wire [389:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[2];
  assign t[145] = t[186] ^ x[10];
  assign t[146] = t[187] ^ x[13];
  assign t[147] = t[188] ^ x[16];
  assign t[148] = t[189] ^ x[19];
  assign t[149] = t[190] ^ x[22];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[27];
  assign t[151] = t[192] ^ x[32];
  assign t[152] = t[193] ^ x[35];
  assign t[153] = t[194] ^ x[38];
  assign t[154] = t[195] ^ x[43];
  assign t[155] = t[196] ^ x[48];
  assign t[156] = t[197] ^ x[51];
  assign t[157] = t[198] ^ x[54];
  assign t[158] = t[199] ^ x[57];
  assign t[159] = t[200] ^ x[62];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[67];
  assign t[161] = t[202] ^ x[70];
  assign t[162] = t[203] ^ x[73];
  assign t[163] = t[204] ^ x[76];
  assign t[164] = t[205] ^ x[79];
  assign t[165] = t[206] ^ x[82];
  assign t[166] = t[207] ^ x[85];
  assign t[167] = t[208] ^ x[88];
  assign t[168] = t[209] ^ x[91];
  assign t[169] = t[210] ^ x[94];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[100];
  assign t[172] = t[213] ^ x[103];
  assign t[173] = t[214] ^ x[106];
  assign t[174] = t[215] ^ x[109];
  assign t[175] = t[216] ^ x[112];
  assign t[176] = t[217] ^ x[115];
  assign t[177] = t[218] ^ x[118];
  assign t[178] = t[219] ^ x[121];
  assign t[179] = t[220] ^ x[124];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[127];
  assign t[181] = t[222] ^ x[130];
  assign t[182] = t[223] ^ x[133];
  assign t[183] = t[224] ^ x[136];
  assign t[184] = t[225] ^ x[139];
  assign t[185] = (t[226] & ~t[227]);
  assign t[186] = (t[228] & ~t[229]);
  assign t[187] = (t[230] & ~t[231]);
  assign t[188] = (t[232] & ~t[233]);
  assign t[189] = (t[234] & ~t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[236] & ~t[237]);
  assign t[191] = (t[238] & ~t[239]);
  assign t[192] = (t[240] & ~t[241]);
  assign t[193] = (t[242] & ~t[243]);
  assign t[194] = (t[244] & ~t[245]);
  assign t[195] = (t[246] & ~t[247]);
  assign t[196] = (t[248] & ~t[249]);
  assign t[197] = (t[250] & ~t[251]);
  assign t[198] = (t[252] & ~t[253]);
  assign t[199] = (t[254] & ~t[255]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[256] & ~t[257]);
  assign t[201] = (t[258] & ~t[259]);
  assign t[202] = (t[260] & ~t[261]);
  assign t[203] = (t[262] & ~t[263]);
  assign t[204] = (t[264] & ~t[265]);
  assign t[205] = (t[266] & ~t[267]);
  assign t[206] = (t[268] & ~t[269]);
  assign t[207] = (t[270] & ~t[271]);
  assign t[208] = (t[272] & ~t[273]);
  assign t[209] = (t[274] & ~t[275]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[276] & ~t[277]);
  assign t[211] = (t[278] & ~t[279]);
  assign t[212] = (t[280] & ~t[281]);
  assign t[213] = (t[282] & ~t[283]);
  assign t[214] = (t[284] & ~t[285]);
  assign t[215] = (t[286] & ~t[287]);
  assign t[216] = (t[288] & ~t[289]);
  assign t[217] = (t[290] & ~t[291]);
  assign t[218] = (t[292] & ~t[293]);
  assign t[219] = (t[294] & ~t[295]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[296] & ~t[297]);
  assign t[221] = (t[298] & ~t[299]);
  assign t[222] = (t[300] & ~t[301]);
  assign t[223] = (t[302] & ~t[303]);
  assign t[224] = (t[304] & ~t[305]);
  assign t[225] = (t[306] & ~t[307]);
  assign t[226] = t[308] ^ x[2];
  assign t[227] = t[309] ^ x[1];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[9];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[12];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[15];
  assign t[234] = t[316] ^ x[19];
  assign t[235] = t[317] ^ x[18];
  assign t[236] = t[318] ^ x[22];
  assign t[237] = t[319] ^ x[21];
  assign t[238] = t[320] ^ x[27];
  assign t[239] = t[321] ^ x[26];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[32];
  assign t[241] = t[323] ^ x[31];
  assign t[242] = t[324] ^ x[35];
  assign t[243] = t[325] ^ x[34];
  assign t[244] = t[326] ^ x[38];
  assign t[245] = t[327] ^ x[37];
  assign t[246] = t[328] ^ x[43];
  assign t[247] = t[329] ^ x[42];
  assign t[248] = t[330] ^ x[48];
  assign t[249] = t[331] ^ x[47];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[51];
  assign t[251] = t[333] ^ x[50];
  assign t[252] = t[334] ^ x[54];
  assign t[253] = t[335] ^ x[53];
  assign t[254] = t[336] ^ x[57];
  assign t[255] = t[337] ^ x[56];
  assign t[256] = t[338] ^ x[62];
  assign t[257] = t[339] ^ x[61];
  assign t[258] = t[340] ^ x[67];
  assign t[259] = t[341] ^ x[66];
  assign t[25] = ~(t[106]);
  assign t[260] = t[342] ^ x[70];
  assign t[261] = t[343] ^ x[69];
  assign t[262] = t[344] ^ x[73];
  assign t[263] = t[345] ^ x[72];
  assign t[264] = t[346] ^ x[76];
  assign t[265] = t[347] ^ x[75];
  assign t[266] = t[348] ^ x[79];
  assign t[267] = t[349] ^ x[78];
  assign t[268] = t[350] ^ x[82];
  assign t[269] = t[351] ^ x[81];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[85];
  assign t[271] = t[353] ^ x[84];
  assign t[272] = t[354] ^ x[88];
  assign t[273] = t[355] ^ x[87];
  assign t[274] = t[356] ^ x[91];
  assign t[275] = t[357] ^ x[90];
  assign t[276] = t[358] ^ x[94];
  assign t[277] = t[359] ^ x[93];
  assign t[278] = t[360] ^ x[97];
  assign t[279] = t[361] ^ x[96];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[100];
  assign t[281] = t[363] ^ x[99];
  assign t[282] = t[364] ^ x[103];
  assign t[283] = t[365] ^ x[102];
  assign t[284] = t[366] ^ x[106];
  assign t[285] = t[367] ^ x[105];
  assign t[286] = t[368] ^ x[109];
  assign t[287] = t[369] ^ x[108];
  assign t[288] = t[370] ^ x[112];
  assign t[289] = t[371] ^ x[111];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[115];
  assign t[291] = t[373] ^ x[114];
  assign t[292] = t[374] ^ x[118];
  assign t[293] = t[375] ^ x[117];
  assign t[294] = t[376] ^ x[121];
  assign t[295] = t[377] ^ x[120];
  assign t[296] = t[378] ^ x[124];
  assign t[297] = t[379] ^ x[123];
  assign t[298] = t[380] ^ x[127];
  assign t[299] = t[381] ^ x[126];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[130];
  assign t[301] = t[383] ^ x[129];
  assign t[302] = t[384] ^ x[133];
  assign t[303] = t[385] ^ x[132];
  assign t[304] = t[386] ^ x[136];
  assign t[305] = t[387] ^ x[135];
  assign t[306] = t[388] ^ x[139];
  assign t[307] = t[389] ^ x[138];
  assign t[308] = (x[0]);
  assign t[309] = (x[0]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[8]);
  assign t[312] = (x[11]);
  assign t[313] = (x[11]);
  assign t[314] = (x[14]);
  assign t[315] = (x[14]);
  assign t[316] = (x[17]);
  assign t[317] = (x[17]);
  assign t[318] = (x[20]);
  assign t[319] = (x[20]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[25]);
  assign t[321] = (x[25]);
  assign t[322] = (x[30]);
  assign t[323] = (x[30]);
  assign t[324] = (x[33]);
  assign t[325] = (x[33]);
  assign t[326] = (x[36]);
  assign t[327] = (x[36]);
  assign t[328] = (x[41]);
  assign t[329] = (x[41]);
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[46]);
  assign t[332] = (x[49]);
  assign t[333] = (x[49]);
  assign t[334] = (x[52]);
  assign t[335] = (x[52]);
  assign t[336] = (x[55]);
  assign t[337] = (x[55]);
  assign t[338] = (x[60]);
  assign t[339] = (x[60]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[65]);
  assign t[342] = (x[68]);
  assign t[343] = (x[68]);
  assign t[344] = (x[71]);
  assign t[345] = (x[71]);
  assign t[346] = (x[74]);
  assign t[347] = (x[74]);
  assign t[348] = (x[77]);
  assign t[349] = (x[77]);
  assign t[34] = t[50] ^ t[43];
  assign t[350] = (x[80]);
  assign t[351] = (x[80]);
  assign t[352] = (x[83]);
  assign t[353] = (x[83]);
  assign t[354] = (x[86]);
  assign t[355] = (x[86]);
  assign t[356] = (x[89]);
  assign t[357] = (x[89]);
  assign t[358] = (x[92]);
  assign t[359] = (x[92]);
  assign t[35] = ~(t[51] & t[52]);
  assign t[360] = (x[95]);
  assign t[361] = (x[95]);
  assign t[362] = (x[98]);
  assign t[363] = (x[98]);
  assign t[364] = (x[101]);
  assign t[365] = (x[101]);
  assign t[366] = (x[104]);
  assign t[367] = (x[104]);
  assign t[368] = (x[107]);
  assign t[369] = (x[107]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[110]);
  assign t[371] = (x[110]);
  assign t[372] = (x[113]);
  assign t[373] = (x[113]);
  assign t[374] = (x[116]);
  assign t[375] = (x[116]);
  assign t[376] = (x[119]);
  assign t[377] = (x[119]);
  assign t[378] = (x[122]);
  assign t[379] = (x[122]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[125]);
  assign t[382] = (x[128]);
  assign t[383] = (x[128]);
  assign t[384] = (x[131]);
  assign t[385] = (x[131]);
  assign t[386] = (x[134]);
  assign t[387] = (x[134]);
  assign t[388] = (x[137]);
  assign t[389] = (x[137]);
  assign t[38] = t[57] | t[109];
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[41];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[112];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[72] ? x[40] : x[39];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = t[75] | t[113];
  assign t[53] = t[18] ? x[45] : x[44];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = ~(t[114]);
  assign t[56] = ~(t[115]);
  assign t[57] = ~(t[78] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[81] | t[116];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[117];
  assign t[63] = t[58] ? x[59] : x[58];
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = t[89] | t[118];
  assign t[67] = t[58] ? x[64] : x[63];
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[91] | t[73]);
  assign t[76] = ~(t[92] & t[93]);
  assign t[77] = t[94] | t[124];
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[95] | t[79]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[96] | t[82]);
  assign t[85] = ~(t[97] & t[98]);
  assign t[86] = t[99] | t[130];
  assign t[87] = ~(t[131]);
  assign t[88] = ~(t[132]);
  assign t[89] = ~(t[100] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[101] | t[92]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[102] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [106:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = t[1] ? t[2] : t[162];
  assign t[100] = t[63] & t[163];
  assign t[101] = ~(t[185]);
  assign t[102] = ~(t[177] | t[178]);
  assign t[103] = ~(t[186]);
  assign t[104] = ~(t[187]);
  assign t[105] = ~(t[126] | t[127]);
  assign t[106] = ~(t[43] | t[128]);
  assign t[107] = ~(t[42] | t[129]);
  assign t[108] = ~(t[188]);
  assign t[109] = ~(t[180] | t[181]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[189]);
  assign t[111] = ~(t[190]);
  assign t[112] = ~(t[130] | t[131]);
  assign t[113] = ~(t[132] | t[133]);
  assign t[114] = ~(t[117] | t[134]);
  assign t[115] = ~(t[191]);
  assign t[116] = ~(t[183] | t[184]);
  assign t[117] = ~(t[63] | t[135]);
  assign t[118] = ~(t[63] | t[136]);
  assign t[119] = t[44] | t[137];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[138] & t[139]);
  assign t[121] = x[4] & t[164];
  assign t[122] = ~(x[4] | t[164]);
  assign t[123] = ~(t[166]);
  assign t[124] = t[163] ? t[95] : t[94];
  assign t[125] = t[163] ? t[141] : t[140];
  assign t[126] = ~(t[192]);
  assign t[127] = ~(t[186] | t[187]);
  assign t[128] = ~(t[63] | t[142]);
  assign t[129] = ~(t[114] & t[139]);
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[193]);
  assign t[131] = ~(t[189] | t[190]);
  assign t[132] = ~(t[106] & t[143]);
  assign t[133] = ~(t[144] & t[139]);
  assign t[134] = ~(t[63] | t[145]);
  assign t[135] = t[163] ? t[93] : t[94];
  assign t[136] = t[163] ? t[140] : t[146];
  assign t[137] = ~(t[63] | t[147]);
  assign t[138] = ~(t[148] | t[149]);
  assign t[139] = t[66] | t[150];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(x[4] & t[151]);
  assign t[141] = ~(t[152] & t[123]);
  assign t[142] = t[163] ? t[141] : t[153];
  assign t[143] = ~(t[66] & t[154]);
  assign t[144] = ~(t[155] & t[156]);
  assign t[145] = t[163] ? t[95] : t[96];
  assign t[146] = ~(t[166] & t[152]);
  assign t[147] = t[163] ? t[146] : t[140];
  assign t[148] = ~(t[157]);
  assign t[149] = ~(t[63] | t[158]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[163] ? t[140] : t[141];
  assign t[151] = ~(t[164] | t[166]);
  assign t[152] = ~(x[4] | t[159]);
  assign t[153] = ~(x[4] & t[99]);
  assign t[154] = ~(t[140] & t[146]);
  assign t[155] = t[166] & t[160];
  assign t[156] = t[122] | t[121];
  assign t[157] = ~(t[160] & t[161]);
  assign t[158] = t[163] ? t[153] : t[141];
  assign t[159] = ~(t[164]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = ~(t[66] | t[163]);
  assign t[161] = ~(t[146] & t[153]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[163] & t[164]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[165] & t[166]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = (t[216]);
  assign t[185] = (t[217]);
  assign t[186] = (t[218]);
  assign t[187] = (t[219]);
  assign t[188] = (t[220]);
  assign t[189] = (t[221]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (t[222]);
  assign t[191] = (t[223]);
  assign t[192] = (t[224]);
  assign t[193] = (t[225]);
  assign t[194] = t[226] ^ x[2];
  assign t[195] = t[227] ^ x[10];
  assign t[196] = t[228] ^ x[13];
  assign t[197] = t[229] ^ x[16];
  assign t[198] = t[230] ^ x[19];
  assign t[199] = t[231] ^ x[22];
  assign t[19] = t[27] ? x[6] : x[7];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[25];
  assign t[201] = t[233] ^ x[28];
  assign t[202] = t[234] ^ x[31];
  assign t[203] = t[235] ^ x[34];
  assign t[204] = t[236] ^ x[37];
  assign t[205] = t[237] ^ x[40];
  assign t[206] = t[238] ^ x[43];
  assign t[207] = t[239] ^ x[46];
  assign t[208] = t[240] ^ x[51];
  assign t[209] = t[241] ^ x[54];
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = t[242] ^ x[57];
  assign t[211] = t[243] ^ x[60];
  assign t[212] = t[244] ^ x[65];
  assign t[213] = t[245] ^ x[68];
  assign t[214] = t[246] ^ x[71];
  assign t[215] = t[247] ^ x[76];
  assign t[216] = t[248] ^ x[79];
  assign t[217] = t[249] ^ x[82];
  assign t[218] = t[250] ^ x[85];
  assign t[219] = t[251] ^ x[88];
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = t[252] ^ x[91];
  assign t[221] = t[253] ^ x[94];
  assign t[222] = t[254] ^ x[97];
  assign t[223] = t[255] ^ x[100];
  assign t[224] = t[256] ^ x[103];
  assign t[225] = t[257] ^ x[106];
  assign t[226] = (t[258] & ~t[259]);
  assign t[227] = (t[260] & ~t[261]);
  assign t[228] = (t[262] & ~t[263]);
  assign t[229] = (t[264] & ~t[265]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (t[266] & ~t[267]);
  assign t[231] = (t[268] & ~t[269]);
  assign t[232] = (t[270] & ~t[271]);
  assign t[233] = (t[272] & ~t[273]);
  assign t[234] = (t[274] & ~t[275]);
  assign t[235] = (t[276] & ~t[277]);
  assign t[236] = (t[278] & ~t[279]);
  assign t[237] = (t[280] & ~t[281]);
  assign t[238] = (t[282] & ~t[283]);
  assign t[239] = (t[284] & ~t[285]);
  assign t[23] = x[4] ? t[33] : t[32];
  assign t[240] = (t[286] & ~t[287]);
  assign t[241] = (t[288] & ~t[289]);
  assign t[242] = (t[290] & ~t[291]);
  assign t[243] = (t[292] & ~t[293]);
  assign t[244] = (t[294] & ~t[295]);
  assign t[245] = (t[296] & ~t[297]);
  assign t[246] = (t[298] & ~t[299]);
  assign t[247] = (t[300] & ~t[301]);
  assign t[248] = (t[302] & ~t[303]);
  assign t[249] = (t[304] & ~t[305]);
  assign t[24] = x[4] ? t[35] : t[34];
  assign t[250] = (t[306] & ~t[307]);
  assign t[251] = (t[308] & ~t[309]);
  assign t[252] = (t[310] & ~t[311]);
  assign t[253] = (t[312] & ~t[313]);
  assign t[254] = (t[314] & ~t[315]);
  assign t[255] = (t[316] & ~t[317]);
  assign t[256] = (t[318] & ~t[319]);
  assign t[257] = (t[320] & ~t[321]);
  assign t[258] = t[322] ^ x[2];
  assign t[259] = t[323] ^ x[1];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[324] ^ x[10];
  assign t[261] = t[325] ^ x[9];
  assign t[262] = t[326] ^ x[13];
  assign t[263] = t[327] ^ x[12];
  assign t[264] = t[328] ^ x[16];
  assign t[265] = t[329] ^ x[15];
  assign t[266] = t[330] ^ x[19];
  assign t[267] = t[331] ^ x[18];
  assign t[268] = t[332] ^ x[22];
  assign t[269] = t[333] ^ x[21];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[334] ^ x[25];
  assign t[271] = t[335] ^ x[24];
  assign t[272] = t[336] ^ x[28];
  assign t[273] = t[337] ^ x[27];
  assign t[274] = t[338] ^ x[31];
  assign t[275] = t[339] ^ x[30];
  assign t[276] = t[340] ^ x[34];
  assign t[277] = t[341] ^ x[33];
  assign t[278] = t[342] ^ x[37];
  assign t[279] = t[343] ^ x[36];
  assign t[27] = ~(t[40]);
  assign t[280] = t[344] ^ x[40];
  assign t[281] = t[345] ^ x[39];
  assign t[282] = t[346] ^ x[43];
  assign t[283] = t[347] ^ x[42];
  assign t[284] = t[348] ^ x[46];
  assign t[285] = t[349] ^ x[45];
  assign t[286] = t[350] ^ x[51];
  assign t[287] = t[351] ^ x[50];
  assign t[288] = t[352] ^ x[54];
  assign t[289] = t[353] ^ x[53];
  assign t[28] = ~(t[41] | t[42]);
  assign t[290] = t[354] ^ x[57];
  assign t[291] = t[355] ^ x[56];
  assign t[292] = t[356] ^ x[60];
  assign t[293] = t[357] ^ x[59];
  assign t[294] = t[358] ^ x[65];
  assign t[295] = t[359] ^ x[64];
  assign t[296] = t[360] ^ x[68];
  assign t[297] = t[361] ^ x[67];
  assign t[298] = t[362] ^ x[71];
  assign t[299] = t[363] ^ x[70];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[364] ^ x[76];
  assign t[301] = t[365] ^ x[75];
  assign t[302] = t[366] ^ x[79];
  assign t[303] = t[367] ^ x[78];
  assign t[304] = t[368] ^ x[82];
  assign t[305] = t[369] ^ x[81];
  assign t[306] = t[370] ^ x[85];
  assign t[307] = t[371] ^ x[84];
  assign t[308] = t[372] ^ x[88];
  assign t[309] = t[373] ^ x[87];
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = t[374] ^ x[91];
  assign t[311] = t[375] ^ x[90];
  assign t[312] = t[376] ^ x[94];
  assign t[313] = t[377] ^ x[93];
  assign t[314] = t[378] ^ x[97];
  assign t[315] = t[379] ^ x[96];
  assign t[316] = t[380] ^ x[100];
  assign t[317] = t[381] ^ x[99];
  assign t[318] = t[382] ^ x[103];
  assign t[319] = t[383] ^ x[102];
  assign t[31] = ~(t[167] | t[47]);
  assign t[320] = t[384] ^ x[106];
  assign t[321] = t[385] ^ x[105];
  assign t[322] = (x[0]);
  assign t[323] = (x[0]);
  assign t[324] = (x[8]);
  assign t[325] = (x[8]);
  assign t[326] = (x[11]);
  assign t[327] = (x[11]);
  assign t[328] = (x[14]);
  assign t[329] = (x[14]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[17]);
  assign t[331] = (x[17]);
  assign t[332] = (x[20]);
  assign t[333] = (x[20]);
  assign t[334] = (x[23]);
  assign t[335] = (x[23]);
  assign t[336] = (x[26]);
  assign t[337] = (x[26]);
  assign t[338] = (x[29]);
  assign t[339] = (x[29]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = (x[32]);
  assign t[341] = (x[32]);
  assign t[342] = (x[35]);
  assign t[343] = (x[35]);
  assign t[344] = (x[38]);
  assign t[345] = (x[38]);
  assign t[346] = (x[41]);
  assign t[347] = (x[41]);
  assign t[348] = (x[44]);
  assign t[349] = (x[44]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = (x[49]);
  assign t[351] = (x[49]);
  assign t[352] = (x[52]);
  assign t[353] = (x[52]);
  assign t[354] = (x[55]);
  assign t[355] = (x[55]);
  assign t[356] = (x[58]);
  assign t[357] = (x[58]);
  assign t[358] = (x[63]);
  assign t[359] = (x[63]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = (x[66]);
  assign t[361] = (x[66]);
  assign t[362] = (x[69]);
  assign t[363] = (x[69]);
  assign t[364] = (x[74]);
  assign t[365] = (x[74]);
  assign t[366] = (x[77]);
  assign t[367] = (x[77]);
  assign t[368] = (x[80]);
  assign t[369] = (x[80]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (x[83]);
  assign t[371] = (x[83]);
  assign t[372] = (x[86]);
  assign t[373] = (x[86]);
  assign t[374] = (x[89]);
  assign t[375] = (x[89]);
  assign t[376] = (x[92]);
  assign t[377] = (x[92]);
  assign t[378] = (x[95]);
  assign t[379] = (x[95]);
  assign t[37] = ~(t[168] | t[58]);
  assign t[380] = (x[98]);
  assign t[381] = (x[98]);
  assign t[382] = (x[101]);
  assign t[383] = (x[101]);
  assign t[384] = (x[104]);
  assign t[385] = (x[104]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[165]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[63] | t[65]);
  assign t[43] = ~(t[66] | t[67]);
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = ~(t[169]);
  assign t[46] = ~(t[170]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[171] | t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[172] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[173]);
  assign t[57] = ~(t[174]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[175] | t[90]);
  assign t[61] = t[27] ? x[48] : x[47];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[66]);
  assign t[64] = t[163] ? t[94] : t[93];
  assign t[65] = t[163] ? t[96] : t[95];
  assign t[66] = ~(t[165]);
  assign t[67] = t[163] ? t[94] : t[95];
  assign t[68] = ~(t[97] | t[98]);
  assign t[69] = ~(t[99] & t[100]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[176]);
  assign t[71] = ~(t[169] | t[170]);
  assign t[72] = ~(t[177]);
  assign t[73] = ~(t[178]);
  assign t[74] = ~(t[101] | t[102]);
  assign t[75] = ~(t[103] | t[104]);
  assign t[76] = ~(t[179] | t[105]);
  assign t[77] = t[27] ? x[62] : x[61];
  assign t[78] = ~(t[106] & t[107]);
  assign t[79] = ~(t[180]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[181]);
  assign t[81] = ~(t[108] | t[109]);
  assign t[82] = ~(t[110] | t[111]);
  assign t[83] = ~(t[182] | t[112]);
  assign t[84] = t[27] ? x[73] : x[72];
  assign t[85] = ~(t[113] & t[114]);
  assign t[86] = ~(t[162]);
  assign t[87] = ~(t[173] | t[174]);
  assign t[88] = ~(t[183]);
  assign t[89] = ~(t[184]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[115] | t[116]);
  assign t[91] = ~(t[117] | t[118]);
  assign t[92] = ~(t[119] | t[120]);
  assign t[93] = ~(t[121] & t[166]);
  assign t[94] = ~(t[122] & t[123]);
  assign t[95] = ~(t[121] & t[123]);
  assign t[96] = ~(t[122] & t[166]);
  assign t[97] = ~(t[66] | t[124]);
  assign t[98] = ~(t[66] | t[125]);
  assign t[99] = ~(t[164] | t[123]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [106:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = t[1] ? t[2] : t[162];
  assign t[100] = t[63] & t[163];
  assign t[101] = ~(t[185]);
  assign t[102] = ~(t[177] | t[178]);
  assign t[103] = ~(t[186]);
  assign t[104] = ~(t[187]);
  assign t[105] = ~(t[126] | t[127]);
  assign t[106] = ~(t[43] | t[128]);
  assign t[107] = ~(t[42] | t[129]);
  assign t[108] = ~(t[188]);
  assign t[109] = ~(t[180] | t[181]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[189]);
  assign t[111] = ~(t[190]);
  assign t[112] = ~(t[130] | t[131]);
  assign t[113] = ~(t[132] | t[133]);
  assign t[114] = ~(t[117] | t[134]);
  assign t[115] = ~(t[191]);
  assign t[116] = ~(t[183] | t[184]);
  assign t[117] = ~(t[63] | t[135]);
  assign t[118] = ~(t[63] | t[136]);
  assign t[119] = t[44] | t[137];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[138] & t[139]);
  assign t[121] = x[4] & t[164];
  assign t[122] = ~(x[4] | t[164]);
  assign t[123] = ~(t[166]);
  assign t[124] = t[163] ? t[95] : t[94];
  assign t[125] = t[163] ? t[141] : t[140];
  assign t[126] = ~(t[192]);
  assign t[127] = ~(t[186] | t[187]);
  assign t[128] = ~(t[63] | t[142]);
  assign t[129] = ~(t[114] & t[139]);
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[193]);
  assign t[131] = ~(t[189] | t[190]);
  assign t[132] = ~(t[106] & t[143]);
  assign t[133] = ~(t[144] & t[139]);
  assign t[134] = ~(t[63] | t[145]);
  assign t[135] = t[163] ? t[93] : t[94];
  assign t[136] = t[163] ? t[140] : t[146];
  assign t[137] = ~(t[63] | t[147]);
  assign t[138] = ~(t[148] | t[149]);
  assign t[139] = t[66] | t[150];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(x[4] & t[151]);
  assign t[141] = ~(t[152] & t[123]);
  assign t[142] = t[163] ? t[141] : t[153];
  assign t[143] = ~(t[66] & t[154]);
  assign t[144] = ~(t[155] & t[156]);
  assign t[145] = t[163] ? t[95] : t[96];
  assign t[146] = ~(t[166] & t[152]);
  assign t[147] = t[163] ? t[146] : t[140];
  assign t[148] = ~(t[157]);
  assign t[149] = ~(t[63] | t[158]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[163] ? t[140] : t[141];
  assign t[151] = ~(t[164] | t[166]);
  assign t[152] = ~(x[4] | t[159]);
  assign t[153] = ~(x[4] & t[99]);
  assign t[154] = ~(t[140] & t[146]);
  assign t[155] = t[166] & t[160];
  assign t[156] = t[122] | t[121];
  assign t[157] = ~(t[160] & t[161]);
  assign t[158] = t[163] ? t[153] : t[141];
  assign t[159] = ~(t[164]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = ~(t[66] | t[163]);
  assign t[161] = ~(t[146] & t[153]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[163] & t[164]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[165] & t[166]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = (t[216]);
  assign t[185] = (t[217]);
  assign t[186] = (t[218]);
  assign t[187] = (t[219]);
  assign t[188] = (t[220]);
  assign t[189] = (t[221]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (t[222]);
  assign t[191] = (t[223]);
  assign t[192] = (t[224]);
  assign t[193] = (t[225]);
  assign t[194] = t[226] ^ x[2];
  assign t[195] = t[227] ^ x[10];
  assign t[196] = t[228] ^ x[13];
  assign t[197] = t[229] ^ x[16];
  assign t[198] = t[230] ^ x[19];
  assign t[199] = t[231] ^ x[22];
  assign t[19] = t[27] ? x[6] : x[7];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[25];
  assign t[201] = t[233] ^ x[28];
  assign t[202] = t[234] ^ x[31];
  assign t[203] = t[235] ^ x[34];
  assign t[204] = t[236] ^ x[37];
  assign t[205] = t[237] ^ x[40];
  assign t[206] = t[238] ^ x[43];
  assign t[207] = t[239] ^ x[46];
  assign t[208] = t[240] ^ x[51];
  assign t[209] = t[241] ^ x[54];
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = t[242] ^ x[57];
  assign t[211] = t[243] ^ x[60];
  assign t[212] = t[244] ^ x[65];
  assign t[213] = t[245] ^ x[68];
  assign t[214] = t[246] ^ x[71];
  assign t[215] = t[247] ^ x[76];
  assign t[216] = t[248] ^ x[79];
  assign t[217] = t[249] ^ x[82];
  assign t[218] = t[250] ^ x[85];
  assign t[219] = t[251] ^ x[88];
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = t[252] ^ x[91];
  assign t[221] = t[253] ^ x[94];
  assign t[222] = t[254] ^ x[97];
  assign t[223] = t[255] ^ x[100];
  assign t[224] = t[256] ^ x[103];
  assign t[225] = t[257] ^ x[106];
  assign t[226] = (t[258] & ~t[259]);
  assign t[227] = (t[260] & ~t[261]);
  assign t[228] = (t[262] & ~t[263]);
  assign t[229] = (t[264] & ~t[265]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (t[266] & ~t[267]);
  assign t[231] = (t[268] & ~t[269]);
  assign t[232] = (t[270] & ~t[271]);
  assign t[233] = (t[272] & ~t[273]);
  assign t[234] = (t[274] & ~t[275]);
  assign t[235] = (t[276] & ~t[277]);
  assign t[236] = (t[278] & ~t[279]);
  assign t[237] = (t[280] & ~t[281]);
  assign t[238] = (t[282] & ~t[283]);
  assign t[239] = (t[284] & ~t[285]);
  assign t[23] = x[4] ? t[33] : t[32];
  assign t[240] = (t[286] & ~t[287]);
  assign t[241] = (t[288] & ~t[289]);
  assign t[242] = (t[290] & ~t[291]);
  assign t[243] = (t[292] & ~t[293]);
  assign t[244] = (t[294] & ~t[295]);
  assign t[245] = (t[296] & ~t[297]);
  assign t[246] = (t[298] & ~t[299]);
  assign t[247] = (t[300] & ~t[301]);
  assign t[248] = (t[302] & ~t[303]);
  assign t[249] = (t[304] & ~t[305]);
  assign t[24] = x[4] ? t[35] : t[34];
  assign t[250] = (t[306] & ~t[307]);
  assign t[251] = (t[308] & ~t[309]);
  assign t[252] = (t[310] & ~t[311]);
  assign t[253] = (t[312] & ~t[313]);
  assign t[254] = (t[314] & ~t[315]);
  assign t[255] = (t[316] & ~t[317]);
  assign t[256] = (t[318] & ~t[319]);
  assign t[257] = (t[320] & ~t[321]);
  assign t[258] = t[322] ^ x[2];
  assign t[259] = t[323] ^ x[1];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[324] ^ x[10];
  assign t[261] = t[325] ^ x[9];
  assign t[262] = t[326] ^ x[13];
  assign t[263] = t[327] ^ x[12];
  assign t[264] = t[328] ^ x[16];
  assign t[265] = t[329] ^ x[15];
  assign t[266] = t[330] ^ x[19];
  assign t[267] = t[331] ^ x[18];
  assign t[268] = t[332] ^ x[22];
  assign t[269] = t[333] ^ x[21];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[334] ^ x[25];
  assign t[271] = t[335] ^ x[24];
  assign t[272] = t[336] ^ x[28];
  assign t[273] = t[337] ^ x[27];
  assign t[274] = t[338] ^ x[31];
  assign t[275] = t[339] ^ x[30];
  assign t[276] = t[340] ^ x[34];
  assign t[277] = t[341] ^ x[33];
  assign t[278] = t[342] ^ x[37];
  assign t[279] = t[343] ^ x[36];
  assign t[27] = ~(t[40]);
  assign t[280] = t[344] ^ x[40];
  assign t[281] = t[345] ^ x[39];
  assign t[282] = t[346] ^ x[43];
  assign t[283] = t[347] ^ x[42];
  assign t[284] = t[348] ^ x[46];
  assign t[285] = t[349] ^ x[45];
  assign t[286] = t[350] ^ x[51];
  assign t[287] = t[351] ^ x[50];
  assign t[288] = t[352] ^ x[54];
  assign t[289] = t[353] ^ x[53];
  assign t[28] = ~(t[41] | t[42]);
  assign t[290] = t[354] ^ x[57];
  assign t[291] = t[355] ^ x[56];
  assign t[292] = t[356] ^ x[60];
  assign t[293] = t[357] ^ x[59];
  assign t[294] = t[358] ^ x[65];
  assign t[295] = t[359] ^ x[64];
  assign t[296] = t[360] ^ x[68];
  assign t[297] = t[361] ^ x[67];
  assign t[298] = t[362] ^ x[71];
  assign t[299] = t[363] ^ x[70];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[364] ^ x[76];
  assign t[301] = t[365] ^ x[75];
  assign t[302] = t[366] ^ x[79];
  assign t[303] = t[367] ^ x[78];
  assign t[304] = t[368] ^ x[82];
  assign t[305] = t[369] ^ x[81];
  assign t[306] = t[370] ^ x[85];
  assign t[307] = t[371] ^ x[84];
  assign t[308] = t[372] ^ x[88];
  assign t[309] = t[373] ^ x[87];
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = t[374] ^ x[91];
  assign t[311] = t[375] ^ x[90];
  assign t[312] = t[376] ^ x[94];
  assign t[313] = t[377] ^ x[93];
  assign t[314] = t[378] ^ x[97];
  assign t[315] = t[379] ^ x[96];
  assign t[316] = t[380] ^ x[100];
  assign t[317] = t[381] ^ x[99];
  assign t[318] = t[382] ^ x[103];
  assign t[319] = t[383] ^ x[102];
  assign t[31] = ~(t[167] | t[47]);
  assign t[320] = t[384] ^ x[106];
  assign t[321] = t[385] ^ x[105];
  assign t[322] = (x[0]);
  assign t[323] = (x[0]);
  assign t[324] = (x[8]);
  assign t[325] = (x[8]);
  assign t[326] = (x[11]);
  assign t[327] = (x[11]);
  assign t[328] = (x[14]);
  assign t[329] = (x[14]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[17]);
  assign t[331] = (x[17]);
  assign t[332] = (x[20]);
  assign t[333] = (x[20]);
  assign t[334] = (x[23]);
  assign t[335] = (x[23]);
  assign t[336] = (x[26]);
  assign t[337] = (x[26]);
  assign t[338] = (x[29]);
  assign t[339] = (x[29]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = (x[32]);
  assign t[341] = (x[32]);
  assign t[342] = (x[35]);
  assign t[343] = (x[35]);
  assign t[344] = (x[38]);
  assign t[345] = (x[38]);
  assign t[346] = (x[41]);
  assign t[347] = (x[41]);
  assign t[348] = (x[44]);
  assign t[349] = (x[44]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = (x[49]);
  assign t[351] = (x[49]);
  assign t[352] = (x[52]);
  assign t[353] = (x[52]);
  assign t[354] = (x[55]);
  assign t[355] = (x[55]);
  assign t[356] = (x[58]);
  assign t[357] = (x[58]);
  assign t[358] = (x[63]);
  assign t[359] = (x[63]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = (x[66]);
  assign t[361] = (x[66]);
  assign t[362] = (x[69]);
  assign t[363] = (x[69]);
  assign t[364] = (x[74]);
  assign t[365] = (x[74]);
  assign t[366] = (x[77]);
  assign t[367] = (x[77]);
  assign t[368] = (x[80]);
  assign t[369] = (x[80]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (x[83]);
  assign t[371] = (x[83]);
  assign t[372] = (x[86]);
  assign t[373] = (x[86]);
  assign t[374] = (x[89]);
  assign t[375] = (x[89]);
  assign t[376] = (x[92]);
  assign t[377] = (x[92]);
  assign t[378] = (x[95]);
  assign t[379] = (x[95]);
  assign t[37] = ~(t[168] | t[58]);
  assign t[380] = (x[98]);
  assign t[381] = (x[98]);
  assign t[382] = (x[101]);
  assign t[383] = (x[101]);
  assign t[384] = (x[104]);
  assign t[385] = (x[104]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[165]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[63] | t[65]);
  assign t[43] = ~(t[66] | t[67]);
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = ~(t[169]);
  assign t[46] = ~(t[170]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[171] | t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[172] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[173]);
  assign t[57] = ~(t[174]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[175] | t[90]);
  assign t[61] = t[27] ? x[48] : x[47];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[66]);
  assign t[64] = t[163] ? t[94] : t[93];
  assign t[65] = t[163] ? t[96] : t[95];
  assign t[66] = ~(t[165]);
  assign t[67] = t[163] ? t[94] : t[95];
  assign t[68] = ~(t[97] | t[98]);
  assign t[69] = ~(t[99] & t[100]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[176]);
  assign t[71] = ~(t[169] | t[170]);
  assign t[72] = ~(t[177]);
  assign t[73] = ~(t[178]);
  assign t[74] = ~(t[101] | t[102]);
  assign t[75] = ~(t[103] | t[104]);
  assign t[76] = ~(t[179] | t[105]);
  assign t[77] = t[27] ? x[62] : x[61];
  assign t[78] = ~(t[106] & t[107]);
  assign t[79] = ~(t[180]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[181]);
  assign t[81] = ~(t[108] | t[109]);
  assign t[82] = ~(t[110] | t[111]);
  assign t[83] = ~(t[182] | t[112]);
  assign t[84] = t[27] ? x[73] : x[72];
  assign t[85] = ~(t[113] & t[114]);
  assign t[86] = ~(t[162]);
  assign t[87] = ~(t[173] | t[174]);
  assign t[88] = ~(t[183]);
  assign t[89] = ~(t[184]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[115] | t[116]);
  assign t[91] = ~(t[117] | t[118]);
  assign t[92] = ~(t[119] | t[120]);
  assign t[93] = ~(t[121] & t[166]);
  assign t[94] = ~(t[122] & t[123]);
  assign t[95] = ~(t[121] & t[123]);
  assign t[96] = ~(t[122] & t[166]);
  assign t[97] = ~(t[66] | t[124]);
  assign t[98] = ~(t[66] | t[125]);
  assign t[99] = ~(t[164] | t[123]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [88:0] x;
 output y;

 wire [255:0] t;
  assign t[0] = t[1] ? t[2] : t[74];
  assign t[100] = t[126] ^ x[2];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[13];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[19];
  assign t[105] = t[131] ^ x[22];
  assign t[106] = t[132] ^ x[25];
  assign t[107] = t[133] ^ x[28];
  assign t[108] = t[134] ^ x[31];
  assign t[109] = t[135] ^ x[36];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[39];
  assign t[111] = t[137] ^ x[42];
  assign t[112] = t[138] ^ x[47];
  assign t[113] = t[139] ^ x[50];
  assign t[114] = t[140] ^ x[55];
  assign t[115] = t[141] ^ x[58];
  assign t[116] = t[142] ^ x[61];
  assign t[117] = t[143] ^ x[64];
  assign t[118] = t[144] ^ x[67];
  assign t[119] = t[145] ^ x[70];
  assign t[11] = ~(x[3]);
  assign t[120] = t[146] ^ x[73];
  assign t[121] = t[147] ^ x[76];
  assign t[122] = t[148] ^ x[79];
  assign t[123] = t[149] ^ x[82];
  assign t[124] = t[150] ^ x[85];
  assign t[125] = t[151] ^ x[88];
  assign t[126] = (t[152] & ~t[153]);
  assign t[127] = (t[154] & ~t[155]);
  assign t[128] = (t[156] & ~t[157]);
  assign t[129] = (t[158] & ~t[159]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[160] & ~t[161]);
  assign t[131] = (t[162] & ~t[163]);
  assign t[132] = (t[164] & ~t[165]);
  assign t[133] = (t[166] & ~t[167]);
  assign t[134] = (t[168] & ~t[169]);
  assign t[135] = (t[170] & ~t[171]);
  assign t[136] = (t[172] & ~t[173]);
  assign t[137] = (t[174] & ~t[175]);
  assign t[138] = (t[176] & ~t[177]);
  assign t[139] = (t[178] & ~t[179]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (t[180] & ~t[181]);
  assign t[141] = (t[182] & ~t[183]);
  assign t[142] = (t[184] & ~t[185]);
  assign t[143] = (t[186] & ~t[187]);
  assign t[144] = (t[188] & ~t[189]);
  assign t[145] = (t[190] & ~t[191]);
  assign t[146] = (t[192] & ~t[193]);
  assign t[147] = (t[194] & ~t[195]);
  assign t[148] = (t[196] & ~t[197]);
  assign t[149] = (t[198] & ~t[199]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[200] & ~t[201]);
  assign t[151] = (t[202] & ~t[203]);
  assign t[152] = t[204] ^ x[2];
  assign t[153] = t[205] ^ x[1];
  assign t[154] = t[206] ^ x[10];
  assign t[155] = t[207] ^ x[9];
  assign t[156] = t[208] ^ x[13];
  assign t[157] = t[209] ^ x[12];
  assign t[158] = t[210] ^ x[16];
  assign t[159] = t[211] ^ x[15];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[212] ^ x[19];
  assign t[161] = t[213] ^ x[18];
  assign t[162] = t[214] ^ x[22];
  assign t[163] = t[215] ^ x[21];
  assign t[164] = t[216] ^ x[25];
  assign t[165] = t[217] ^ x[24];
  assign t[166] = t[218] ^ x[28];
  assign t[167] = t[219] ^ x[27];
  assign t[168] = t[220] ^ x[31];
  assign t[169] = t[221] ^ x[30];
  assign t[16] = ~(t[75] & t[76]);
  assign t[170] = t[222] ^ x[36];
  assign t[171] = t[223] ^ x[35];
  assign t[172] = t[224] ^ x[39];
  assign t[173] = t[225] ^ x[38];
  assign t[174] = t[226] ^ x[42];
  assign t[175] = t[227] ^ x[41];
  assign t[176] = t[228] ^ x[47];
  assign t[177] = t[229] ^ x[46];
  assign t[178] = t[230] ^ x[50];
  assign t[179] = t[231] ^ x[49];
  assign t[17] = ~(t[77] & t[78]);
  assign t[180] = t[232] ^ x[55];
  assign t[181] = t[233] ^ x[54];
  assign t[182] = t[234] ^ x[58];
  assign t[183] = t[235] ^ x[57];
  assign t[184] = t[236] ^ x[61];
  assign t[185] = t[237] ^ x[60];
  assign t[186] = t[238] ^ x[64];
  assign t[187] = t[239] ^ x[63];
  assign t[188] = t[240] ^ x[67];
  assign t[189] = t[241] ^ x[66];
  assign t[18] = ~(t[24]);
  assign t[190] = t[242] ^ x[70];
  assign t[191] = t[243] ^ x[69];
  assign t[192] = t[244] ^ x[73];
  assign t[193] = t[245] ^ x[72];
  assign t[194] = t[246] ^ x[76];
  assign t[195] = t[247] ^ x[75];
  assign t[196] = t[248] ^ x[79];
  assign t[197] = t[249] ^ x[78];
  assign t[198] = t[250] ^ x[82];
  assign t[199] = t[251] ^ x[81];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[252] ^ x[85];
  assign t[201] = t[253] ^ x[84];
  assign t[202] = t[254] ^ x[88];
  assign t[203] = t[255] ^ x[87];
  assign t[204] = (x[0]);
  assign t[205] = (x[0]);
  assign t[206] = (x[8]);
  assign t[207] = (x[8]);
  assign t[208] = (x[11]);
  assign t[209] = (x[11]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[14]);
  assign t[211] = (x[14]);
  assign t[212] = (x[17]);
  assign t[213] = (x[17]);
  assign t[214] = (x[20]);
  assign t[215] = (x[20]);
  assign t[216] = (x[23]);
  assign t[217] = (x[23]);
  assign t[218] = (x[26]);
  assign t[219] = (x[26]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[29]);
  assign t[221] = (x[29]);
  assign t[222] = (x[34]);
  assign t[223] = (x[34]);
  assign t[224] = (x[37]);
  assign t[225] = (x[37]);
  assign t[226] = (x[40]);
  assign t[227] = (x[40]);
  assign t[228] = (x[45]);
  assign t[229] = (x[45]);
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = (x[48]);
  assign t[231] = (x[48]);
  assign t[232] = (x[53]);
  assign t[233] = (x[53]);
  assign t[234] = (x[56]);
  assign t[235] = (x[56]);
  assign t[236] = (x[59]);
  assign t[237] = (x[59]);
  assign t[238] = (x[62]);
  assign t[239] = (x[62]);
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[65]);
  assign t[241] = (x[65]);
  assign t[242] = (x[68]);
  assign t[243] = (x[68]);
  assign t[244] = (x[71]);
  assign t[245] = (x[71]);
  assign t[246] = (x[74]);
  assign t[247] = (x[74]);
  assign t[248] = (x[77]);
  assign t[249] = (x[77]);
  assign t[24] = ~(t[77]);
  assign t[250] = (x[80]);
  assign t[251] = (x[80]);
  assign t[252] = (x[83]);
  assign t[253] = (x[83]);
  assign t[254] = (x[86]);
  assign t[255] = (x[86]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[79] & t[37]);
  assign t[28] = ~(t[80] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[81] & t[47]);
  assign t[34] = ~(t[82] & t[48]);
  assign t[35] = t[49] ? x[33] : x[32];
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[83]);
  assign t[38] = ~(t[83] & t[52]);
  assign t[39] = ~(t[84] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[85] & t[54]);
  assign t[41] = t[55] ? x[44] : x[43];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[86] & t[58]);
  assign t[44] = ~(t[87] & t[59]);
  assign t[45] = t[49] ? x[52] : x[51];
  assign t[46] = ~(t[60] & t[61]);
  assign t[47] = ~(t[88]);
  assign t[48] = ~(t[88] & t[62]);
  assign t[49] = ~(t[24]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[90] & t[64]);
  assign t[52] = ~(t[79]);
  assign t[53] = ~(t[91]);
  assign t[54] = ~(t[91] & t[65]);
  assign t[55] = ~(t[24]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93] & t[67]);
  assign t[58] = ~(t[94]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[96] & t[70]);
  assign t[62] = ~(t[81]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[97] & t[71]);
  assign t[65] = ~(t[84]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[98] & t[72]);
  assign t[68] = ~(t[86]);
  assign t[69] = ~(t[99]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[99] & t[73]);
  assign t[71] = ~(t[89]);
  assign t[72] = ~(t[92]);
  assign t[73] = ~(t[95]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = (t[125]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind191(x, y);
 input [88:0] x;
 output y;

 wire [255:0] t;
  assign t[0] = t[1] ? t[2] : t[74];
  assign t[100] = t[126] ^ x[2];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[13];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[19];
  assign t[105] = t[131] ^ x[22];
  assign t[106] = t[132] ^ x[25];
  assign t[107] = t[133] ^ x[28];
  assign t[108] = t[134] ^ x[31];
  assign t[109] = t[135] ^ x[36];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[39];
  assign t[111] = t[137] ^ x[42];
  assign t[112] = t[138] ^ x[47];
  assign t[113] = t[139] ^ x[50];
  assign t[114] = t[140] ^ x[55];
  assign t[115] = t[141] ^ x[58];
  assign t[116] = t[142] ^ x[61];
  assign t[117] = t[143] ^ x[64];
  assign t[118] = t[144] ^ x[67];
  assign t[119] = t[145] ^ x[70];
  assign t[11] = ~(x[3]);
  assign t[120] = t[146] ^ x[73];
  assign t[121] = t[147] ^ x[76];
  assign t[122] = t[148] ^ x[79];
  assign t[123] = t[149] ^ x[82];
  assign t[124] = t[150] ^ x[85];
  assign t[125] = t[151] ^ x[88];
  assign t[126] = (t[152] & ~t[153]);
  assign t[127] = (t[154] & ~t[155]);
  assign t[128] = (t[156] & ~t[157]);
  assign t[129] = (t[158] & ~t[159]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[160] & ~t[161]);
  assign t[131] = (t[162] & ~t[163]);
  assign t[132] = (t[164] & ~t[165]);
  assign t[133] = (t[166] & ~t[167]);
  assign t[134] = (t[168] & ~t[169]);
  assign t[135] = (t[170] & ~t[171]);
  assign t[136] = (t[172] & ~t[173]);
  assign t[137] = (t[174] & ~t[175]);
  assign t[138] = (t[176] & ~t[177]);
  assign t[139] = (t[178] & ~t[179]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (t[180] & ~t[181]);
  assign t[141] = (t[182] & ~t[183]);
  assign t[142] = (t[184] & ~t[185]);
  assign t[143] = (t[186] & ~t[187]);
  assign t[144] = (t[188] & ~t[189]);
  assign t[145] = (t[190] & ~t[191]);
  assign t[146] = (t[192] & ~t[193]);
  assign t[147] = (t[194] & ~t[195]);
  assign t[148] = (t[196] & ~t[197]);
  assign t[149] = (t[198] & ~t[199]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[200] & ~t[201]);
  assign t[151] = (t[202] & ~t[203]);
  assign t[152] = t[204] ^ x[2];
  assign t[153] = t[205] ^ x[1];
  assign t[154] = t[206] ^ x[10];
  assign t[155] = t[207] ^ x[9];
  assign t[156] = t[208] ^ x[13];
  assign t[157] = t[209] ^ x[12];
  assign t[158] = t[210] ^ x[16];
  assign t[159] = t[211] ^ x[15];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[212] ^ x[19];
  assign t[161] = t[213] ^ x[18];
  assign t[162] = t[214] ^ x[22];
  assign t[163] = t[215] ^ x[21];
  assign t[164] = t[216] ^ x[25];
  assign t[165] = t[217] ^ x[24];
  assign t[166] = t[218] ^ x[28];
  assign t[167] = t[219] ^ x[27];
  assign t[168] = t[220] ^ x[31];
  assign t[169] = t[221] ^ x[30];
  assign t[16] = ~(t[75] & t[76]);
  assign t[170] = t[222] ^ x[36];
  assign t[171] = t[223] ^ x[35];
  assign t[172] = t[224] ^ x[39];
  assign t[173] = t[225] ^ x[38];
  assign t[174] = t[226] ^ x[42];
  assign t[175] = t[227] ^ x[41];
  assign t[176] = t[228] ^ x[47];
  assign t[177] = t[229] ^ x[46];
  assign t[178] = t[230] ^ x[50];
  assign t[179] = t[231] ^ x[49];
  assign t[17] = ~(t[77] & t[78]);
  assign t[180] = t[232] ^ x[55];
  assign t[181] = t[233] ^ x[54];
  assign t[182] = t[234] ^ x[58];
  assign t[183] = t[235] ^ x[57];
  assign t[184] = t[236] ^ x[61];
  assign t[185] = t[237] ^ x[60];
  assign t[186] = t[238] ^ x[64];
  assign t[187] = t[239] ^ x[63];
  assign t[188] = t[240] ^ x[67];
  assign t[189] = t[241] ^ x[66];
  assign t[18] = ~(t[24]);
  assign t[190] = t[242] ^ x[70];
  assign t[191] = t[243] ^ x[69];
  assign t[192] = t[244] ^ x[73];
  assign t[193] = t[245] ^ x[72];
  assign t[194] = t[246] ^ x[76];
  assign t[195] = t[247] ^ x[75];
  assign t[196] = t[248] ^ x[79];
  assign t[197] = t[249] ^ x[78];
  assign t[198] = t[250] ^ x[82];
  assign t[199] = t[251] ^ x[81];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[252] ^ x[85];
  assign t[201] = t[253] ^ x[84];
  assign t[202] = t[254] ^ x[88];
  assign t[203] = t[255] ^ x[87];
  assign t[204] = (x[0]);
  assign t[205] = (x[0]);
  assign t[206] = (x[8]);
  assign t[207] = (x[8]);
  assign t[208] = (x[11]);
  assign t[209] = (x[11]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[14]);
  assign t[211] = (x[14]);
  assign t[212] = (x[17]);
  assign t[213] = (x[17]);
  assign t[214] = (x[20]);
  assign t[215] = (x[20]);
  assign t[216] = (x[23]);
  assign t[217] = (x[23]);
  assign t[218] = (x[26]);
  assign t[219] = (x[26]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[29]);
  assign t[221] = (x[29]);
  assign t[222] = (x[34]);
  assign t[223] = (x[34]);
  assign t[224] = (x[37]);
  assign t[225] = (x[37]);
  assign t[226] = (x[40]);
  assign t[227] = (x[40]);
  assign t[228] = (x[45]);
  assign t[229] = (x[45]);
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = (x[48]);
  assign t[231] = (x[48]);
  assign t[232] = (x[53]);
  assign t[233] = (x[53]);
  assign t[234] = (x[56]);
  assign t[235] = (x[56]);
  assign t[236] = (x[59]);
  assign t[237] = (x[59]);
  assign t[238] = (x[62]);
  assign t[239] = (x[62]);
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[65]);
  assign t[241] = (x[65]);
  assign t[242] = (x[68]);
  assign t[243] = (x[68]);
  assign t[244] = (x[71]);
  assign t[245] = (x[71]);
  assign t[246] = (x[74]);
  assign t[247] = (x[74]);
  assign t[248] = (x[77]);
  assign t[249] = (x[77]);
  assign t[24] = ~(t[77]);
  assign t[250] = (x[80]);
  assign t[251] = (x[80]);
  assign t[252] = (x[83]);
  assign t[253] = (x[83]);
  assign t[254] = (x[86]);
  assign t[255] = (x[86]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[79] & t[37]);
  assign t[28] = ~(t[80] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[81] & t[47]);
  assign t[34] = ~(t[82] & t[48]);
  assign t[35] = t[49] ? x[33] : x[32];
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[83]);
  assign t[38] = ~(t[83] & t[52]);
  assign t[39] = ~(t[84] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[85] & t[54]);
  assign t[41] = t[55] ? x[44] : x[43];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[86] & t[58]);
  assign t[44] = ~(t[87] & t[59]);
  assign t[45] = t[49] ? x[52] : x[51];
  assign t[46] = ~(t[60] & t[61]);
  assign t[47] = ~(t[88]);
  assign t[48] = ~(t[88] & t[62]);
  assign t[49] = ~(t[24]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[90] & t[64]);
  assign t[52] = ~(t[79]);
  assign t[53] = ~(t[91]);
  assign t[54] = ~(t[91] & t[65]);
  assign t[55] = ~(t[24]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93] & t[67]);
  assign t[58] = ~(t[94]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[96] & t[70]);
  assign t[62] = ~(t[81]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[97] & t[71]);
  assign t[65] = ~(t[84]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[98] & t[72]);
  assign t[68] = ~(t[86]);
  assign t[69] = ~(t[99]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[99] & t[73]);
  assign t[71] = ~(t[89]);
  assign t[72] = ~(t[92]);
  assign t[73] = ~(t[95]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = (t[125]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [106:0] x;
 output y;

 wire [310:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[2];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[10];
  assign t[121] = t[153] ^ x[13];
  assign t[122] = t[154] ^ x[16];
  assign t[123] = t[155] ^ x[19];
  assign t[124] = t[156] ^ x[22];
  assign t[125] = t[157] ^ x[25];
  assign t[126] = t[158] ^ x[30];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[36];
  assign t[129] = t[161] ^ x[41];
  assign t[12] = t[88] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[46];
  assign t[131] = t[163] ^ x[49];
  assign t[132] = t[164] ^ x[52];
  assign t[133] = t[165] ^ x[55];
  assign t[134] = t[166] ^ x[58];
  assign t[135] = t[167] ^ x[61];
  assign t[136] = t[168] ^ x[64];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[70];
  assign t[139] = t[171] ^ x[73];
  assign t[13] = ~(t[18] ^ t[15]);
  assign t[140] = t[172] ^ x[76];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[82];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = t[176] ^ x[88];
  assign t[145] = t[177] ^ x[91];
  assign t[146] = t[178] ^ x[94];
  assign t[147] = t[179] ^ x[97];
  assign t[148] = t[180] ^ x[100];
  assign t[149] = t[181] ^ x[103];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[182] ^ x[106];
  assign t[151] = (t[183] & ~t[184]);
  assign t[152] = (t[185] & ~t[186]);
  assign t[153] = (t[187] & ~t[188]);
  assign t[154] = (t[189] & ~t[190]);
  assign t[155] = (t[191] & ~t[192]);
  assign t[156] = (t[193] & ~t[194]);
  assign t[157] = (t[195] & ~t[196]);
  assign t[158] = (t[197] & ~t[198]);
  assign t[159] = (t[199] & ~t[200]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[201] & ~t[202]);
  assign t[161] = (t[203] & ~t[204]);
  assign t[162] = (t[205] & ~t[206]);
  assign t[163] = (t[207] & ~t[208]);
  assign t[164] = (t[209] & ~t[210]);
  assign t[165] = (t[211] & ~t[212]);
  assign t[166] = (t[213] & ~t[214]);
  assign t[167] = (t[215] & ~t[216]);
  assign t[168] = (t[217] & ~t[218]);
  assign t[169] = (t[219] & ~t[220]);
  assign t[16] = ~(t[89] & t[90]);
  assign t[170] = (t[221] & ~t[222]);
  assign t[171] = (t[223] & ~t[224]);
  assign t[172] = (t[225] & ~t[226]);
  assign t[173] = (t[227] & ~t[228]);
  assign t[174] = (t[229] & ~t[230]);
  assign t[175] = (t[231] & ~t[232]);
  assign t[176] = (t[233] & ~t[234]);
  assign t[177] = (t[235] & ~t[236]);
  assign t[178] = (t[237] & ~t[238]);
  assign t[179] = (t[239] & ~t[240]);
  assign t[17] = ~(t[88] & t[91]);
  assign t[180] = (t[241] & ~t[242]);
  assign t[181] = (t[243] & ~t[244]);
  assign t[182] = (t[245] & ~t[246]);
  assign t[183] = t[247] ^ x[2];
  assign t[184] = t[248] ^ x[1];
  assign t[185] = t[249] ^ x[10];
  assign t[186] = t[250] ^ x[9];
  assign t[187] = t[251] ^ x[13];
  assign t[188] = t[252] ^ x[12];
  assign t[189] = t[253] ^ x[16];
  assign t[18] = x[4] ? t[24] : t[23];
  assign t[190] = t[254] ^ x[15];
  assign t[191] = t[255] ^ x[19];
  assign t[192] = t[256] ^ x[18];
  assign t[193] = t[257] ^ x[22];
  assign t[194] = t[258] ^ x[21];
  assign t[195] = t[259] ^ x[25];
  assign t[196] = t[260] ^ x[24];
  assign t[197] = t[261] ^ x[30];
  assign t[198] = t[262] ^ x[29];
  assign t[199] = t[263] ^ x[33];
  assign t[19] = ~(t[25] & t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[32];
  assign t[201] = t[265] ^ x[36];
  assign t[202] = t[266] ^ x[35];
  assign t[203] = t[267] ^ x[41];
  assign t[204] = t[268] ^ x[40];
  assign t[205] = t[269] ^ x[46];
  assign t[206] = t[270] ^ x[45];
  assign t[207] = t[271] ^ x[49];
  assign t[208] = t[272] ^ x[48];
  assign t[209] = t[273] ^ x[52];
  assign t[20] = t[12] ^ t[23];
  assign t[210] = t[274] ^ x[51];
  assign t[211] = t[275] ^ x[55];
  assign t[212] = t[276] ^ x[54];
  assign t[213] = t[277] ^ x[58];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[61];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[64];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[67];
  assign t[21] = x[4] ? t[28] : t[27];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[70];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[73];
  assign t[224] = t[288] ^ x[72];
  assign t[225] = t[289] ^ x[76];
  assign t[226] = t[290] ^ x[75];
  assign t[227] = t[291] ^ x[79];
  assign t[228] = t[292] ^ x[78];
  assign t[229] = t[293] ^ x[82];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[81];
  assign t[231] = t[295] ^ x[85];
  assign t[232] = t[296] ^ x[84];
  assign t[233] = t[297] ^ x[88];
  assign t[234] = t[298] ^ x[87];
  assign t[235] = t[299] ^ x[91];
  assign t[236] = t[300] ^ x[90];
  assign t[237] = t[301] ^ x[94];
  assign t[238] = t[302] ^ x[93];
  assign t[239] = t[303] ^ x[97];
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = t[304] ^ x[96];
  assign t[241] = t[305] ^ x[100];
  assign t[242] = t[306] ^ x[99];
  assign t[243] = t[307] ^ x[103];
  assign t[244] = t[308] ^ x[102];
  assign t[245] = t[309] ^ x[106];
  assign t[246] = t[310] ^ x[105];
  assign t[247] = (x[0]);
  assign t[248] = (x[0]);
  assign t[249] = (x[8]);
  assign t[24] = t[33] ^ t[34];
  assign t[250] = (x[8]);
  assign t[251] = (x[11]);
  assign t[252] = (x[11]);
  assign t[253] = (x[14]);
  assign t[254] = (x[14]);
  assign t[255] = (x[17]);
  assign t[256] = (x[17]);
  assign t[257] = (x[20]);
  assign t[258] = (x[20]);
  assign t[259] = (x[23]);
  assign t[25] = ~(t[35] & t[36]);
  assign t[260] = (x[23]);
  assign t[261] = (x[28]);
  assign t[262] = (x[28]);
  assign t[263] = (x[31]);
  assign t[264] = (x[31]);
  assign t[265] = (x[34]);
  assign t[266] = (x[34]);
  assign t[267] = (x[39]);
  assign t[268] = (x[39]);
  assign t[269] = (x[44]);
  assign t[26] = ~(t[37] & t[92]);
  assign t[270] = (x[44]);
  assign t[271] = (x[47]);
  assign t[272] = (x[47]);
  assign t[273] = (x[50]);
  assign t[274] = (x[50]);
  assign t[275] = (x[53]);
  assign t[276] = (x[53]);
  assign t[277] = (x[56]);
  assign t[278] = (x[56]);
  assign t[279] = (x[59]);
  assign t[27] = ~(t[38] & t[39]);
  assign t[280] = (x[59]);
  assign t[281] = (x[62]);
  assign t[282] = (x[62]);
  assign t[283] = (x[65]);
  assign t[284] = (x[65]);
  assign t[285] = (x[68]);
  assign t[286] = (x[68]);
  assign t[287] = (x[71]);
  assign t[288] = (x[71]);
  assign t[289] = (x[74]);
  assign t[28] = t[40] ^ t[41];
  assign t[290] = (x[74]);
  assign t[291] = (x[77]);
  assign t[292] = (x[77]);
  assign t[293] = (x[80]);
  assign t[294] = (x[80]);
  assign t[295] = (x[83]);
  assign t[296] = (x[83]);
  assign t[297] = (x[86]);
  assign t[298] = (x[86]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[42] & t[43]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[89]);
  assign t[301] = (x[92]);
  assign t[302] = (x[92]);
  assign t[303] = (x[95]);
  assign t[304] = (x[95]);
  assign t[305] = (x[98]);
  assign t[306] = (x[98]);
  assign t[307] = (x[101]);
  assign t[308] = (x[101]);
  assign t[309] = (x[104]);
  assign t[30] = t[44] ^ t[45];
  assign t[310] = (x[104]);
  assign t[31] = ~(t[46] & t[47]);
  assign t[32] = ~(t[48] & t[93]);
  assign t[33] = t[49] ? x[27] : x[26];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = ~(t[94]);
  assign t[36] = ~(t[95]);
  assign t[37] = ~(t[52] & t[53]);
  assign t[38] = ~(t[54] & t[55]);
  assign t[39] = ~(t[56] & t[96]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[49] ? x[38] : x[37];
  assign t[41] = ~(t[57] & t[58]);
  assign t[42] = ~(t[59] & t[60]);
  assign t[43] = ~(t[61] & t[97]);
  assign t[44] = t[62] ? x[43] : x[42];
  assign t[45] = ~(t[63] & t[64]);
  assign t[46] = ~(t[98]);
  assign t[47] = ~(t[99]);
  assign t[48] = ~(t[65] & t[66]);
  assign t[49] = ~(t[67]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[70] & t[100]);
  assign t[52] = ~(t[95] & t[94]);
  assign t[53] = ~(t[101]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(t[103]);
  assign t[56] = ~(t[71] & t[72]);
  assign t[57] = ~(t[73] & t[74]);
  assign t[58] = ~(t[75] & t[104]);
  assign t[59] = ~(t[105]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[106]);
  assign t[61] = ~(t[76] & t[77]);
  assign t[62] = ~(t[67]);
  assign t[63] = ~(t[78] & t[79]);
  assign t[64] = ~(t[80] & t[107]);
  assign t[65] = ~(t[99] & t[98]);
  assign t[66] = ~(t[87]);
  assign t[67] = ~(t[88]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [106:0] x;
 output y;

 wire [310:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[2];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[10];
  assign t[121] = t[153] ^ x[13];
  assign t[122] = t[154] ^ x[16];
  assign t[123] = t[155] ^ x[19];
  assign t[124] = t[156] ^ x[22];
  assign t[125] = t[157] ^ x[25];
  assign t[126] = t[158] ^ x[30];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[36];
  assign t[129] = t[161] ^ x[41];
  assign t[12] = t[88] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[46];
  assign t[131] = t[163] ^ x[49];
  assign t[132] = t[164] ^ x[52];
  assign t[133] = t[165] ^ x[55];
  assign t[134] = t[166] ^ x[58];
  assign t[135] = t[167] ^ x[61];
  assign t[136] = t[168] ^ x[64];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[70];
  assign t[139] = t[171] ^ x[73];
  assign t[13] = ~(t[18] ^ t[15]);
  assign t[140] = t[172] ^ x[76];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[82];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = t[176] ^ x[88];
  assign t[145] = t[177] ^ x[91];
  assign t[146] = t[178] ^ x[94];
  assign t[147] = t[179] ^ x[97];
  assign t[148] = t[180] ^ x[100];
  assign t[149] = t[181] ^ x[103];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[182] ^ x[106];
  assign t[151] = (t[183] & ~t[184]);
  assign t[152] = (t[185] & ~t[186]);
  assign t[153] = (t[187] & ~t[188]);
  assign t[154] = (t[189] & ~t[190]);
  assign t[155] = (t[191] & ~t[192]);
  assign t[156] = (t[193] & ~t[194]);
  assign t[157] = (t[195] & ~t[196]);
  assign t[158] = (t[197] & ~t[198]);
  assign t[159] = (t[199] & ~t[200]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[201] & ~t[202]);
  assign t[161] = (t[203] & ~t[204]);
  assign t[162] = (t[205] & ~t[206]);
  assign t[163] = (t[207] & ~t[208]);
  assign t[164] = (t[209] & ~t[210]);
  assign t[165] = (t[211] & ~t[212]);
  assign t[166] = (t[213] & ~t[214]);
  assign t[167] = (t[215] & ~t[216]);
  assign t[168] = (t[217] & ~t[218]);
  assign t[169] = (t[219] & ~t[220]);
  assign t[16] = ~(t[89] & t[90]);
  assign t[170] = (t[221] & ~t[222]);
  assign t[171] = (t[223] & ~t[224]);
  assign t[172] = (t[225] & ~t[226]);
  assign t[173] = (t[227] & ~t[228]);
  assign t[174] = (t[229] & ~t[230]);
  assign t[175] = (t[231] & ~t[232]);
  assign t[176] = (t[233] & ~t[234]);
  assign t[177] = (t[235] & ~t[236]);
  assign t[178] = (t[237] & ~t[238]);
  assign t[179] = (t[239] & ~t[240]);
  assign t[17] = ~(t[88] & t[91]);
  assign t[180] = (t[241] & ~t[242]);
  assign t[181] = (t[243] & ~t[244]);
  assign t[182] = (t[245] & ~t[246]);
  assign t[183] = t[247] ^ x[2];
  assign t[184] = t[248] ^ x[1];
  assign t[185] = t[249] ^ x[10];
  assign t[186] = t[250] ^ x[9];
  assign t[187] = t[251] ^ x[13];
  assign t[188] = t[252] ^ x[12];
  assign t[189] = t[253] ^ x[16];
  assign t[18] = x[4] ? t[24] : t[23];
  assign t[190] = t[254] ^ x[15];
  assign t[191] = t[255] ^ x[19];
  assign t[192] = t[256] ^ x[18];
  assign t[193] = t[257] ^ x[22];
  assign t[194] = t[258] ^ x[21];
  assign t[195] = t[259] ^ x[25];
  assign t[196] = t[260] ^ x[24];
  assign t[197] = t[261] ^ x[30];
  assign t[198] = t[262] ^ x[29];
  assign t[199] = t[263] ^ x[33];
  assign t[19] = ~(t[25] & t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[32];
  assign t[201] = t[265] ^ x[36];
  assign t[202] = t[266] ^ x[35];
  assign t[203] = t[267] ^ x[41];
  assign t[204] = t[268] ^ x[40];
  assign t[205] = t[269] ^ x[46];
  assign t[206] = t[270] ^ x[45];
  assign t[207] = t[271] ^ x[49];
  assign t[208] = t[272] ^ x[48];
  assign t[209] = t[273] ^ x[52];
  assign t[20] = t[12] ^ t[23];
  assign t[210] = t[274] ^ x[51];
  assign t[211] = t[275] ^ x[55];
  assign t[212] = t[276] ^ x[54];
  assign t[213] = t[277] ^ x[58];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[61];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[64];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[67];
  assign t[21] = x[4] ? t[28] : t[27];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[70];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[73];
  assign t[224] = t[288] ^ x[72];
  assign t[225] = t[289] ^ x[76];
  assign t[226] = t[290] ^ x[75];
  assign t[227] = t[291] ^ x[79];
  assign t[228] = t[292] ^ x[78];
  assign t[229] = t[293] ^ x[82];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[81];
  assign t[231] = t[295] ^ x[85];
  assign t[232] = t[296] ^ x[84];
  assign t[233] = t[297] ^ x[88];
  assign t[234] = t[298] ^ x[87];
  assign t[235] = t[299] ^ x[91];
  assign t[236] = t[300] ^ x[90];
  assign t[237] = t[301] ^ x[94];
  assign t[238] = t[302] ^ x[93];
  assign t[239] = t[303] ^ x[97];
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = t[304] ^ x[96];
  assign t[241] = t[305] ^ x[100];
  assign t[242] = t[306] ^ x[99];
  assign t[243] = t[307] ^ x[103];
  assign t[244] = t[308] ^ x[102];
  assign t[245] = t[309] ^ x[106];
  assign t[246] = t[310] ^ x[105];
  assign t[247] = (x[0]);
  assign t[248] = (x[0]);
  assign t[249] = (x[8]);
  assign t[24] = t[33] ^ t[34];
  assign t[250] = (x[8]);
  assign t[251] = (x[11]);
  assign t[252] = (x[11]);
  assign t[253] = (x[14]);
  assign t[254] = (x[14]);
  assign t[255] = (x[17]);
  assign t[256] = (x[17]);
  assign t[257] = (x[20]);
  assign t[258] = (x[20]);
  assign t[259] = (x[23]);
  assign t[25] = ~(t[35] & t[36]);
  assign t[260] = (x[23]);
  assign t[261] = (x[28]);
  assign t[262] = (x[28]);
  assign t[263] = (x[31]);
  assign t[264] = (x[31]);
  assign t[265] = (x[34]);
  assign t[266] = (x[34]);
  assign t[267] = (x[39]);
  assign t[268] = (x[39]);
  assign t[269] = (x[44]);
  assign t[26] = ~(t[37] & t[92]);
  assign t[270] = (x[44]);
  assign t[271] = (x[47]);
  assign t[272] = (x[47]);
  assign t[273] = (x[50]);
  assign t[274] = (x[50]);
  assign t[275] = (x[53]);
  assign t[276] = (x[53]);
  assign t[277] = (x[56]);
  assign t[278] = (x[56]);
  assign t[279] = (x[59]);
  assign t[27] = ~(t[38] & t[39]);
  assign t[280] = (x[59]);
  assign t[281] = (x[62]);
  assign t[282] = (x[62]);
  assign t[283] = (x[65]);
  assign t[284] = (x[65]);
  assign t[285] = (x[68]);
  assign t[286] = (x[68]);
  assign t[287] = (x[71]);
  assign t[288] = (x[71]);
  assign t[289] = (x[74]);
  assign t[28] = t[40] ^ t[41];
  assign t[290] = (x[74]);
  assign t[291] = (x[77]);
  assign t[292] = (x[77]);
  assign t[293] = (x[80]);
  assign t[294] = (x[80]);
  assign t[295] = (x[83]);
  assign t[296] = (x[83]);
  assign t[297] = (x[86]);
  assign t[298] = (x[86]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[42] & t[43]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[89]);
  assign t[301] = (x[92]);
  assign t[302] = (x[92]);
  assign t[303] = (x[95]);
  assign t[304] = (x[95]);
  assign t[305] = (x[98]);
  assign t[306] = (x[98]);
  assign t[307] = (x[101]);
  assign t[308] = (x[101]);
  assign t[309] = (x[104]);
  assign t[30] = t[44] ^ t[45];
  assign t[310] = (x[104]);
  assign t[31] = ~(t[46] & t[47]);
  assign t[32] = ~(t[48] & t[93]);
  assign t[33] = t[49] ? x[27] : x[26];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = ~(t[94]);
  assign t[36] = ~(t[95]);
  assign t[37] = ~(t[52] & t[53]);
  assign t[38] = ~(t[54] & t[55]);
  assign t[39] = ~(t[56] & t[96]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[49] ? x[38] : x[37];
  assign t[41] = ~(t[57] & t[58]);
  assign t[42] = ~(t[59] & t[60]);
  assign t[43] = ~(t[61] & t[97]);
  assign t[44] = t[62] ? x[43] : x[42];
  assign t[45] = ~(t[63] & t[64]);
  assign t[46] = ~(t[98]);
  assign t[47] = ~(t[99]);
  assign t[48] = ~(t[65] & t[66]);
  assign t[49] = ~(t[67]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[70] & t[100]);
  assign t[52] = ~(t[95] & t[94]);
  assign t[53] = ~(t[101]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(t[103]);
  assign t[56] = ~(t[71] & t[72]);
  assign t[57] = ~(t[73] & t[74]);
  assign t[58] = ~(t[75] & t[104]);
  assign t[59] = ~(t[105]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[106]);
  assign t[61] = ~(t[76] & t[77]);
  assign t[62] = ~(t[67]);
  assign t[63] = ~(t[78] & t[79]);
  assign t[64] = ~(t[80] & t[107]);
  assign t[65] = ~(t[99] & t[98]);
  assign t[66] = ~(t[87]);
  assign t[67] = ~(t[88]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [106:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[2];
  assign t[113] = t[145] ^ x[10];
  assign t[114] = t[146] ^ x[13];
  assign t[115] = t[147] ^ x[16];
  assign t[116] = t[148] ^ x[19];
  assign t[117] = t[149] ^ x[22];
  assign t[118] = t[150] ^ x[25];
  assign t[119] = t[151] ^ x[30];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[36];
  assign t[122] = t[154] ^ x[41];
  assign t[123] = t[155] ^ x[46];
  assign t[124] = t[156] ^ x[49];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[55];
  assign t[127] = t[159] ^ x[58];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[70];
  assign t[132] = t[164] ^ x[73];
  assign t[133] = t[165] ^ x[76];
  assign t[134] = t[166] ^ x[79];
  assign t[135] = t[167] ^ x[82];
  assign t[136] = t[168] ^ x[85];
  assign t[137] = t[169] ^ x[88];
  assign t[138] = t[170] ^ x[91];
  assign t[139] = t[171] ^ x[94];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[97];
  assign t[141] = t[173] ^ x[100];
  assign t[142] = t[174] ^ x[103];
  assign t[143] = t[175] ^ x[106];
  assign t[144] = (t[176] & ~t[177]);
  assign t[145] = (t[178] & ~t[179]);
  assign t[146] = (t[180] & ~t[181]);
  assign t[147] = (t[182] & ~t[183]);
  assign t[148] = (t[184] & ~t[185]);
  assign t[149] = (t[186] & ~t[187]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[188] & ~t[189]);
  assign t[151] = (t[190] & ~t[191]);
  assign t[152] = (t[192] & ~t[193]);
  assign t[153] = (t[194] & ~t[195]);
  assign t[154] = (t[196] & ~t[197]);
  assign t[155] = (t[198] & ~t[199]);
  assign t[156] = (t[200] & ~t[201]);
  assign t[157] = (t[202] & ~t[203]);
  assign t[158] = (t[204] & ~t[205]);
  assign t[159] = (t[206] & ~t[207]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[208] & ~t[209]);
  assign t[161] = (t[210] & ~t[211]);
  assign t[162] = (t[212] & ~t[213]);
  assign t[163] = (t[214] & ~t[215]);
  assign t[164] = (t[216] & ~t[217]);
  assign t[165] = (t[218] & ~t[219]);
  assign t[166] = (t[220] & ~t[221]);
  assign t[167] = (t[222] & ~t[223]);
  assign t[168] = (t[224] & ~t[225]);
  assign t[169] = (t[226] & ~t[227]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (t[228] & ~t[229]);
  assign t[171] = (t[230] & ~t[231]);
  assign t[172] = (t[232] & ~t[233]);
  assign t[173] = (t[234] & ~t[235]);
  assign t[174] = (t[236] & ~t[237]);
  assign t[175] = (t[238] & ~t[239]);
  assign t[176] = t[240] ^ x[2];
  assign t[177] = t[241] ^ x[1];
  assign t[178] = t[242] ^ x[10];
  assign t[179] = t[243] ^ x[9];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[244] ^ x[13];
  assign t[181] = t[245] ^ x[12];
  assign t[182] = t[246] ^ x[16];
  assign t[183] = t[247] ^ x[15];
  assign t[184] = t[248] ^ x[19];
  assign t[185] = t[249] ^ x[18];
  assign t[186] = t[250] ^ x[22];
  assign t[187] = t[251] ^ x[21];
  assign t[188] = t[252] ^ x[25];
  assign t[189] = t[253] ^ x[24];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[30];
  assign t[191] = t[255] ^ x[29];
  assign t[192] = t[256] ^ x[33];
  assign t[193] = t[257] ^ x[32];
  assign t[194] = t[258] ^ x[36];
  assign t[195] = t[259] ^ x[35];
  assign t[196] = t[260] ^ x[41];
  assign t[197] = t[261] ^ x[40];
  assign t[198] = t[262] ^ x[46];
  assign t[199] = t[263] ^ x[45];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[49];
  assign t[201] = t[265] ^ x[48];
  assign t[202] = t[266] ^ x[52];
  assign t[203] = t[267] ^ x[51];
  assign t[204] = t[268] ^ x[55];
  assign t[205] = t[269] ^ x[54];
  assign t[206] = t[270] ^ x[58];
  assign t[207] = t[271] ^ x[57];
  assign t[208] = t[272] ^ x[61];
  assign t[209] = t[273] ^ x[60];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[64];
  assign t[211] = t[275] ^ x[63];
  assign t[212] = t[276] ^ x[67];
  assign t[213] = t[277] ^ x[66];
  assign t[214] = t[278] ^ x[70];
  assign t[215] = t[279] ^ x[69];
  assign t[216] = t[280] ^ x[73];
  assign t[217] = t[281] ^ x[72];
  assign t[218] = t[282] ^ x[76];
  assign t[219] = t[283] ^ x[75];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[79];
  assign t[221] = t[285] ^ x[78];
  assign t[222] = t[286] ^ x[82];
  assign t[223] = t[287] ^ x[81];
  assign t[224] = t[288] ^ x[85];
  assign t[225] = t[289] ^ x[84];
  assign t[226] = t[290] ^ x[88];
  assign t[227] = t[291] ^ x[87];
  assign t[228] = t[292] ^ x[91];
  assign t[229] = t[293] ^ x[90];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[94];
  assign t[231] = t[295] ^ x[93];
  assign t[232] = t[296] ^ x[97];
  assign t[233] = t[297] ^ x[96];
  assign t[234] = t[298] ^ x[100];
  assign t[235] = t[299] ^ x[99];
  assign t[236] = t[300] ^ x[103];
  assign t[237] = t[301] ^ x[102];
  assign t[238] = t[302] ^ x[106];
  assign t[239] = t[303] ^ x[105];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[0]);
  assign t[241] = (x[0]);
  assign t[242] = (x[8]);
  assign t[243] = (x[8]);
  assign t[244] = (x[11]);
  assign t[245] = (x[11]);
  assign t[246] = (x[14]);
  assign t[247] = (x[14]);
  assign t[248] = (x[17]);
  assign t[249] = (x[17]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[20]);
  assign t[251] = (x[20]);
  assign t[252] = (x[23]);
  assign t[253] = (x[23]);
  assign t[254] = (x[28]);
  assign t[255] = (x[28]);
  assign t[256] = (x[31]);
  assign t[257] = (x[31]);
  assign t[258] = (x[34]);
  assign t[259] = (x[34]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[39]);
  assign t[261] = (x[39]);
  assign t[262] = (x[44]);
  assign t[263] = (x[44]);
  assign t[264] = (x[47]);
  assign t[265] = (x[47]);
  assign t[266] = (x[50]);
  assign t[267] = (x[50]);
  assign t[268] = (x[53]);
  assign t[269] = (x[53]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[56]);
  assign t[271] = (x[56]);
  assign t[272] = (x[59]);
  assign t[273] = (x[59]);
  assign t[274] = (x[62]);
  assign t[275] = (x[62]);
  assign t[276] = (x[65]);
  assign t[277] = (x[65]);
  assign t[278] = (x[68]);
  assign t[279] = (x[68]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[71]);
  assign t[281] = (x[71]);
  assign t[282] = (x[74]);
  assign t[283] = (x[74]);
  assign t[284] = (x[77]);
  assign t[285] = (x[77]);
  assign t[286] = (x[80]);
  assign t[287] = (x[80]);
  assign t[288] = (x[83]);
  assign t[289] = (x[83]);
  assign t[28] = t[39] | t[85];
  assign t[290] = (x[86]);
  assign t[291] = (x[86]);
  assign t[292] = (x[89]);
  assign t[293] = (x[89]);
  assign t[294] = (x[92]);
  assign t[295] = (x[92]);
  assign t[296] = (x[95]);
  assign t[297] = (x[95]);
  assign t[298] = (x[98]);
  assign t[299] = (x[98]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[101]);
  assign t[301] = (x[101]);
  assign t[302] = (x[104]);
  assign t[303] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[18] ? x[38] : x[37];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[59] & t[60]);
  assign t[45] = t[61] | t[90];
  assign t[46] = t[62] ? x[43] : x[42];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[70] & t[71]);
  assign t[58] = t[72] | t[96];
  assign t[59] = ~(t[97]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[98]);
  assign t[61] = ~(t[73] | t[59]);
  assign t[62] = ~(t[24]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [106:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[2];
  assign t[113] = t[145] ^ x[10];
  assign t[114] = t[146] ^ x[13];
  assign t[115] = t[147] ^ x[16];
  assign t[116] = t[148] ^ x[19];
  assign t[117] = t[149] ^ x[22];
  assign t[118] = t[150] ^ x[25];
  assign t[119] = t[151] ^ x[30];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[36];
  assign t[122] = t[154] ^ x[41];
  assign t[123] = t[155] ^ x[46];
  assign t[124] = t[156] ^ x[49];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[55];
  assign t[127] = t[159] ^ x[58];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[70];
  assign t[132] = t[164] ^ x[73];
  assign t[133] = t[165] ^ x[76];
  assign t[134] = t[166] ^ x[79];
  assign t[135] = t[167] ^ x[82];
  assign t[136] = t[168] ^ x[85];
  assign t[137] = t[169] ^ x[88];
  assign t[138] = t[170] ^ x[91];
  assign t[139] = t[171] ^ x[94];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[97];
  assign t[141] = t[173] ^ x[100];
  assign t[142] = t[174] ^ x[103];
  assign t[143] = t[175] ^ x[106];
  assign t[144] = (t[176] & ~t[177]);
  assign t[145] = (t[178] & ~t[179]);
  assign t[146] = (t[180] & ~t[181]);
  assign t[147] = (t[182] & ~t[183]);
  assign t[148] = (t[184] & ~t[185]);
  assign t[149] = (t[186] & ~t[187]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[188] & ~t[189]);
  assign t[151] = (t[190] & ~t[191]);
  assign t[152] = (t[192] & ~t[193]);
  assign t[153] = (t[194] & ~t[195]);
  assign t[154] = (t[196] & ~t[197]);
  assign t[155] = (t[198] & ~t[199]);
  assign t[156] = (t[200] & ~t[201]);
  assign t[157] = (t[202] & ~t[203]);
  assign t[158] = (t[204] & ~t[205]);
  assign t[159] = (t[206] & ~t[207]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[208] & ~t[209]);
  assign t[161] = (t[210] & ~t[211]);
  assign t[162] = (t[212] & ~t[213]);
  assign t[163] = (t[214] & ~t[215]);
  assign t[164] = (t[216] & ~t[217]);
  assign t[165] = (t[218] & ~t[219]);
  assign t[166] = (t[220] & ~t[221]);
  assign t[167] = (t[222] & ~t[223]);
  assign t[168] = (t[224] & ~t[225]);
  assign t[169] = (t[226] & ~t[227]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (t[228] & ~t[229]);
  assign t[171] = (t[230] & ~t[231]);
  assign t[172] = (t[232] & ~t[233]);
  assign t[173] = (t[234] & ~t[235]);
  assign t[174] = (t[236] & ~t[237]);
  assign t[175] = (t[238] & ~t[239]);
  assign t[176] = t[240] ^ x[2];
  assign t[177] = t[241] ^ x[1];
  assign t[178] = t[242] ^ x[10];
  assign t[179] = t[243] ^ x[9];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[244] ^ x[13];
  assign t[181] = t[245] ^ x[12];
  assign t[182] = t[246] ^ x[16];
  assign t[183] = t[247] ^ x[15];
  assign t[184] = t[248] ^ x[19];
  assign t[185] = t[249] ^ x[18];
  assign t[186] = t[250] ^ x[22];
  assign t[187] = t[251] ^ x[21];
  assign t[188] = t[252] ^ x[25];
  assign t[189] = t[253] ^ x[24];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[30];
  assign t[191] = t[255] ^ x[29];
  assign t[192] = t[256] ^ x[33];
  assign t[193] = t[257] ^ x[32];
  assign t[194] = t[258] ^ x[36];
  assign t[195] = t[259] ^ x[35];
  assign t[196] = t[260] ^ x[41];
  assign t[197] = t[261] ^ x[40];
  assign t[198] = t[262] ^ x[46];
  assign t[199] = t[263] ^ x[45];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[49];
  assign t[201] = t[265] ^ x[48];
  assign t[202] = t[266] ^ x[52];
  assign t[203] = t[267] ^ x[51];
  assign t[204] = t[268] ^ x[55];
  assign t[205] = t[269] ^ x[54];
  assign t[206] = t[270] ^ x[58];
  assign t[207] = t[271] ^ x[57];
  assign t[208] = t[272] ^ x[61];
  assign t[209] = t[273] ^ x[60];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[64];
  assign t[211] = t[275] ^ x[63];
  assign t[212] = t[276] ^ x[67];
  assign t[213] = t[277] ^ x[66];
  assign t[214] = t[278] ^ x[70];
  assign t[215] = t[279] ^ x[69];
  assign t[216] = t[280] ^ x[73];
  assign t[217] = t[281] ^ x[72];
  assign t[218] = t[282] ^ x[76];
  assign t[219] = t[283] ^ x[75];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[79];
  assign t[221] = t[285] ^ x[78];
  assign t[222] = t[286] ^ x[82];
  assign t[223] = t[287] ^ x[81];
  assign t[224] = t[288] ^ x[85];
  assign t[225] = t[289] ^ x[84];
  assign t[226] = t[290] ^ x[88];
  assign t[227] = t[291] ^ x[87];
  assign t[228] = t[292] ^ x[91];
  assign t[229] = t[293] ^ x[90];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[94];
  assign t[231] = t[295] ^ x[93];
  assign t[232] = t[296] ^ x[97];
  assign t[233] = t[297] ^ x[96];
  assign t[234] = t[298] ^ x[100];
  assign t[235] = t[299] ^ x[99];
  assign t[236] = t[300] ^ x[103];
  assign t[237] = t[301] ^ x[102];
  assign t[238] = t[302] ^ x[106];
  assign t[239] = t[303] ^ x[105];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[0]);
  assign t[241] = (x[0]);
  assign t[242] = (x[8]);
  assign t[243] = (x[8]);
  assign t[244] = (x[11]);
  assign t[245] = (x[11]);
  assign t[246] = (x[14]);
  assign t[247] = (x[14]);
  assign t[248] = (x[17]);
  assign t[249] = (x[17]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[20]);
  assign t[251] = (x[20]);
  assign t[252] = (x[23]);
  assign t[253] = (x[23]);
  assign t[254] = (x[28]);
  assign t[255] = (x[28]);
  assign t[256] = (x[31]);
  assign t[257] = (x[31]);
  assign t[258] = (x[34]);
  assign t[259] = (x[34]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[39]);
  assign t[261] = (x[39]);
  assign t[262] = (x[44]);
  assign t[263] = (x[44]);
  assign t[264] = (x[47]);
  assign t[265] = (x[47]);
  assign t[266] = (x[50]);
  assign t[267] = (x[50]);
  assign t[268] = (x[53]);
  assign t[269] = (x[53]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[56]);
  assign t[271] = (x[56]);
  assign t[272] = (x[59]);
  assign t[273] = (x[59]);
  assign t[274] = (x[62]);
  assign t[275] = (x[62]);
  assign t[276] = (x[65]);
  assign t[277] = (x[65]);
  assign t[278] = (x[68]);
  assign t[279] = (x[68]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[71]);
  assign t[281] = (x[71]);
  assign t[282] = (x[74]);
  assign t[283] = (x[74]);
  assign t[284] = (x[77]);
  assign t[285] = (x[77]);
  assign t[286] = (x[80]);
  assign t[287] = (x[80]);
  assign t[288] = (x[83]);
  assign t[289] = (x[83]);
  assign t[28] = t[39] | t[85];
  assign t[290] = (x[86]);
  assign t[291] = (x[86]);
  assign t[292] = (x[89]);
  assign t[293] = (x[89]);
  assign t[294] = (x[92]);
  assign t[295] = (x[92]);
  assign t[296] = (x[95]);
  assign t[297] = (x[95]);
  assign t[298] = (x[98]);
  assign t[299] = (x[98]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[101]);
  assign t[301] = (x[101]);
  assign t[302] = (x[104]);
  assign t[303] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[18] ? x[38] : x[37];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[59] & t[60]);
  assign t[45] = t[61] | t[90];
  assign t[46] = t[62] ? x[43] : x[42];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[70] & t[71]);
  assign t[58] = t[72] | t[96];
  assign t[59] = ~(t[97]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[98]);
  assign t[61] = ~(t[73] | t[59]);
  assign t[62] = ~(t[24]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind196(x, y);
 input [151:0] x;
 output y;

 wire [526:0] t;
  assign t[0] = t[1] ? t[2] : t[212];
  assign t[100] = ~(t[147] & t[148]);
  assign t[101] = ~(t[234]);
  assign t[102] = ~(t[235]);
  assign t[103] = ~(t[149] | t[150]);
  assign t[104] = t[215] ? x[84] : x[83];
  assign t[105] = t[151] | t[152];
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[224] | t[225]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[153] | t[154]);
  assign t[111] = ~(t[140] | t[155]);
  assign t[112] = ~(t[156] | t[85]);
  assign t[113] = ~(t[239]);
  assign t[114] = ~(t[240]);
  assign t[115] = ~(t[157] | t[158]);
  assign t[116] = ~(t[159] | t[160]);
  assign t[117] = ~(t[241] | t[161]);
  assign t[118] = t[30] ? x[104] : x[103];
  assign t[119] = ~(t[162] & t[163]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[243]);
  assign t[122] = ~(t[164] | t[165]);
  assign t[123] = ~(t[166] | t[167]);
  assign t[124] = ~(t[244] | t[168]);
  assign t[125] = t[30] ? x[115] : x[114];
  assign t[126] = ~(t[169] & t[170]);
  assign t[127] = ~(t[215]);
  assign t[128] = ~(t[171] & t[172]);
  assign t[129] = ~(t[173] & t[216]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[216] & t[174]);
  assign t[131] = ~(x[4] & t[175]);
  assign t[132] = ~(t[176] | t[142]);
  assign t[133] = ~(t[177] & t[178]);
  assign t[134] = t[213] ? t[130] : t[131];
  assign t[135] = ~(t[179]);
  assign t[136] = ~(t[82] | t[180]);
  assign t[137] = t[213] ? t[131] : t[181];
  assign t[138] = ~(t[245]);
  assign t[139] = ~(t[230] | t[231]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[82] | t[182]);
  assign t[141] = ~(t[31] & t[183]);
  assign t[142] = ~(t[127] | t[184]);
  assign t[143] = t[155] | t[135];
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[232] | t[233]);
  assign t[146] = ~(t[49]);
  assign t[147] = ~(t[151] | t[185]);
  assign t[148] = ~(t[140]);
  assign t[149] = ~(t[247]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[234] | t[235]);
  assign t[151] = ~(t[179] & t[133]);
  assign t[152] = ~(t[111] & t[186]);
  assign t[153] = ~(t[248]);
  assign t[154] = ~(t[237] | t[238]);
  assign t[155] = ~(t[82] | t[187]);
  assign t[156] = ~(t[127] | t[188]);
  assign t[157] = ~(t[249]);
  assign t[158] = ~(t[239] | t[240]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[189] | t[190]);
  assign t[162] = ~(t[156] | t[191]);
  assign t[163] = ~(t[155] | t[192]);
  assign t[164] = ~(t[252]);
  assign t[165] = ~(t[242] | t[243]);
  assign t[166] = ~(t[253]);
  assign t[167] = ~(t[254]);
  assign t[168] = ~(t[193] | t[194]);
  assign t[169] = ~(t[195] | t[196]);
  assign t[16] = ~(t[213] & t[214]);
  assign t[170] = ~(t[50] | t[197]);
  assign t[171] = ~(x[4] | t[214]);
  assign t[172] = ~(t[216]);
  assign t[173] = x[4] & t[214];
  assign t[174] = ~(x[4] | t[198]);
  assign t[175] = ~(t[214] | t[216]);
  assign t[176] = ~(t[127] | t[199]);
  assign t[177] = ~(t[214] | t[172]);
  assign t[178] = t[82] & t[213];
  assign t[179] = ~(t[200] & t[201]);
  assign t[17] = ~(t[215] & t[216]);
  assign t[180] = t[213] ? t[202] : t[181];
  assign t[181] = ~(t[174] & t[172]);
  assign t[182] = t[213] ? t[128] : t[129];
  assign t[183] = ~(t[203] & t[204]);
  assign t[184] = t[213] ? t[181] : t[131];
  assign t[185] = ~(t[205] & t[88]);
  assign t[186] = ~(t[51] | t[197]);
  assign t[187] = t[213] ? t[207] : t[206];
  assign t[188] = t[213] ? t[128] : t[206];
  assign t[189] = ~(t[255]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[250] | t[251]);
  assign t[191] = ~(t[82] | t[208]);
  assign t[192] = ~(t[170] & t[88]);
  assign t[193] = ~(t[256]);
  assign t[194] = ~(t[253] | t[254]);
  assign t[195] = ~(t[162] & t[209]);
  assign t[196] = ~(t[183] & t[88]);
  assign t[197] = ~(t[82] | t[210]);
  assign t[198] = ~(t[214]);
  assign t[199] = t[213] ? t[206] : t[128];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[127] | t[213]);
  assign t[201] = ~(t[130] & t[202]);
  assign t[202] = ~(x[4] & t[177]);
  assign t[203] = t[216] & t[200];
  assign t[204] = t[171] | t[173];
  assign t[205] = ~(t[142]);
  assign t[206] = ~(t[173] & t[172]);
  assign t[207] = ~(t[171] & t[216]);
  assign t[208] = t[213] ? t[181] : t[202];
  assign t[209] = ~(t[127] & t[211]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = t[213] ? t[206] : t[207];
  assign t[211] = ~(t[131] & t[130]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = (t[301]);
  assign t[257] = t[302] ^ x[2];
  assign t[258] = t[303] ^ x[10];
  assign t[259] = t[304] ^ x[13];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[16];
  assign t[261] = t[306] ^ x[19];
  assign t[262] = t[307] ^ x[22];
  assign t[263] = t[308] ^ x[25];
  assign t[264] = t[309] ^ x[28];
  assign t[265] = t[310] ^ x[31];
  assign t[266] = t[311] ^ x[34];
  assign t[267] = t[312] ^ x[39];
  assign t[268] = t[313] ^ x[42];
  assign t[269] = t[314] ^ x[45];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[48];
  assign t[271] = t[316] ^ x[51];
  assign t[272] = t[317] ^ x[56];
  assign t[273] = t[318] ^ x[59];
  assign t[274] = t[319] ^ x[62];
  assign t[275] = t[320] ^ x[65];
  assign t[276] = t[321] ^ x[68];
  assign t[277] = t[322] ^ x[71];
  assign t[278] = t[323] ^ x[74];
  assign t[279] = t[324] ^ x[79];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[82];
  assign t[281] = t[326] ^ x[87];
  assign t[282] = t[327] ^ x[90];
  assign t[283] = t[328] ^ x[93];
  assign t[284] = t[329] ^ x[96];
  assign t[285] = t[330] ^ x[99];
  assign t[286] = t[331] ^ x[102];
  assign t[287] = t[332] ^ x[107];
  assign t[288] = t[333] ^ x[110];
  assign t[289] = t[334] ^ x[113];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[118];
  assign t[291] = t[336] ^ x[121];
  assign t[292] = t[337] ^ x[124];
  assign t[293] = t[338] ^ x[127];
  assign t[294] = t[339] ^ x[130];
  assign t[295] = t[340] ^ x[133];
  assign t[296] = t[341] ^ x[136];
  assign t[297] = t[342] ^ x[139];
  assign t[298] = t[343] ^ x[142];
  assign t[299] = t[344] ^ x[145];
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[148];
  assign t[301] = t[346] ^ x[151];
  assign t[302] = (t[347] & ~t[348]);
  assign t[303] = (t[349] & ~t[350]);
  assign t[304] = (t[351] & ~t[352]);
  assign t[305] = (t[353] & ~t[354]);
  assign t[306] = (t[355] & ~t[356]);
  assign t[307] = (t[357] & ~t[358]);
  assign t[308] = (t[359] & ~t[360]);
  assign t[309] = (t[361] & ~t[362]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[363] & ~t[364]);
  assign t[311] = (t[365] & ~t[366]);
  assign t[312] = (t[367] & ~t[368]);
  assign t[313] = (t[369] & ~t[370]);
  assign t[314] = (t[371] & ~t[372]);
  assign t[315] = (t[373] & ~t[374]);
  assign t[316] = (t[375] & ~t[376]);
  assign t[317] = (t[377] & ~t[378]);
  assign t[318] = (t[379] & ~t[380]);
  assign t[319] = (t[381] & ~t[382]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[383] & ~t[384]);
  assign t[321] = (t[385] & ~t[386]);
  assign t[322] = (t[387] & ~t[388]);
  assign t[323] = (t[389] & ~t[390]);
  assign t[324] = (t[391] & ~t[392]);
  assign t[325] = (t[393] & ~t[394]);
  assign t[326] = (t[395] & ~t[396]);
  assign t[327] = (t[397] & ~t[398]);
  assign t[328] = (t[399] & ~t[400]);
  assign t[329] = (t[401] & ~t[402]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[403] & ~t[404]);
  assign t[331] = (t[405] & ~t[406]);
  assign t[332] = (t[407] & ~t[408]);
  assign t[333] = (t[409] & ~t[410]);
  assign t[334] = (t[411] & ~t[412]);
  assign t[335] = (t[413] & ~t[414]);
  assign t[336] = (t[415] & ~t[416]);
  assign t[337] = (t[417] & ~t[418]);
  assign t[338] = (t[419] & ~t[420]);
  assign t[339] = (t[421] & ~t[422]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (t[423] & ~t[424]);
  assign t[341] = (t[425] & ~t[426]);
  assign t[342] = (t[427] & ~t[428]);
  assign t[343] = (t[429] & ~t[430]);
  assign t[344] = (t[431] & ~t[432]);
  assign t[345] = (t[433] & ~t[434]);
  assign t[346] = (t[435] & ~t[436]);
  assign t[347] = t[437] ^ x[2];
  assign t[348] = t[438] ^ x[1];
  assign t[349] = t[439] ^ x[10];
  assign t[34] = ~(t[217] | t[56]);
  assign t[350] = t[440] ^ x[9];
  assign t[351] = t[441] ^ x[13];
  assign t[352] = t[442] ^ x[12];
  assign t[353] = t[443] ^ x[16];
  assign t[354] = t[444] ^ x[15];
  assign t[355] = t[445] ^ x[19];
  assign t[356] = t[446] ^ x[18];
  assign t[357] = t[447] ^ x[22];
  assign t[358] = t[448] ^ x[21];
  assign t[359] = t[449] ^ x[25];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[24];
  assign t[361] = t[451] ^ x[28];
  assign t[362] = t[452] ^ x[27];
  assign t[363] = t[453] ^ x[31];
  assign t[364] = t[454] ^ x[30];
  assign t[365] = t[455] ^ x[34];
  assign t[366] = t[456] ^ x[33];
  assign t[367] = t[457] ^ x[39];
  assign t[368] = t[458] ^ x[38];
  assign t[369] = t[459] ^ x[42];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[41];
  assign t[371] = t[461] ^ x[45];
  assign t[372] = t[462] ^ x[44];
  assign t[373] = t[463] ^ x[48];
  assign t[374] = t[464] ^ x[47];
  assign t[375] = t[465] ^ x[51];
  assign t[376] = t[466] ^ x[50];
  assign t[377] = t[467] ^ x[56];
  assign t[378] = t[468] ^ x[55];
  assign t[379] = t[469] ^ x[59];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[58];
  assign t[381] = t[471] ^ x[62];
  assign t[382] = t[472] ^ x[61];
  assign t[383] = t[473] ^ x[65];
  assign t[384] = t[474] ^ x[64];
  assign t[385] = t[475] ^ x[68];
  assign t[386] = t[476] ^ x[67];
  assign t[387] = t[477] ^ x[71];
  assign t[388] = t[478] ^ x[70];
  assign t[389] = t[479] ^ x[74];
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[390] = t[480] ^ x[73];
  assign t[391] = t[481] ^ x[79];
  assign t[392] = t[482] ^ x[78];
  assign t[393] = t[483] ^ x[82];
  assign t[394] = t[484] ^ x[81];
  assign t[395] = t[485] ^ x[87];
  assign t[396] = t[486] ^ x[86];
  assign t[397] = t[487] ^ x[90];
  assign t[398] = t[488] ^ x[89];
  assign t[399] = t[489] ^ x[93];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[92];
  assign t[401] = t[491] ^ x[96];
  assign t[402] = t[492] ^ x[95];
  assign t[403] = t[493] ^ x[99];
  assign t[404] = t[494] ^ x[98];
  assign t[405] = t[495] ^ x[102];
  assign t[406] = t[496] ^ x[101];
  assign t[407] = t[497] ^ x[107];
  assign t[408] = t[498] ^ x[106];
  assign t[409] = t[499] ^ x[110];
  assign t[40] = ~(t[39] ^ t[66]);
  assign t[410] = t[500] ^ x[109];
  assign t[411] = t[501] ^ x[113];
  assign t[412] = t[502] ^ x[112];
  assign t[413] = t[503] ^ x[118];
  assign t[414] = t[504] ^ x[117];
  assign t[415] = t[505] ^ x[121];
  assign t[416] = t[506] ^ x[120];
  assign t[417] = t[507] ^ x[124];
  assign t[418] = t[508] ^ x[123];
  assign t[419] = t[509] ^ x[127];
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = t[510] ^ x[126];
  assign t[421] = t[511] ^ x[130];
  assign t[422] = t[512] ^ x[129];
  assign t[423] = t[513] ^ x[133];
  assign t[424] = t[514] ^ x[132];
  assign t[425] = t[515] ^ x[136];
  assign t[426] = t[516] ^ x[135];
  assign t[427] = t[517] ^ x[139];
  assign t[428] = t[518] ^ x[138];
  assign t[429] = t[519] ^ x[142];
  assign t[42] = ~(t[218] | t[69]);
  assign t[430] = t[520] ^ x[141];
  assign t[431] = t[521] ^ x[145];
  assign t[432] = t[522] ^ x[144];
  assign t[433] = t[523] ^ x[148];
  assign t[434] = t[524] ^ x[147];
  assign t[435] = t[525] ^ x[151];
  assign t[436] = t[526] ^ x[150];
  assign t[437] = (x[0]);
  assign t[438] = (x[0]);
  assign t[439] = (x[8]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[8]);
  assign t[441] = (x[11]);
  assign t[442] = (x[11]);
  assign t[443] = (x[14]);
  assign t[444] = (x[14]);
  assign t[445] = (x[17]);
  assign t[446] = (x[17]);
  assign t[447] = (x[20]);
  assign t[448] = (x[20]);
  assign t[449] = (x[23]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[23]);
  assign t[451] = (x[26]);
  assign t[452] = (x[26]);
  assign t[453] = (x[29]);
  assign t[454] = (x[29]);
  assign t[455] = (x[32]);
  assign t[456] = (x[32]);
  assign t[457] = (x[37]);
  assign t[458] = (x[37]);
  assign t[459] = (x[40]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[40]);
  assign t[461] = (x[43]);
  assign t[462] = (x[43]);
  assign t[463] = (x[46]);
  assign t[464] = (x[46]);
  assign t[465] = (x[49]);
  assign t[466] = (x[49]);
  assign t[467] = (x[54]);
  assign t[468] = (x[54]);
  assign t[469] = (x[57]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[470] = (x[57]);
  assign t[471] = (x[60]);
  assign t[472] = (x[60]);
  assign t[473] = (x[63]);
  assign t[474] = (x[63]);
  assign t[475] = (x[66]);
  assign t[476] = (x[66]);
  assign t[477] = (x[69]);
  assign t[478] = (x[69]);
  assign t[479] = (x[72]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = (x[72]);
  assign t[481] = (x[77]);
  assign t[482] = (x[77]);
  assign t[483] = (x[80]);
  assign t[484] = (x[80]);
  assign t[485] = (x[85]);
  assign t[486] = (x[85]);
  assign t[487] = (x[88]);
  assign t[488] = (x[88]);
  assign t[489] = (x[91]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = (x[91]);
  assign t[491] = (x[94]);
  assign t[492] = (x[94]);
  assign t[493] = (x[97]);
  assign t[494] = (x[97]);
  assign t[495] = (x[100]);
  assign t[496] = (x[100]);
  assign t[497] = (x[105]);
  assign t[498] = (x[105]);
  assign t[499] = (x[108]);
  assign t[49] = ~(t[215]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[108]);
  assign t[501] = (x[111]);
  assign t[502] = (x[111]);
  assign t[503] = (x[116]);
  assign t[504] = (x[116]);
  assign t[505] = (x[119]);
  assign t[506] = (x[119]);
  assign t[507] = (x[122]);
  assign t[508] = (x[122]);
  assign t[509] = (x[125]);
  assign t[50] = ~(t[82] | t[83]);
  assign t[510] = (x[125]);
  assign t[511] = (x[128]);
  assign t[512] = (x[128]);
  assign t[513] = (x[131]);
  assign t[514] = (x[131]);
  assign t[515] = (x[134]);
  assign t[516] = (x[134]);
  assign t[517] = (x[137]);
  assign t[518] = (x[137]);
  assign t[519] = (x[140]);
  assign t[51] = ~(t[82] | t[84]);
  assign t[520] = (x[140]);
  assign t[521] = (x[143]);
  assign t[522] = (x[143]);
  assign t[523] = (x[146]);
  assign t[524] = (x[146]);
  assign t[525] = (x[149]);
  assign t[526] = (x[149]);
  assign t[52] = t[85] | t[86];
  assign t[53] = ~(t[87] & t[88]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[220]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[221] | t[93]);
  assign t[59] = t[215] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[222] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[223] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[224]);
  assign t[68] = ~(t[225]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[226] | t[110]);
  assign t[72] = t[30] ? x[53] : x[52];
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[227] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[228] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] | t[124]);
  assign t[81] = ~(t[125] ^ t[126]);
  assign t[82] = ~(t[127]);
  assign t[83] = t[213] ? t[129] : t[128];
  assign t[84] = t[213] ? t[131] : t[130];
  assign t[85] = ~(t[132] & t[133]);
  assign t[86] = ~(t[82] | t[134]);
  assign t[87] = ~(t[135] | t[136]);
  assign t[88] = t[127] | t[137];
  assign t[89] = ~(t[229]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[219] | t[220]);
  assign t[91] = ~(t[230]);
  assign t[92] = ~(t[231]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[140] | t[141]);
  assign t[95] = ~(t[142] | t[143]);
  assign t[96] = ~(t[232]);
  assign t[97] = ~(t[233]);
  assign t[98] = ~(t[144] | t[145]);
  assign t[99] = t[146] ? x[76] : x[75];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [151:0] x;
 output y;

 wire [526:0] t;
  assign t[0] = t[1] ? t[2] : t[212];
  assign t[100] = ~(t[147] & t[148]);
  assign t[101] = ~(t[234]);
  assign t[102] = ~(t[235]);
  assign t[103] = ~(t[149] | t[150]);
  assign t[104] = t[215] ? x[84] : x[83];
  assign t[105] = t[151] | t[152];
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[224] | t[225]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[153] | t[154]);
  assign t[111] = ~(t[140] | t[155]);
  assign t[112] = ~(t[156] | t[85]);
  assign t[113] = ~(t[239]);
  assign t[114] = ~(t[240]);
  assign t[115] = ~(t[157] | t[158]);
  assign t[116] = ~(t[159] | t[160]);
  assign t[117] = ~(t[241] | t[161]);
  assign t[118] = t[30] ? x[104] : x[103];
  assign t[119] = ~(t[162] & t[163]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[243]);
  assign t[122] = ~(t[164] | t[165]);
  assign t[123] = ~(t[166] | t[167]);
  assign t[124] = ~(t[244] | t[168]);
  assign t[125] = t[30] ? x[115] : x[114];
  assign t[126] = ~(t[169] & t[170]);
  assign t[127] = ~(t[215]);
  assign t[128] = ~(t[171] & t[172]);
  assign t[129] = ~(t[173] & t[216]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[216] & t[174]);
  assign t[131] = ~(x[4] & t[175]);
  assign t[132] = ~(t[176] | t[142]);
  assign t[133] = ~(t[177] & t[178]);
  assign t[134] = t[213] ? t[130] : t[131];
  assign t[135] = ~(t[179]);
  assign t[136] = ~(t[82] | t[180]);
  assign t[137] = t[213] ? t[131] : t[181];
  assign t[138] = ~(t[245]);
  assign t[139] = ~(t[230] | t[231]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[82] | t[182]);
  assign t[141] = ~(t[31] & t[183]);
  assign t[142] = ~(t[127] | t[184]);
  assign t[143] = t[155] | t[135];
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[232] | t[233]);
  assign t[146] = ~(t[49]);
  assign t[147] = ~(t[151] | t[185]);
  assign t[148] = ~(t[140]);
  assign t[149] = ~(t[247]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[234] | t[235]);
  assign t[151] = ~(t[179] & t[133]);
  assign t[152] = ~(t[111] & t[186]);
  assign t[153] = ~(t[248]);
  assign t[154] = ~(t[237] | t[238]);
  assign t[155] = ~(t[82] | t[187]);
  assign t[156] = ~(t[127] | t[188]);
  assign t[157] = ~(t[249]);
  assign t[158] = ~(t[239] | t[240]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[189] | t[190]);
  assign t[162] = ~(t[156] | t[191]);
  assign t[163] = ~(t[155] | t[192]);
  assign t[164] = ~(t[252]);
  assign t[165] = ~(t[242] | t[243]);
  assign t[166] = ~(t[253]);
  assign t[167] = ~(t[254]);
  assign t[168] = ~(t[193] | t[194]);
  assign t[169] = ~(t[195] | t[196]);
  assign t[16] = ~(t[213] & t[214]);
  assign t[170] = ~(t[50] | t[197]);
  assign t[171] = ~(x[4] | t[214]);
  assign t[172] = ~(t[216]);
  assign t[173] = x[4] & t[214];
  assign t[174] = ~(x[4] | t[198]);
  assign t[175] = ~(t[214] | t[216]);
  assign t[176] = ~(t[127] | t[199]);
  assign t[177] = ~(t[214] | t[172]);
  assign t[178] = t[82] & t[213];
  assign t[179] = ~(t[200] & t[201]);
  assign t[17] = ~(t[215] & t[216]);
  assign t[180] = t[213] ? t[202] : t[181];
  assign t[181] = ~(t[174] & t[172]);
  assign t[182] = t[213] ? t[128] : t[129];
  assign t[183] = ~(t[203] & t[204]);
  assign t[184] = t[213] ? t[181] : t[131];
  assign t[185] = ~(t[205] & t[88]);
  assign t[186] = ~(t[51] | t[197]);
  assign t[187] = t[213] ? t[207] : t[206];
  assign t[188] = t[213] ? t[128] : t[206];
  assign t[189] = ~(t[255]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[250] | t[251]);
  assign t[191] = ~(t[82] | t[208]);
  assign t[192] = ~(t[170] & t[88]);
  assign t[193] = ~(t[256]);
  assign t[194] = ~(t[253] | t[254]);
  assign t[195] = ~(t[162] & t[209]);
  assign t[196] = ~(t[183] & t[88]);
  assign t[197] = ~(t[82] | t[210]);
  assign t[198] = ~(t[214]);
  assign t[199] = t[213] ? t[206] : t[128];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[127] | t[213]);
  assign t[201] = ~(t[130] & t[202]);
  assign t[202] = ~(x[4] & t[177]);
  assign t[203] = t[216] & t[200];
  assign t[204] = t[171] | t[173];
  assign t[205] = ~(t[142]);
  assign t[206] = ~(t[173] & t[172]);
  assign t[207] = ~(t[171] & t[216]);
  assign t[208] = t[213] ? t[181] : t[202];
  assign t[209] = ~(t[127] & t[211]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = t[213] ? t[206] : t[207];
  assign t[211] = ~(t[131] & t[130]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = (t[301]);
  assign t[257] = t[302] ^ x[2];
  assign t[258] = t[303] ^ x[10];
  assign t[259] = t[304] ^ x[13];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[16];
  assign t[261] = t[306] ^ x[19];
  assign t[262] = t[307] ^ x[22];
  assign t[263] = t[308] ^ x[25];
  assign t[264] = t[309] ^ x[28];
  assign t[265] = t[310] ^ x[31];
  assign t[266] = t[311] ^ x[34];
  assign t[267] = t[312] ^ x[39];
  assign t[268] = t[313] ^ x[42];
  assign t[269] = t[314] ^ x[45];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[48];
  assign t[271] = t[316] ^ x[51];
  assign t[272] = t[317] ^ x[56];
  assign t[273] = t[318] ^ x[59];
  assign t[274] = t[319] ^ x[62];
  assign t[275] = t[320] ^ x[65];
  assign t[276] = t[321] ^ x[68];
  assign t[277] = t[322] ^ x[71];
  assign t[278] = t[323] ^ x[74];
  assign t[279] = t[324] ^ x[79];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[82];
  assign t[281] = t[326] ^ x[87];
  assign t[282] = t[327] ^ x[90];
  assign t[283] = t[328] ^ x[93];
  assign t[284] = t[329] ^ x[96];
  assign t[285] = t[330] ^ x[99];
  assign t[286] = t[331] ^ x[102];
  assign t[287] = t[332] ^ x[107];
  assign t[288] = t[333] ^ x[110];
  assign t[289] = t[334] ^ x[113];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[118];
  assign t[291] = t[336] ^ x[121];
  assign t[292] = t[337] ^ x[124];
  assign t[293] = t[338] ^ x[127];
  assign t[294] = t[339] ^ x[130];
  assign t[295] = t[340] ^ x[133];
  assign t[296] = t[341] ^ x[136];
  assign t[297] = t[342] ^ x[139];
  assign t[298] = t[343] ^ x[142];
  assign t[299] = t[344] ^ x[145];
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[148];
  assign t[301] = t[346] ^ x[151];
  assign t[302] = (t[347] & ~t[348]);
  assign t[303] = (t[349] & ~t[350]);
  assign t[304] = (t[351] & ~t[352]);
  assign t[305] = (t[353] & ~t[354]);
  assign t[306] = (t[355] & ~t[356]);
  assign t[307] = (t[357] & ~t[358]);
  assign t[308] = (t[359] & ~t[360]);
  assign t[309] = (t[361] & ~t[362]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[363] & ~t[364]);
  assign t[311] = (t[365] & ~t[366]);
  assign t[312] = (t[367] & ~t[368]);
  assign t[313] = (t[369] & ~t[370]);
  assign t[314] = (t[371] & ~t[372]);
  assign t[315] = (t[373] & ~t[374]);
  assign t[316] = (t[375] & ~t[376]);
  assign t[317] = (t[377] & ~t[378]);
  assign t[318] = (t[379] & ~t[380]);
  assign t[319] = (t[381] & ~t[382]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[383] & ~t[384]);
  assign t[321] = (t[385] & ~t[386]);
  assign t[322] = (t[387] & ~t[388]);
  assign t[323] = (t[389] & ~t[390]);
  assign t[324] = (t[391] & ~t[392]);
  assign t[325] = (t[393] & ~t[394]);
  assign t[326] = (t[395] & ~t[396]);
  assign t[327] = (t[397] & ~t[398]);
  assign t[328] = (t[399] & ~t[400]);
  assign t[329] = (t[401] & ~t[402]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (t[403] & ~t[404]);
  assign t[331] = (t[405] & ~t[406]);
  assign t[332] = (t[407] & ~t[408]);
  assign t[333] = (t[409] & ~t[410]);
  assign t[334] = (t[411] & ~t[412]);
  assign t[335] = (t[413] & ~t[414]);
  assign t[336] = (t[415] & ~t[416]);
  assign t[337] = (t[417] & ~t[418]);
  assign t[338] = (t[419] & ~t[420]);
  assign t[339] = (t[421] & ~t[422]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (t[423] & ~t[424]);
  assign t[341] = (t[425] & ~t[426]);
  assign t[342] = (t[427] & ~t[428]);
  assign t[343] = (t[429] & ~t[430]);
  assign t[344] = (t[431] & ~t[432]);
  assign t[345] = (t[433] & ~t[434]);
  assign t[346] = (t[435] & ~t[436]);
  assign t[347] = t[437] ^ x[2];
  assign t[348] = t[438] ^ x[1];
  assign t[349] = t[439] ^ x[10];
  assign t[34] = ~(t[217] | t[56]);
  assign t[350] = t[440] ^ x[9];
  assign t[351] = t[441] ^ x[13];
  assign t[352] = t[442] ^ x[12];
  assign t[353] = t[443] ^ x[16];
  assign t[354] = t[444] ^ x[15];
  assign t[355] = t[445] ^ x[19];
  assign t[356] = t[446] ^ x[18];
  assign t[357] = t[447] ^ x[22];
  assign t[358] = t[448] ^ x[21];
  assign t[359] = t[449] ^ x[25];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[24];
  assign t[361] = t[451] ^ x[28];
  assign t[362] = t[452] ^ x[27];
  assign t[363] = t[453] ^ x[31];
  assign t[364] = t[454] ^ x[30];
  assign t[365] = t[455] ^ x[34];
  assign t[366] = t[456] ^ x[33];
  assign t[367] = t[457] ^ x[39];
  assign t[368] = t[458] ^ x[38];
  assign t[369] = t[459] ^ x[42];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[41];
  assign t[371] = t[461] ^ x[45];
  assign t[372] = t[462] ^ x[44];
  assign t[373] = t[463] ^ x[48];
  assign t[374] = t[464] ^ x[47];
  assign t[375] = t[465] ^ x[51];
  assign t[376] = t[466] ^ x[50];
  assign t[377] = t[467] ^ x[56];
  assign t[378] = t[468] ^ x[55];
  assign t[379] = t[469] ^ x[59];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[58];
  assign t[381] = t[471] ^ x[62];
  assign t[382] = t[472] ^ x[61];
  assign t[383] = t[473] ^ x[65];
  assign t[384] = t[474] ^ x[64];
  assign t[385] = t[475] ^ x[68];
  assign t[386] = t[476] ^ x[67];
  assign t[387] = t[477] ^ x[71];
  assign t[388] = t[478] ^ x[70];
  assign t[389] = t[479] ^ x[74];
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[390] = t[480] ^ x[73];
  assign t[391] = t[481] ^ x[79];
  assign t[392] = t[482] ^ x[78];
  assign t[393] = t[483] ^ x[82];
  assign t[394] = t[484] ^ x[81];
  assign t[395] = t[485] ^ x[87];
  assign t[396] = t[486] ^ x[86];
  assign t[397] = t[487] ^ x[90];
  assign t[398] = t[488] ^ x[89];
  assign t[399] = t[489] ^ x[93];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[92];
  assign t[401] = t[491] ^ x[96];
  assign t[402] = t[492] ^ x[95];
  assign t[403] = t[493] ^ x[99];
  assign t[404] = t[494] ^ x[98];
  assign t[405] = t[495] ^ x[102];
  assign t[406] = t[496] ^ x[101];
  assign t[407] = t[497] ^ x[107];
  assign t[408] = t[498] ^ x[106];
  assign t[409] = t[499] ^ x[110];
  assign t[40] = ~(t[39] ^ t[66]);
  assign t[410] = t[500] ^ x[109];
  assign t[411] = t[501] ^ x[113];
  assign t[412] = t[502] ^ x[112];
  assign t[413] = t[503] ^ x[118];
  assign t[414] = t[504] ^ x[117];
  assign t[415] = t[505] ^ x[121];
  assign t[416] = t[506] ^ x[120];
  assign t[417] = t[507] ^ x[124];
  assign t[418] = t[508] ^ x[123];
  assign t[419] = t[509] ^ x[127];
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = t[510] ^ x[126];
  assign t[421] = t[511] ^ x[130];
  assign t[422] = t[512] ^ x[129];
  assign t[423] = t[513] ^ x[133];
  assign t[424] = t[514] ^ x[132];
  assign t[425] = t[515] ^ x[136];
  assign t[426] = t[516] ^ x[135];
  assign t[427] = t[517] ^ x[139];
  assign t[428] = t[518] ^ x[138];
  assign t[429] = t[519] ^ x[142];
  assign t[42] = ~(t[218] | t[69]);
  assign t[430] = t[520] ^ x[141];
  assign t[431] = t[521] ^ x[145];
  assign t[432] = t[522] ^ x[144];
  assign t[433] = t[523] ^ x[148];
  assign t[434] = t[524] ^ x[147];
  assign t[435] = t[525] ^ x[151];
  assign t[436] = t[526] ^ x[150];
  assign t[437] = (x[0]);
  assign t[438] = (x[0]);
  assign t[439] = (x[8]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[8]);
  assign t[441] = (x[11]);
  assign t[442] = (x[11]);
  assign t[443] = (x[14]);
  assign t[444] = (x[14]);
  assign t[445] = (x[17]);
  assign t[446] = (x[17]);
  assign t[447] = (x[20]);
  assign t[448] = (x[20]);
  assign t[449] = (x[23]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[23]);
  assign t[451] = (x[26]);
  assign t[452] = (x[26]);
  assign t[453] = (x[29]);
  assign t[454] = (x[29]);
  assign t[455] = (x[32]);
  assign t[456] = (x[32]);
  assign t[457] = (x[37]);
  assign t[458] = (x[37]);
  assign t[459] = (x[40]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[40]);
  assign t[461] = (x[43]);
  assign t[462] = (x[43]);
  assign t[463] = (x[46]);
  assign t[464] = (x[46]);
  assign t[465] = (x[49]);
  assign t[466] = (x[49]);
  assign t[467] = (x[54]);
  assign t[468] = (x[54]);
  assign t[469] = (x[57]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[470] = (x[57]);
  assign t[471] = (x[60]);
  assign t[472] = (x[60]);
  assign t[473] = (x[63]);
  assign t[474] = (x[63]);
  assign t[475] = (x[66]);
  assign t[476] = (x[66]);
  assign t[477] = (x[69]);
  assign t[478] = (x[69]);
  assign t[479] = (x[72]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = (x[72]);
  assign t[481] = (x[77]);
  assign t[482] = (x[77]);
  assign t[483] = (x[80]);
  assign t[484] = (x[80]);
  assign t[485] = (x[85]);
  assign t[486] = (x[85]);
  assign t[487] = (x[88]);
  assign t[488] = (x[88]);
  assign t[489] = (x[91]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = (x[91]);
  assign t[491] = (x[94]);
  assign t[492] = (x[94]);
  assign t[493] = (x[97]);
  assign t[494] = (x[97]);
  assign t[495] = (x[100]);
  assign t[496] = (x[100]);
  assign t[497] = (x[105]);
  assign t[498] = (x[105]);
  assign t[499] = (x[108]);
  assign t[49] = ~(t[215]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[108]);
  assign t[501] = (x[111]);
  assign t[502] = (x[111]);
  assign t[503] = (x[116]);
  assign t[504] = (x[116]);
  assign t[505] = (x[119]);
  assign t[506] = (x[119]);
  assign t[507] = (x[122]);
  assign t[508] = (x[122]);
  assign t[509] = (x[125]);
  assign t[50] = ~(t[82] | t[83]);
  assign t[510] = (x[125]);
  assign t[511] = (x[128]);
  assign t[512] = (x[128]);
  assign t[513] = (x[131]);
  assign t[514] = (x[131]);
  assign t[515] = (x[134]);
  assign t[516] = (x[134]);
  assign t[517] = (x[137]);
  assign t[518] = (x[137]);
  assign t[519] = (x[140]);
  assign t[51] = ~(t[82] | t[84]);
  assign t[520] = (x[140]);
  assign t[521] = (x[143]);
  assign t[522] = (x[143]);
  assign t[523] = (x[146]);
  assign t[524] = (x[146]);
  assign t[525] = (x[149]);
  assign t[526] = (x[149]);
  assign t[52] = t[85] | t[86];
  assign t[53] = ~(t[87] & t[88]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[220]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[221] | t[93]);
  assign t[59] = t[215] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[222] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[223] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[224]);
  assign t[68] = ~(t[225]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[226] | t[110]);
  assign t[72] = t[30] ? x[53] : x[52];
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[227] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[228] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] | t[124]);
  assign t[81] = ~(t[125] ^ t[126]);
  assign t[82] = ~(t[127]);
  assign t[83] = t[213] ? t[129] : t[128];
  assign t[84] = t[213] ? t[131] : t[130];
  assign t[85] = ~(t[132] & t[133]);
  assign t[86] = ~(t[82] | t[134]);
  assign t[87] = ~(t[135] | t[136]);
  assign t[88] = t[127] | t[137];
  assign t[89] = ~(t[229]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[219] | t[220]);
  assign t[91] = ~(t[230]);
  assign t[92] = ~(t[231]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[140] | t[141]);
  assign t[95] = ~(t[142] | t[143]);
  assign t[96] = ~(t[232]);
  assign t[97] = ~(t[233]);
  assign t[98] = ~(t[144] | t[145]);
  assign t[99] = t[146] ? x[76] : x[75];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[44];
  assign t[38] = ~(t[107] & t[57]);
  assign t[39] = ~(t[108] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[59] ? x[35] : x[34];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[103] ? x[52] : x[51];
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = ~(t[115] & t[76]);
  assign t[56] = t[103] ? x[60] : x[59];
  assign t[57] = ~(t[116]);
  assign t[58] = ~(t[116] & t[77]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[78]);
  assign t[61] = ~(t[118] & t[79]);
  assign t[62] = ~(t[119] & t[80]);
  assign t[63] = ~(t[120] & t[81]);
  assign t[64] = t[48] ? x[77] : x[76];
  assign t[65] = ~(t[82] & t[83]);
  assign t[66] = ~(t[121] & t[84]);
  assign t[67] = ~(t[122] & t[85]);
  assign t[68] = t[18] ? x[85] : x[84];
  assign t[69] = ~(t[86] & t[87]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[107]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[114]);
  assign t[91] = ~(t[117]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[133]);
  assign t[94] = ~(t[133] & t[98]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[128]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[44];
  assign t[38] = ~(t[107] & t[57]);
  assign t[39] = ~(t[108] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[59] ? x[35] : x[34];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[103] ? x[52] : x[51];
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = ~(t[115] & t[76]);
  assign t[56] = t[103] ? x[60] : x[59];
  assign t[57] = ~(t[116]);
  assign t[58] = ~(t[116] & t[77]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[78]);
  assign t[61] = ~(t[118] & t[79]);
  assign t[62] = ~(t[119] & t[80]);
  assign t[63] = ~(t[120] & t[81]);
  assign t[64] = t[48] ? x[77] : x[76];
  assign t[65] = ~(t[82] & t[83]);
  assign t[66] = ~(t[121] & t[84]);
  assign t[67] = ~(t[122] & t[85]);
  assign t[68] = t[18] ? x[85] : x[84];
  assign t[69] = ~(t[86] & t[87]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[107]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[114]);
  assign t[91] = ~(t[117]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[133]);
  assign t[94] = ~(t[133] & t[98]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[128]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[145] & t[144]);
  assign t[104] = ~(t[155]);
  assign t[105] = ~(t[147] & t[146]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[115] & t[116]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[53] ^ t[44];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[56] ^ t[36];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[59] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[122] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[128]);
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = ~(t[77] & t[129]);
  assign t[53] = t[122] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[130]);
  assign t[56] = t[122] ? x[48] : x[47];
  assign t[57] = ~(t[131]);
  assign t[58] = ~(t[132]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[133]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[134]);
  assign t[64] = t[18] ? x[62] : x[61];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[135]);
  assign t[68] = t[94] ? x[67] : x[66];
  assign t[69] = ~(t[95] & t[96]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127] & t[126]);
  assign t[71] = ~(t[136]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[97] & t[98]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[140]);
  assign t[77] = ~(t[99] & t[100]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[142]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[132] & t[131]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[145]);
  assign t[85] = ~(t[103] & t[104]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[147]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[109] & t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[150]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[25]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind201(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[145] & t[144]);
  assign t[104] = ~(t[155]);
  assign t[105] = ~(t[147] & t[146]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[115] & t[116]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[53] ^ t[44];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[56] ^ t[36];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[59] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[122] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[128]);
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = ~(t[77] & t[129]);
  assign t[53] = t[122] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[130]);
  assign t[56] = t[122] ? x[48] : x[47];
  assign t[57] = ~(t[131]);
  assign t[58] = ~(t[132]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[133]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[134]);
  assign t[64] = t[18] ? x[62] : x[61];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[135]);
  assign t[68] = t[94] ? x[67] : x[66];
  assign t[69] = ~(t[95] & t[96]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127] & t[126]);
  assign t[71] = ~(t[136]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[97] & t[98]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[140]);
  assign t[77] = ~(t[99] & t[100]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[142]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[132] & t[131]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[145]);
  assign t[85] = ~(t[103] & t[104]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[147]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[109] & t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[150]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[25]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[44];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[57] ^ t[36];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[113] ? x[43] : x[42];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = t[80] | t[121];
  assign t[57] = t[113] ? x[48] : x[47];
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] | t[58]);
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[124];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[125];
  assign t[65] = t[18] ? x[62] : x[61];
  assign t[66] = ~(t[88] & t[89]);
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = t[92] | t[126];
  assign t[69] = t[93] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[139];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[140]);
  assign t[91] = ~(t[141]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[25]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[44];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[57] ^ t[36];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[58] & t[59]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[113] ? x[43] : x[42];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = t[80] | t[121];
  assign t[57] = t[113] ? x[48] : x[47];
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] | t[58]);
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[124];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[125];
  assign t[65] = t[18] ? x[62] : x[61];
  assign t[66] = ~(t[88] & t[89]);
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = t[92] | t[126];
  assign t[69] = t[93] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[139];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[140]);
  assign t[91] = ~(t[141]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[25]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [139:0] x;
 output y;

 wire [481:0] t;
  assign t[0] = t[1] ? t[2] : t[195];
  assign t[100] = ~(t[217]);
  assign t[101] = ~(t[206] | t[207]);
  assign t[102] = ~(t[218]);
  assign t[103] = ~(t[219]);
  assign t[104] = ~(t[138] | t[139]);
  assign t[105] = ~(t[86] | t[140]);
  assign t[106] = ~(t[141] & t[142]);
  assign t[107] = ~(t[220]);
  assign t[108] = ~(t[221]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[145] ? x[95] : x[94];
  assign t[111] = t[146] | t[147];
  assign t[112] = ~(t[222]);
  assign t[113] = ~(t[223]);
  assign t[114] = ~(t[148] | t[149]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[224] | t[152]);
  assign t[117] = t[145] ? x[106] : x[105];
  assign t[118] = ~(t[153] & t[154]);
  assign t[119] = ~(t[198]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[155] & t[83]);
  assign t[121] = ~(t[156] & t[199]);
  assign t[122] = ~(t[119] | t[157]);
  assign t[123] = ~(t[79] | t[158]);
  assign t[124] = ~(t[159] & t[160]);
  assign t[125] = ~(t[161] & t[162]);
  assign t[126] = ~(t[163] | t[164]);
  assign t[127] = ~(t[165] | t[166]);
  assign t[128] = ~(t[225]);
  assign t[129] = ~(t[212] | t[213]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[163] | t[167]);
  assign t[131] = ~(t[168] | t[169]);
  assign t[132] = ~(t[226]);
  assign t[133] = ~(t[214] | t[215]);
  assign t[134] = ~(t[227]);
  assign t[135] = ~(t[228]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[166]);
  assign t[138] = ~(t[229]);
  assign t[139] = ~(t[218] | t[219]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[147] | t[164];
  assign t[141] = t[199] & t[161];
  assign t[142] = t[155] | t[156];
  assign t[143] = ~(t[230]);
  assign t[144] = ~(t[220] | t[221]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[173] & t[32]);
  assign t[147] = ~(t[79] | t[174]);
  assign t[148] = ~(t[231]);
  assign t[149] = ~(t[222] | t[223]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[232]);
  assign t[151] = ~(t[233]);
  assign t[152] = ~(t[175] | t[176]);
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[177] | t[147]);
  assign t[155] = ~(x[4] | t[197]);
  assign t[156] = x[4] & t[197];
  assign t[157] = t[196] ? t[120] : t[178];
  assign t[158] = t[196] ? t[180] : t[179];
  assign t[159] = ~(x[4] & t[181]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[199] & t[182]);
  assign t[161] = ~(t[119] | t[196]);
  assign t[162] = ~(t[160] & t[179]);
  assign t[163] = ~(t[79] | t[183]);
  assign t[164] = ~(t[79] | t[184]);
  assign t[165] = ~(t[79] | t[185]);
  assign t[166] = ~(t[79] | t[186]);
  assign t[167] = ~(t[187] & t[106]);
  assign t[168] = ~(t[119] | t[188]);
  assign t[169] = t[164] | t[189];
  assign t[16] = ~(t[196] & t[197]);
  assign t[170] = ~(t[234]);
  assign t[171] = ~(t[227] | t[228]);
  assign t[172] = ~(t[79] | t[190]);
  assign t[173] = ~(t[191] | t[168]);
  assign t[174] = t[196] ? t[160] : t[159];
  assign t[175] = ~(t[235]);
  assign t[176] = ~(t[232] | t[233]);
  assign t[177] = ~(t[137]);
  assign t[178] = ~(t[156] & t[83]);
  assign t[179] = ~(x[4] & t[51]);
  assign t[17] = ~(t[198] & t[199]);
  assign t[180] = ~(t[182] & t[83]);
  assign t[181] = ~(t[197] | t[199]);
  assign t[182] = ~(x[4] | t[192]);
  assign t[183] = t[196] ? t[120] : t[121];
  assign t[184] = t[196] ? t[193] : t[178];
  assign t[185] = t[196] ? t[159] : t[160];
  assign t[186] = t[196] ? t[178] : t[193];
  assign t[187] = ~(t[49] | t[165]);
  assign t[188] = t[196] ? t[180] : t[159];
  assign t[189] = ~(t[125]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[196] ? t[179] : t[180];
  assign t[191] = ~(t[119] | t[194]);
  assign t[192] = ~(t[197]);
  assign t[193] = ~(t[155] & t[199]);
  assign t[194] = t[196] ? t[178] : t[120];
  assign t[195] = (t[236]);
  assign t[196] = (t[237]);
  assign t[197] = (t[238]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = t[277] ^ x[2];
  assign t[237] = t[278] ^ x[10];
  assign t[238] = t[279] ^ x[13];
  assign t[239] = t[280] ^ x[16];
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = t[281] ^ x[19];
  assign t[241] = t[282] ^ x[22];
  assign t[242] = t[283] ^ x[25];
  assign t[243] = t[284] ^ x[28];
  assign t[244] = t[285] ^ x[31];
  assign t[245] = t[286] ^ x[36];
  assign t[246] = t[287] ^ x[39];
  assign t[247] = t[288] ^ x[42];
  assign t[248] = t[289] ^ x[45];
  assign t[249] = t[290] ^ x[48];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[53];
  assign t[251] = t[292] ^ x[56];
  assign t[252] = t[293] ^ x[59];
  assign t[253] = t[294] ^ x[62];
  assign t[254] = t[295] ^ x[65];
  assign t[255] = t[296] ^ x[70];
  assign t[256] = t[297] ^ x[73];
  assign t[257] = t[298] ^ x[76];
  assign t[258] = t[299] ^ x[81];
  assign t[259] = t[300] ^ x[84];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[87];
  assign t[261] = t[302] ^ x[90];
  assign t[262] = t[303] ^ x[93];
  assign t[263] = t[304] ^ x[98];
  assign t[264] = t[305] ^ x[101];
  assign t[265] = t[306] ^ x[104];
  assign t[266] = t[307] ^ x[109];
  assign t[267] = t[308] ^ x[112];
  assign t[268] = t[309] ^ x[115];
  assign t[269] = t[310] ^ x[118];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[121];
  assign t[271] = t[312] ^ x[124];
  assign t[272] = t[313] ^ x[127];
  assign t[273] = t[314] ^ x[130];
  assign t[274] = t[315] ^ x[133];
  assign t[275] = t[316] ^ x[136];
  assign t[276] = t[317] ^ x[139];
  assign t[277] = (t[318] & ~t[319]);
  assign t[278] = (t[320] & ~t[321]);
  assign t[279] = (t[322] & ~t[323]);
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = (t[324] & ~t[325]);
  assign t[281] = (t[326] & ~t[327]);
  assign t[282] = (t[328] & ~t[329]);
  assign t[283] = (t[330] & ~t[331]);
  assign t[284] = (t[332] & ~t[333]);
  assign t[285] = (t[334] & ~t[335]);
  assign t[286] = (t[336] & ~t[337]);
  assign t[287] = (t[338] & ~t[339]);
  assign t[288] = (t[340] & ~t[341]);
  assign t[289] = (t[342] & ~t[343]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[344] & ~t[345]);
  assign t[291] = (t[346] & ~t[347]);
  assign t[292] = (t[348] & ~t[349]);
  assign t[293] = (t[350] & ~t[351]);
  assign t[294] = (t[352] & ~t[353]);
  assign t[295] = (t[354] & ~t[355]);
  assign t[296] = (t[356] & ~t[357]);
  assign t[297] = (t[358] & ~t[359]);
  assign t[298] = (t[360] & ~t[361]);
  assign t[299] = (t[362] & ~t[363]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[364] & ~t[365]);
  assign t[301] = (t[366] & ~t[367]);
  assign t[302] = (t[368] & ~t[369]);
  assign t[303] = (t[370] & ~t[371]);
  assign t[304] = (t[372] & ~t[373]);
  assign t[305] = (t[374] & ~t[375]);
  assign t[306] = (t[376] & ~t[377]);
  assign t[307] = (t[378] & ~t[379]);
  assign t[308] = (t[380] & ~t[381]);
  assign t[309] = (t[382] & ~t[383]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[384] & ~t[385]);
  assign t[311] = (t[386] & ~t[387]);
  assign t[312] = (t[388] & ~t[389]);
  assign t[313] = (t[390] & ~t[391]);
  assign t[314] = (t[392] & ~t[393]);
  assign t[315] = (t[394] & ~t[395]);
  assign t[316] = (t[396] & ~t[397]);
  assign t[317] = (t[398] & ~t[399]);
  assign t[318] = t[400] ^ x[2];
  assign t[319] = t[401] ^ x[1];
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = t[402] ^ x[10];
  assign t[321] = t[403] ^ x[9];
  assign t[322] = t[404] ^ x[13];
  assign t[323] = t[405] ^ x[12];
  assign t[324] = t[406] ^ x[16];
  assign t[325] = t[407] ^ x[15];
  assign t[326] = t[408] ^ x[19];
  assign t[327] = t[409] ^ x[18];
  assign t[328] = t[410] ^ x[22];
  assign t[329] = t[411] ^ x[21];
  assign t[32] = ~(t[51] & t[52]);
  assign t[330] = t[412] ^ x[25];
  assign t[331] = t[413] ^ x[24];
  assign t[332] = t[414] ^ x[28];
  assign t[333] = t[415] ^ x[27];
  assign t[334] = t[416] ^ x[31];
  assign t[335] = t[417] ^ x[30];
  assign t[336] = t[418] ^ x[36];
  assign t[337] = t[419] ^ x[35];
  assign t[338] = t[420] ^ x[39];
  assign t[339] = t[421] ^ x[38];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[42];
  assign t[341] = t[423] ^ x[41];
  assign t[342] = t[424] ^ x[45];
  assign t[343] = t[425] ^ x[44];
  assign t[344] = t[426] ^ x[48];
  assign t[345] = t[427] ^ x[47];
  assign t[346] = t[428] ^ x[53];
  assign t[347] = t[429] ^ x[52];
  assign t[348] = t[430] ^ x[56];
  assign t[349] = t[431] ^ x[55];
  assign t[34] = ~(t[200] | t[55]);
  assign t[350] = t[432] ^ x[59];
  assign t[351] = t[433] ^ x[58];
  assign t[352] = t[434] ^ x[62];
  assign t[353] = t[435] ^ x[61];
  assign t[354] = t[436] ^ x[65];
  assign t[355] = t[437] ^ x[64];
  assign t[356] = t[438] ^ x[70];
  assign t[357] = t[439] ^ x[69];
  assign t[358] = t[440] ^ x[73];
  assign t[359] = t[441] ^ x[72];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[76];
  assign t[361] = t[443] ^ x[75];
  assign t[362] = t[444] ^ x[81];
  assign t[363] = t[445] ^ x[80];
  assign t[364] = t[446] ^ x[84];
  assign t[365] = t[447] ^ x[83];
  assign t[366] = t[448] ^ x[87];
  assign t[367] = t[449] ^ x[86];
  assign t[368] = t[450] ^ x[90];
  assign t[369] = t[451] ^ x[89];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[93];
  assign t[371] = t[453] ^ x[92];
  assign t[372] = t[454] ^ x[98];
  assign t[373] = t[455] ^ x[97];
  assign t[374] = t[456] ^ x[101];
  assign t[375] = t[457] ^ x[100];
  assign t[376] = t[458] ^ x[104];
  assign t[377] = t[459] ^ x[103];
  assign t[378] = t[460] ^ x[109];
  assign t[379] = t[461] ^ x[108];
  assign t[37] = ~(t[44] ^ t[60]);
  assign t[380] = t[462] ^ x[112];
  assign t[381] = t[463] ^ x[111];
  assign t[382] = t[464] ^ x[115];
  assign t[383] = t[465] ^ x[114];
  assign t[384] = t[466] ^ x[118];
  assign t[385] = t[467] ^ x[117];
  assign t[386] = t[468] ^ x[121];
  assign t[387] = t[469] ^ x[120];
  assign t[388] = t[470] ^ x[124];
  assign t[389] = t[471] ^ x[123];
  assign t[38] = ~(t[61] | t[62]);
  assign t[390] = t[472] ^ x[127];
  assign t[391] = t[473] ^ x[126];
  assign t[392] = t[474] ^ x[130];
  assign t[393] = t[475] ^ x[129];
  assign t[394] = t[476] ^ x[133];
  assign t[395] = t[477] ^ x[132];
  assign t[396] = t[478] ^ x[136];
  assign t[397] = t[479] ^ x[135];
  assign t[398] = t[480] ^ x[139];
  assign t[399] = t[481] ^ x[138];
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[0]);
  assign t[401] = (x[0]);
  assign t[402] = (x[8]);
  assign t[403] = (x[8]);
  assign t[404] = (x[11]);
  assign t[405] = (x[11]);
  assign t[406] = (x[14]);
  assign t[407] = (x[14]);
  assign t[408] = (x[17]);
  assign t[409] = (x[17]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[20]);
  assign t[411] = (x[20]);
  assign t[412] = (x[23]);
  assign t[413] = (x[23]);
  assign t[414] = (x[26]);
  assign t[415] = (x[26]);
  assign t[416] = (x[29]);
  assign t[417] = (x[29]);
  assign t[418] = (x[34]);
  assign t[419] = (x[34]);
  assign t[41] = ~(t[201] | t[67]);
  assign t[420] = (x[37]);
  assign t[421] = (x[37]);
  assign t[422] = (x[40]);
  assign t[423] = (x[40]);
  assign t[424] = (x[43]);
  assign t[425] = (x[43]);
  assign t[426] = (x[46]);
  assign t[427] = (x[46]);
  assign t[428] = (x[51]);
  assign t[429] = (x[51]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[54]);
  assign t[431] = (x[54]);
  assign t[432] = (x[57]);
  assign t[433] = (x[57]);
  assign t[434] = (x[60]);
  assign t[435] = (x[60]);
  assign t[436] = (x[63]);
  assign t[437] = (x[63]);
  assign t[438] = (x[68]);
  assign t[439] = (x[68]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[71]);
  assign t[441] = (x[71]);
  assign t[442] = (x[74]);
  assign t[443] = (x[74]);
  assign t[444] = (x[79]);
  assign t[445] = (x[79]);
  assign t[446] = (x[82]);
  assign t[447] = (x[82]);
  assign t[448] = (x[85]);
  assign t[449] = (x[85]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[88]);
  assign t[451] = (x[88]);
  assign t[452] = (x[91]);
  assign t[453] = (x[91]);
  assign t[454] = (x[96]);
  assign t[455] = (x[96]);
  assign t[456] = (x[99]);
  assign t[457] = (x[99]);
  assign t[458] = (x[102]);
  assign t[459] = (x[102]);
  assign t[45] = ~(t[46] ^ t[74]);
  assign t[460] = (x[107]);
  assign t[461] = (x[107]);
  assign t[462] = (x[110]);
  assign t[463] = (x[110]);
  assign t[464] = (x[113]);
  assign t[465] = (x[113]);
  assign t[466] = (x[116]);
  assign t[467] = (x[116]);
  assign t[468] = (x[119]);
  assign t[469] = (x[119]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[122]);
  assign t[471] = (x[122]);
  assign t[472] = (x[125]);
  assign t[473] = (x[125]);
  assign t[474] = (x[128]);
  assign t[475] = (x[128]);
  assign t[476] = (x[131]);
  assign t[477] = (x[131]);
  assign t[478] = (x[134]);
  assign t[479] = (x[134]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[137]);
  assign t[481] = (x[137]);
  assign t[48] = ~(t[198]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[82]);
  assign t[51] = ~(t[197] | t[83]);
  assign t[52] = t[79] & t[196];
  assign t[53] = ~(t[202]);
  assign t[54] = ~(t[203]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[198] ? x[33] : x[32];
  assign t[57] = t[86] | t[87];
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[204] | t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[61] = ~(t[93] | t[94]);
  assign t[62] = ~(t[205] | t[95]);
  assign t[63] = ~(t[96] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[206]);
  assign t[66] = ~(t[207]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[208] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[50] : x[49];
  assign t[71] = ~(t[105] & t[106]);
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[209] | t[109]);
  assign t[74] = ~(t[110] ^ t[111]);
  assign t[75] = ~(t[112] | t[113]);
  assign t[76] = ~(t[210] | t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[117] ^ t[118]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[196] ? t[121] : t[120];
  assign t[81] = ~(t[122] | t[123]);
  assign t[82] = ~(t[119] & t[124]);
  assign t[83] = ~(t[199]);
  assign t[84] = ~(t[211]);
  assign t[85] = ~(t[202] | t[203]);
  assign t[86] = ~(t[125] & t[32]);
  assign t[87] = ~(t[126] & t[127]);
  assign t[88] = ~(t[212]);
  assign t[89] = ~(t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[128] | t[129]);
  assign t[91] = t[198] ? x[67] : x[66];
  assign t[92] = ~(t[130] & t[131]);
  assign t[93] = ~(t[214]);
  assign t[94] = ~(t[215]);
  assign t[95] = ~(t[132] | t[133]);
  assign t[96] = ~(t[134] | t[135]);
  assign t[97] = ~(t[216] | t[136]);
  assign t[98] = t[198] ? x[78] : x[77];
  assign t[99] = ~(t[130] & t[137]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [139:0] x;
 output y;

 wire [481:0] t;
  assign t[0] = t[1] ? t[2] : t[195];
  assign t[100] = ~(t[217]);
  assign t[101] = ~(t[206] | t[207]);
  assign t[102] = ~(t[218]);
  assign t[103] = ~(t[219]);
  assign t[104] = ~(t[138] | t[139]);
  assign t[105] = ~(t[86] | t[140]);
  assign t[106] = ~(t[141] & t[142]);
  assign t[107] = ~(t[220]);
  assign t[108] = ~(t[221]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[145] ? x[95] : x[94];
  assign t[111] = t[146] | t[147];
  assign t[112] = ~(t[222]);
  assign t[113] = ~(t[223]);
  assign t[114] = ~(t[148] | t[149]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[224] | t[152]);
  assign t[117] = t[145] ? x[106] : x[105];
  assign t[118] = ~(t[153] & t[154]);
  assign t[119] = ~(t[198]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[155] & t[83]);
  assign t[121] = ~(t[156] & t[199]);
  assign t[122] = ~(t[119] | t[157]);
  assign t[123] = ~(t[79] | t[158]);
  assign t[124] = ~(t[159] & t[160]);
  assign t[125] = ~(t[161] & t[162]);
  assign t[126] = ~(t[163] | t[164]);
  assign t[127] = ~(t[165] | t[166]);
  assign t[128] = ~(t[225]);
  assign t[129] = ~(t[212] | t[213]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[163] | t[167]);
  assign t[131] = ~(t[168] | t[169]);
  assign t[132] = ~(t[226]);
  assign t[133] = ~(t[214] | t[215]);
  assign t[134] = ~(t[227]);
  assign t[135] = ~(t[228]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[166]);
  assign t[138] = ~(t[229]);
  assign t[139] = ~(t[218] | t[219]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[147] | t[164];
  assign t[141] = t[199] & t[161];
  assign t[142] = t[155] | t[156];
  assign t[143] = ~(t[230]);
  assign t[144] = ~(t[220] | t[221]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[173] & t[32]);
  assign t[147] = ~(t[79] | t[174]);
  assign t[148] = ~(t[231]);
  assign t[149] = ~(t[222] | t[223]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[232]);
  assign t[151] = ~(t[233]);
  assign t[152] = ~(t[175] | t[176]);
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[177] | t[147]);
  assign t[155] = ~(x[4] | t[197]);
  assign t[156] = x[4] & t[197];
  assign t[157] = t[196] ? t[120] : t[178];
  assign t[158] = t[196] ? t[180] : t[179];
  assign t[159] = ~(x[4] & t[181]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[199] & t[182]);
  assign t[161] = ~(t[119] | t[196]);
  assign t[162] = ~(t[160] & t[179]);
  assign t[163] = ~(t[79] | t[183]);
  assign t[164] = ~(t[79] | t[184]);
  assign t[165] = ~(t[79] | t[185]);
  assign t[166] = ~(t[79] | t[186]);
  assign t[167] = ~(t[187] & t[106]);
  assign t[168] = ~(t[119] | t[188]);
  assign t[169] = t[164] | t[189];
  assign t[16] = ~(t[196] & t[197]);
  assign t[170] = ~(t[234]);
  assign t[171] = ~(t[227] | t[228]);
  assign t[172] = ~(t[79] | t[190]);
  assign t[173] = ~(t[191] | t[168]);
  assign t[174] = t[196] ? t[160] : t[159];
  assign t[175] = ~(t[235]);
  assign t[176] = ~(t[232] | t[233]);
  assign t[177] = ~(t[137]);
  assign t[178] = ~(t[156] & t[83]);
  assign t[179] = ~(x[4] & t[51]);
  assign t[17] = ~(t[198] & t[199]);
  assign t[180] = ~(t[182] & t[83]);
  assign t[181] = ~(t[197] | t[199]);
  assign t[182] = ~(x[4] | t[192]);
  assign t[183] = t[196] ? t[120] : t[121];
  assign t[184] = t[196] ? t[193] : t[178];
  assign t[185] = t[196] ? t[159] : t[160];
  assign t[186] = t[196] ? t[178] : t[193];
  assign t[187] = ~(t[49] | t[165]);
  assign t[188] = t[196] ? t[180] : t[159];
  assign t[189] = ~(t[125]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[196] ? t[179] : t[180];
  assign t[191] = ~(t[119] | t[194]);
  assign t[192] = ~(t[197]);
  assign t[193] = ~(t[155] & t[199]);
  assign t[194] = t[196] ? t[178] : t[120];
  assign t[195] = (t[236]);
  assign t[196] = (t[237]);
  assign t[197] = (t[238]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[6] : x[7];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = t[277] ^ x[2];
  assign t[237] = t[278] ^ x[10];
  assign t[238] = t[279] ^ x[13];
  assign t[239] = t[280] ^ x[16];
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = t[281] ^ x[19];
  assign t[241] = t[282] ^ x[22];
  assign t[242] = t[283] ^ x[25];
  assign t[243] = t[284] ^ x[28];
  assign t[244] = t[285] ^ x[31];
  assign t[245] = t[286] ^ x[36];
  assign t[246] = t[287] ^ x[39];
  assign t[247] = t[288] ^ x[42];
  assign t[248] = t[289] ^ x[45];
  assign t[249] = t[290] ^ x[48];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[53];
  assign t[251] = t[292] ^ x[56];
  assign t[252] = t[293] ^ x[59];
  assign t[253] = t[294] ^ x[62];
  assign t[254] = t[295] ^ x[65];
  assign t[255] = t[296] ^ x[70];
  assign t[256] = t[297] ^ x[73];
  assign t[257] = t[298] ^ x[76];
  assign t[258] = t[299] ^ x[81];
  assign t[259] = t[300] ^ x[84];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[87];
  assign t[261] = t[302] ^ x[90];
  assign t[262] = t[303] ^ x[93];
  assign t[263] = t[304] ^ x[98];
  assign t[264] = t[305] ^ x[101];
  assign t[265] = t[306] ^ x[104];
  assign t[266] = t[307] ^ x[109];
  assign t[267] = t[308] ^ x[112];
  assign t[268] = t[309] ^ x[115];
  assign t[269] = t[310] ^ x[118];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[121];
  assign t[271] = t[312] ^ x[124];
  assign t[272] = t[313] ^ x[127];
  assign t[273] = t[314] ^ x[130];
  assign t[274] = t[315] ^ x[133];
  assign t[275] = t[316] ^ x[136];
  assign t[276] = t[317] ^ x[139];
  assign t[277] = (t[318] & ~t[319]);
  assign t[278] = (t[320] & ~t[321]);
  assign t[279] = (t[322] & ~t[323]);
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = (t[324] & ~t[325]);
  assign t[281] = (t[326] & ~t[327]);
  assign t[282] = (t[328] & ~t[329]);
  assign t[283] = (t[330] & ~t[331]);
  assign t[284] = (t[332] & ~t[333]);
  assign t[285] = (t[334] & ~t[335]);
  assign t[286] = (t[336] & ~t[337]);
  assign t[287] = (t[338] & ~t[339]);
  assign t[288] = (t[340] & ~t[341]);
  assign t[289] = (t[342] & ~t[343]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[344] & ~t[345]);
  assign t[291] = (t[346] & ~t[347]);
  assign t[292] = (t[348] & ~t[349]);
  assign t[293] = (t[350] & ~t[351]);
  assign t[294] = (t[352] & ~t[353]);
  assign t[295] = (t[354] & ~t[355]);
  assign t[296] = (t[356] & ~t[357]);
  assign t[297] = (t[358] & ~t[359]);
  assign t[298] = (t[360] & ~t[361]);
  assign t[299] = (t[362] & ~t[363]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[364] & ~t[365]);
  assign t[301] = (t[366] & ~t[367]);
  assign t[302] = (t[368] & ~t[369]);
  assign t[303] = (t[370] & ~t[371]);
  assign t[304] = (t[372] & ~t[373]);
  assign t[305] = (t[374] & ~t[375]);
  assign t[306] = (t[376] & ~t[377]);
  assign t[307] = (t[378] & ~t[379]);
  assign t[308] = (t[380] & ~t[381]);
  assign t[309] = (t[382] & ~t[383]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[384] & ~t[385]);
  assign t[311] = (t[386] & ~t[387]);
  assign t[312] = (t[388] & ~t[389]);
  assign t[313] = (t[390] & ~t[391]);
  assign t[314] = (t[392] & ~t[393]);
  assign t[315] = (t[394] & ~t[395]);
  assign t[316] = (t[396] & ~t[397]);
  assign t[317] = (t[398] & ~t[399]);
  assign t[318] = t[400] ^ x[2];
  assign t[319] = t[401] ^ x[1];
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = t[402] ^ x[10];
  assign t[321] = t[403] ^ x[9];
  assign t[322] = t[404] ^ x[13];
  assign t[323] = t[405] ^ x[12];
  assign t[324] = t[406] ^ x[16];
  assign t[325] = t[407] ^ x[15];
  assign t[326] = t[408] ^ x[19];
  assign t[327] = t[409] ^ x[18];
  assign t[328] = t[410] ^ x[22];
  assign t[329] = t[411] ^ x[21];
  assign t[32] = ~(t[51] & t[52]);
  assign t[330] = t[412] ^ x[25];
  assign t[331] = t[413] ^ x[24];
  assign t[332] = t[414] ^ x[28];
  assign t[333] = t[415] ^ x[27];
  assign t[334] = t[416] ^ x[31];
  assign t[335] = t[417] ^ x[30];
  assign t[336] = t[418] ^ x[36];
  assign t[337] = t[419] ^ x[35];
  assign t[338] = t[420] ^ x[39];
  assign t[339] = t[421] ^ x[38];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[42];
  assign t[341] = t[423] ^ x[41];
  assign t[342] = t[424] ^ x[45];
  assign t[343] = t[425] ^ x[44];
  assign t[344] = t[426] ^ x[48];
  assign t[345] = t[427] ^ x[47];
  assign t[346] = t[428] ^ x[53];
  assign t[347] = t[429] ^ x[52];
  assign t[348] = t[430] ^ x[56];
  assign t[349] = t[431] ^ x[55];
  assign t[34] = ~(t[200] | t[55]);
  assign t[350] = t[432] ^ x[59];
  assign t[351] = t[433] ^ x[58];
  assign t[352] = t[434] ^ x[62];
  assign t[353] = t[435] ^ x[61];
  assign t[354] = t[436] ^ x[65];
  assign t[355] = t[437] ^ x[64];
  assign t[356] = t[438] ^ x[70];
  assign t[357] = t[439] ^ x[69];
  assign t[358] = t[440] ^ x[73];
  assign t[359] = t[441] ^ x[72];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[76];
  assign t[361] = t[443] ^ x[75];
  assign t[362] = t[444] ^ x[81];
  assign t[363] = t[445] ^ x[80];
  assign t[364] = t[446] ^ x[84];
  assign t[365] = t[447] ^ x[83];
  assign t[366] = t[448] ^ x[87];
  assign t[367] = t[449] ^ x[86];
  assign t[368] = t[450] ^ x[90];
  assign t[369] = t[451] ^ x[89];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[93];
  assign t[371] = t[453] ^ x[92];
  assign t[372] = t[454] ^ x[98];
  assign t[373] = t[455] ^ x[97];
  assign t[374] = t[456] ^ x[101];
  assign t[375] = t[457] ^ x[100];
  assign t[376] = t[458] ^ x[104];
  assign t[377] = t[459] ^ x[103];
  assign t[378] = t[460] ^ x[109];
  assign t[379] = t[461] ^ x[108];
  assign t[37] = ~(t[44] ^ t[60]);
  assign t[380] = t[462] ^ x[112];
  assign t[381] = t[463] ^ x[111];
  assign t[382] = t[464] ^ x[115];
  assign t[383] = t[465] ^ x[114];
  assign t[384] = t[466] ^ x[118];
  assign t[385] = t[467] ^ x[117];
  assign t[386] = t[468] ^ x[121];
  assign t[387] = t[469] ^ x[120];
  assign t[388] = t[470] ^ x[124];
  assign t[389] = t[471] ^ x[123];
  assign t[38] = ~(t[61] | t[62]);
  assign t[390] = t[472] ^ x[127];
  assign t[391] = t[473] ^ x[126];
  assign t[392] = t[474] ^ x[130];
  assign t[393] = t[475] ^ x[129];
  assign t[394] = t[476] ^ x[133];
  assign t[395] = t[477] ^ x[132];
  assign t[396] = t[478] ^ x[136];
  assign t[397] = t[479] ^ x[135];
  assign t[398] = t[480] ^ x[139];
  assign t[399] = t[481] ^ x[138];
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[0]);
  assign t[401] = (x[0]);
  assign t[402] = (x[8]);
  assign t[403] = (x[8]);
  assign t[404] = (x[11]);
  assign t[405] = (x[11]);
  assign t[406] = (x[14]);
  assign t[407] = (x[14]);
  assign t[408] = (x[17]);
  assign t[409] = (x[17]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[20]);
  assign t[411] = (x[20]);
  assign t[412] = (x[23]);
  assign t[413] = (x[23]);
  assign t[414] = (x[26]);
  assign t[415] = (x[26]);
  assign t[416] = (x[29]);
  assign t[417] = (x[29]);
  assign t[418] = (x[34]);
  assign t[419] = (x[34]);
  assign t[41] = ~(t[201] | t[67]);
  assign t[420] = (x[37]);
  assign t[421] = (x[37]);
  assign t[422] = (x[40]);
  assign t[423] = (x[40]);
  assign t[424] = (x[43]);
  assign t[425] = (x[43]);
  assign t[426] = (x[46]);
  assign t[427] = (x[46]);
  assign t[428] = (x[51]);
  assign t[429] = (x[51]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[54]);
  assign t[431] = (x[54]);
  assign t[432] = (x[57]);
  assign t[433] = (x[57]);
  assign t[434] = (x[60]);
  assign t[435] = (x[60]);
  assign t[436] = (x[63]);
  assign t[437] = (x[63]);
  assign t[438] = (x[68]);
  assign t[439] = (x[68]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[71]);
  assign t[441] = (x[71]);
  assign t[442] = (x[74]);
  assign t[443] = (x[74]);
  assign t[444] = (x[79]);
  assign t[445] = (x[79]);
  assign t[446] = (x[82]);
  assign t[447] = (x[82]);
  assign t[448] = (x[85]);
  assign t[449] = (x[85]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[88]);
  assign t[451] = (x[88]);
  assign t[452] = (x[91]);
  assign t[453] = (x[91]);
  assign t[454] = (x[96]);
  assign t[455] = (x[96]);
  assign t[456] = (x[99]);
  assign t[457] = (x[99]);
  assign t[458] = (x[102]);
  assign t[459] = (x[102]);
  assign t[45] = ~(t[46] ^ t[74]);
  assign t[460] = (x[107]);
  assign t[461] = (x[107]);
  assign t[462] = (x[110]);
  assign t[463] = (x[110]);
  assign t[464] = (x[113]);
  assign t[465] = (x[113]);
  assign t[466] = (x[116]);
  assign t[467] = (x[116]);
  assign t[468] = (x[119]);
  assign t[469] = (x[119]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[122]);
  assign t[471] = (x[122]);
  assign t[472] = (x[125]);
  assign t[473] = (x[125]);
  assign t[474] = (x[128]);
  assign t[475] = (x[128]);
  assign t[476] = (x[131]);
  assign t[477] = (x[131]);
  assign t[478] = (x[134]);
  assign t[479] = (x[134]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[137]);
  assign t[481] = (x[137]);
  assign t[48] = ~(t[198]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[82]);
  assign t[51] = ~(t[197] | t[83]);
  assign t[52] = t[79] & t[196];
  assign t[53] = ~(t[202]);
  assign t[54] = ~(t[203]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[198] ? x[33] : x[32];
  assign t[57] = t[86] | t[87];
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[204] | t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[61] = ~(t[93] | t[94]);
  assign t[62] = ~(t[205] | t[95]);
  assign t[63] = ~(t[96] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[206]);
  assign t[66] = ~(t[207]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[208] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[50] : x[49];
  assign t[71] = ~(t[105] & t[106]);
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[209] | t[109]);
  assign t[74] = ~(t[110] ^ t[111]);
  assign t[75] = ~(t[112] | t[113]);
  assign t[76] = ~(t[210] | t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[117] ^ t[118]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[196] ? t[121] : t[120];
  assign t[81] = ~(t[122] | t[123]);
  assign t[82] = ~(t[119] & t[124]);
  assign t[83] = ~(t[199]);
  assign t[84] = ~(t[211]);
  assign t[85] = ~(t[202] | t[203]);
  assign t[86] = ~(t[125] & t[32]);
  assign t[87] = ~(t[126] & t[127]);
  assign t[88] = ~(t[212]);
  assign t[89] = ~(t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[128] | t[129]);
  assign t[91] = t[198] ? x[67] : x[66];
  assign t[92] = ~(t[130] & t[131]);
  assign t[93] = ~(t[214]);
  assign t[94] = ~(t[215]);
  assign t[95] = ~(t[132] | t[133]);
  assign t[96] = ~(t[134] | t[135]);
  assign t[97] = ~(t[216] | t[136]);
  assign t[98] = t[198] ? x[78] : x[77];
  assign t[99] = ~(t[130] & t[137]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind206(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[49];
  assign t[139] = t[171] ^ x[52];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[57];
  assign t[141] = t[173] ^ x[60];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[49];
  assign t[215] = t[279] ^ x[48];
  assign t[216] = t[280] ^ x[52];
  assign t[217] = t[281] ^ x[51];
  assign t[218] = t[282] ^ x[57];
  assign t[219] = t[283] ^ x[56];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[60];
  assign t[221] = t[285] ^ x[59];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[47]);
  assign t[279] = (x[47]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[50]);
  assign t[282] = (x[55]);
  assign t[283] = (x[55]);
  assign t[284] = (x[58]);
  assign t[285] = (x[58]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[97] ? x[27] : x[26];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[50];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[43];
  assign t[37] = ~(t[101] & t[54]);
  assign t[38] = ~(t[102] & t[55]);
  assign t[39] = t[18] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[56] & t[57]);
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[41];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[65]);
  assign t[47] = ~(t[104] & t[66]);
  assign t[48] = ~(t[105] & t[67]);
  assign t[49] = t[97] ? x[46] : x[45];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[72] ? x[54] : x[53];
  assign t[54] = ~(t[108]);
  assign t[55] = ~(t[108] & t[73]);
  assign t[56] = ~(t[109] & t[74]);
  assign t[57] = ~(t[110] & t[75]);
  assign t[58] = ~(t[111] & t[76]);
  assign t[59] = ~(t[112] & t[77]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[78] ? x[71] : x[70];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[113] & t[81]);
  assign t[63] = ~(t[114] & t[82]);
  assign t[64] = t[78] ? x[79] : x[78];
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[115]);
  assign t[67] = ~(t[115] & t[83]);
  assign t[68] = ~(t[116] & t[84]);
  assign t[69] = ~(t[117] & t[85]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[118]);
  assign t[71] = ~(t[118] & t[86]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[101]);
  assign t[74] = ~(t[119]);
  assign t[75] = ~(t[119] & t[87]);
  assign t[76] = ~(t[120]);
  assign t[77] = ~(t[120] & t[88]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122] & t[90]);
  assign t[81] = ~(t[123]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[124]);
  assign t[85] = ~(t[124] & t[92]);
  assign t[86] = ~(t[106]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[125]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] & t[93]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[121]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[49];
  assign t[139] = t[171] ^ x[52];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[57];
  assign t[141] = t[173] ^ x[60];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[49];
  assign t[215] = t[279] ^ x[48];
  assign t[216] = t[280] ^ x[52];
  assign t[217] = t[281] ^ x[51];
  assign t[218] = t[282] ^ x[57];
  assign t[219] = t[283] ^ x[56];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[60];
  assign t[221] = t[285] ^ x[59];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[47]);
  assign t[279] = (x[47]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[50]);
  assign t[282] = (x[55]);
  assign t[283] = (x[55]);
  assign t[284] = (x[58]);
  assign t[285] = (x[58]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[97] ? x[27] : x[26];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[50];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[43];
  assign t[37] = ~(t[101] & t[54]);
  assign t[38] = ~(t[102] & t[55]);
  assign t[39] = t[18] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[56] & t[57]);
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[41];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[65]);
  assign t[47] = ~(t[104] & t[66]);
  assign t[48] = ~(t[105] & t[67]);
  assign t[49] = t[97] ? x[46] : x[45];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[72] ? x[54] : x[53];
  assign t[54] = ~(t[108]);
  assign t[55] = ~(t[108] & t[73]);
  assign t[56] = ~(t[109] & t[74]);
  assign t[57] = ~(t[110] & t[75]);
  assign t[58] = ~(t[111] & t[76]);
  assign t[59] = ~(t[112] & t[77]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[78] ? x[71] : x[70];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[113] & t[81]);
  assign t[63] = ~(t[114] & t[82]);
  assign t[64] = t[78] ? x[79] : x[78];
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[115]);
  assign t[67] = ~(t[115] & t[83]);
  assign t[68] = ~(t[116] & t[84]);
  assign t[69] = ~(t[117] & t[85]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[118]);
  assign t[71] = ~(t[118] & t[86]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[101]);
  assign t[74] = ~(t[119]);
  assign t[75] = ~(t[119] & t[87]);
  assign t[76] = ~(t[120]);
  assign t[77] = ~(t[120] & t[88]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122] & t[90]);
  assign t[81] = ~(t[123]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[124]);
  assign t[85] = ~(t[124] & t[92]);
  assign t[86] = ~(t[106]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[125]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] & t[93]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[121]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = ~(t[114]);
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[114] ? x[24] : x[23];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[41];
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = t[18] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[67] & t[68]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = ~(t[71] & t[120]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[114] ? x[40] : x[39];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[121]);
  assign t[54] = t[18] ? x[45] : x[44];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[77] & t[78]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[124]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[125]);
  assign t[62] = t[85] ? x[59] : x[58];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[126]);
  assign t[65] = t[85] ? x[64] : x[63];
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[91] & t[92]);
  assign t[72] = ~(t[93] & t[94]);
  assign t[73] = ~(t[95] & t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[96] & t[97]);
  assign t[77] = ~(t[123] & t[122]);
  assign t[78] = ~(t[133]);
  assign t[79] = ~(t[134]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[135]);
  assign t[81] = ~(t[98] & t[99]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[100] & t[101]);
  assign t[85] = ~(t[25]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = ~(t[114]);
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[114] ? x[24] : x[23];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[41];
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = t[18] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[67] & t[68]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = ~(t[71] & t[120]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[114] ? x[40] : x[39];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[121]);
  assign t[54] = t[18] ? x[45] : x[44];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[77] & t[78]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[124]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[125]);
  assign t[62] = t[85] ? x[59] : x[58];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[126]);
  assign t[65] = t[85] ? x[64] : x[63];
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[91] & t[92]);
  assign t[72] = ~(t[93] & t[94]);
  assign t[73] = ~(t[95] & t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[96] & t[97]);
  assign t[77] = ~(t[123] & t[122]);
  assign t[78] = ~(t[133]);
  assign t[79] = ~(t[134]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[135]);
  assign t[81] = ~(t[98] & t[99]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[100] & t[101]);
  assign t[85] = ~(t[25]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [139:0] x;
 output y;

 wire [388:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[2];
  assign t[144] = t[185] ^ x[10];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[27];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[32];
  assign t[151] = t[192] ^ x[35];
  assign t[152] = t[193] ^ x[38];
  assign t[153] = t[194] ^ x[43];
  assign t[154] = t[195] ^ x[48];
  assign t[155] = t[196] ^ x[51];
  assign t[156] = t[197] ^ x[54];
  assign t[157] = t[198] ^ x[57];
  assign t[158] = t[199] ^ x[62];
  assign t[159] = t[200] ^ x[67];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[70];
  assign t[161] = t[202] ^ x[73];
  assign t[162] = t[203] ^ x[76];
  assign t[163] = t[204] ^ x[79];
  assign t[164] = t[205] ^ x[82];
  assign t[165] = t[206] ^ x[85];
  assign t[166] = t[207] ^ x[88];
  assign t[167] = t[208] ^ x[91];
  assign t[168] = t[209] ^ x[94];
  assign t[169] = t[210] ^ x[97];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[100];
  assign t[171] = t[212] ^ x[103];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[109];
  assign t[174] = t[215] ^ x[112];
  assign t[175] = t[216] ^ x[115];
  assign t[176] = t[217] ^ x[118];
  assign t[177] = t[218] ^ x[121];
  assign t[178] = t[219] ^ x[124];
  assign t[179] = t[220] ^ x[127];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[130];
  assign t[181] = t[222] ^ x[133];
  assign t[182] = t[223] ^ x[136];
  assign t[183] = t[224] ^ x[139];
  assign t[184] = (t[225] & ~t[226]);
  assign t[185] = (t[227] & ~t[228]);
  assign t[186] = (t[229] & ~t[230]);
  assign t[187] = (t[231] & ~t[232]);
  assign t[188] = (t[233] & ~t[234]);
  assign t[189] = (t[235] & ~t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[237] & ~t[238]);
  assign t[191] = (t[239] & ~t[240]);
  assign t[192] = (t[241] & ~t[242]);
  assign t[193] = (t[243] & ~t[244]);
  assign t[194] = (t[245] & ~t[246]);
  assign t[195] = (t[247] & ~t[248]);
  assign t[196] = (t[249] & ~t[250]);
  assign t[197] = (t[251] & ~t[252]);
  assign t[198] = (t[253] & ~t[254]);
  assign t[199] = (t[255] & ~t[256]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[257] & ~t[258]);
  assign t[201] = (t[259] & ~t[260]);
  assign t[202] = (t[261] & ~t[262]);
  assign t[203] = (t[263] & ~t[264]);
  assign t[204] = (t[265] & ~t[266]);
  assign t[205] = (t[267] & ~t[268]);
  assign t[206] = (t[269] & ~t[270]);
  assign t[207] = (t[271] & ~t[272]);
  assign t[208] = (t[273] & ~t[274]);
  assign t[209] = (t[275] & ~t[276]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[277] & ~t[278]);
  assign t[211] = (t[279] & ~t[280]);
  assign t[212] = (t[281] & ~t[282]);
  assign t[213] = (t[283] & ~t[284]);
  assign t[214] = (t[285] & ~t[286]);
  assign t[215] = (t[287] & ~t[288]);
  assign t[216] = (t[289] & ~t[290]);
  assign t[217] = (t[291] & ~t[292]);
  assign t[218] = (t[293] & ~t[294]);
  assign t[219] = (t[295] & ~t[296]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[297] & ~t[298]);
  assign t[221] = (t[299] & ~t[300]);
  assign t[222] = (t[301] & ~t[302]);
  assign t[223] = (t[303] & ~t[304]);
  assign t[224] = (t[305] & ~t[306]);
  assign t[225] = t[307] ^ x[2];
  assign t[226] = t[308] ^ x[1];
  assign t[227] = t[309] ^ x[10];
  assign t[228] = t[310] ^ x[9];
  assign t[229] = t[311] ^ x[13];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[312] ^ x[12];
  assign t[231] = t[313] ^ x[16];
  assign t[232] = t[314] ^ x[15];
  assign t[233] = t[315] ^ x[19];
  assign t[234] = t[316] ^ x[18];
  assign t[235] = t[317] ^ x[22];
  assign t[236] = t[318] ^ x[21];
  assign t[237] = t[319] ^ x[27];
  assign t[238] = t[320] ^ x[26];
  assign t[239] = t[321] ^ x[32];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[31];
  assign t[241] = t[323] ^ x[35];
  assign t[242] = t[324] ^ x[34];
  assign t[243] = t[325] ^ x[38];
  assign t[244] = t[326] ^ x[37];
  assign t[245] = t[327] ^ x[43];
  assign t[246] = t[328] ^ x[42];
  assign t[247] = t[329] ^ x[48];
  assign t[248] = t[330] ^ x[47];
  assign t[249] = t[331] ^ x[51];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[50];
  assign t[251] = t[333] ^ x[54];
  assign t[252] = t[334] ^ x[53];
  assign t[253] = t[335] ^ x[57];
  assign t[254] = t[336] ^ x[56];
  assign t[255] = t[337] ^ x[62];
  assign t[256] = t[338] ^ x[61];
  assign t[257] = t[339] ^ x[67];
  assign t[258] = t[340] ^ x[66];
  assign t[259] = t[341] ^ x[70];
  assign t[25] = ~(t[105]);
  assign t[260] = t[342] ^ x[69];
  assign t[261] = t[343] ^ x[73];
  assign t[262] = t[344] ^ x[72];
  assign t[263] = t[345] ^ x[76];
  assign t[264] = t[346] ^ x[75];
  assign t[265] = t[347] ^ x[79];
  assign t[266] = t[348] ^ x[78];
  assign t[267] = t[349] ^ x[82];
  assign t[268] = t[350] ^ x[81];
  assign t[269] = t[351] ^ x[85];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[84];
  assign t[271] = t[353] ^ x[88];
  assign t[272] = t[354] ^ x[87];
  assign t[273] = t[355] ^ x[91];
  assign t[274] = t[356] ^ x[90];
  assign t[275] = t[357] ^ x[94];
  assign t[276] = t[358] ^ x[93];
  assign t[277] = t[359] ^ x[97];
  assign t[278] = t[360] ^ x[96];
  assign t[279] = t[361] ^ x[100];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[99];
  assign t[281] = t[363] ^ x[103];
  assign t[282] = t[364] ^ x[102];
  assign t[283] = t[365] ^ x[106];
  assign t[284] = t[366] ^ x[105];
  assign t[285] = t[367] ^ x[109];
  assign t[286] = t[368] ^ x[108];
  assign t[287] = t[369] ^ x[112];
  assign t[288] = t[370] ^ x[111];
  assign t[289] = t[371] ^ x[115];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[114];
  assign t[291] = t[373] ^ x[118];
  assign t[292] = t[374] ^ x[117];
  assign t[293] = t[375] ^ x[121];
  assign t[294] = t[376] ^ x[120];
  assign t[295] = t[377] ^ x[124];
  assign t[296] = t[378] ^ x[123];
  assign t[297] = t[379] ^ x[127];
  assign t[298] = t[380] ^ x[126];
  assign t[299] = t[381] ^ x[130];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[129];
  assign t[301] = t[383] ^ x[133];
  assign t[302] = t[384] ^ x[132];
  assign t[303] = t[385] ^ x[136];
  assign t[304] = t[386] ^ x[135];
  assign t[305] = t[387] ^ x[139];
  assign t[306] = t[388] ^ x[138];
  assign t[307] = (x[0]);
  assign t[308] = (x[0]);
  assign t[309] = (x[8]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[11]);
  assign t[312] = (x[11]);
  assign t[313] = (x[14]);
  assign t[314] = (x[14]);
  assign t[315] = (x[17]);
  assign t[316] = (x[17]);
  assign t[317] = (x[20]);
  assign t[318] = (x[20]);
  assign t[319] = (x[25]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[25]);
  assign t[321] = (x[30]);
  assign t[322] = (x[30]);
  assign t[323] = (x[33]);
  assign t[324] = (x[33]);
  assign t[325] = (x[36]);
  assign t[326] = (x[36]);
  assign t[327] = (x[41]);
  assign t[328] = (x[41]);
  assign t[329] = (x[46]);
  assign t[32] = t[105] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[49]);
  assign t[332] = (x[49]);
  assign t[333] = (x[52]);
  assign t[334] = (x[52]);
  assign t[335] = (x[55]);
  assign t[336] = (x[55]);
  assign t[337] = (x[60]);
  assign t[338] = (x[60]);
  assign t[339] = (x[65]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[68]);
  assign t[342] = (x[68]);
  assign t[343] = (x[71]);
  assign t[344] = (x[71]);
  assign t[345] = (x[74]);
  assign t[346] = (x[74]);
  assign t[347] = (x[77]);
  assign t[348] = (x[77]);
  assign t[349] = (x[80]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[80]);
  assign t[351] = (x[83]);
  assign t[352] = (x[83]);
  assign t[353] = (x[86]);
  assign t[354] = (x[86]);
  assign t[355] = (x[89]);
  assign t[356] = (x[89]);
  assign t[357] = (x[92]);
  assign t[358] = (x[92]);
  assign t[359] = (x[95]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[95]);
  assign t[361] = (x[98]);
  assign t[362] = (x[98]);
  assign t[363] = (x[101]);
  assign t[364] = (x[101]);
  assign t[365] = (x[104]);
  assign t[366] = (x[104]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[54] ^ t[41];
  assign t[370] = (x[110]);
  assign t[371] = (x[113]);
  assign t[372] = (x[113]);
  assign t[373] = (x[116]);
  assign t[374] = (x[116]);
  assign t[375] = (x[119]);
  assign t[376] = (x[119]);
  assign t[377] = (x[122]);
  assign t[378] = (x[122]);
  assign t[379] = (x[125]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[128]);
  assign t[382] = (x[128]);
  assign t[383] = (x[131]);
  assign t[384] = (x[131]);
  assign t[385] = (x[134]);
  assign t[386] = (x[134]);
  assign t[387] = (x[137]);
  assign t[388] = (x[137]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[18] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[67] | t[45]);
  assign t[48] = ~(t[68] & t[69]);
  assign t[49] = t[70] | t[111];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[105] ? x[40] : x[39];
  assign t[51] = ~(t[71] & t[72]);
  assign t[52] = ~(t[73] & t[74]);
  assign t[53] = t[75] | t[112];
  assign t[54] = t[76] ? x[45] : x[44];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = t[80] | t[115];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[116];
  assign t[62] = t[76] ? x[59] : x[58];
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = t[86] | t[117];
  assign t[65] = t[76] ? x[64] : x[63];
  assign t[66] = ~(t[87] & t[88]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = t[92] | t[121];
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[93] | t[73]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind211(x, y);
 input [139:0] x;
 output y;

 wire [388:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[6] : x[7];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[2];
  assign t[144] = t[185] ^ x[10];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[27];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[32];
  assign t[151] = t[192] ^ x[35];
  assign t[152] = t[193] ^ x[38];
  assign t[153] = t[194] ^ x[43];
  assign t[154] = t[195] ^ x[48];
  assign t[155] = t[196] ^ x[51];
  assign t[156] = t[197] ^ x[54];
  assign t[157] = t[198] ^ x[57];
  assign t[158] = t[199] ^ x[62];
  assign t[159] = t[200] ^ x[67];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[70];
  assign t[161] = t[202] ^ x[73];
  assign t[162] = t[203] ^ x[76];
  assign t[163] = t[204] ^ x[79];
  assign t[164] = t[205] ^ x[82];
  assign t[165] = t[206] ^ x[85];
  assign t[166] = t[207] ^ x[88];
  assign t[167] = t[208] ^ x[91];
  assign t[168] = t[209] ^ x[94];
  assign t[169] = t[210] ^ x[97];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[100];
  assign t[171] = t[212] ^ x[103];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[109];
  assign t[174] = t[215] ^ x[112];
  assign t[175] = t[216] ^ x[115];
  assign t[176] = t[217] ^ x[118];
  assign t[177] = t[218] ^ x[121];
  assign t[178] = t[219] ^ x[124];
  assign t[179] = t[220] ^ x[127];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[130];
  assign t[181] = t[222] ^ x[133];
  assign t[182] = t[223] ^ x[136];
  assign t[183] = t[224] ^ x[139];
  assign t[184] = (t[225] & ~t[226]);
  assign t[185] = (t[227] & ~t[228]);
  assign t[186] = (t[229] & ~t[230]);
  assign t[187] = (t[231] & ~t[232]);
  assign t[188] = (t[233] & ~t[234]);
  assign t[189] = (t[235] & ~t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[237] & ~t[238]);
  assign t[191] = (t[239] & ~t[240]);
  assign t[192] = (t[241] & ~t[242]);
  assign t[193] = (t[243] & ~t[244]);
  assign t[194] = (t[245] & ~t[246]);
  assign t[195] = (t[247] & ~t[248]);
  assign t[196] = (t[249] & ~t[250]);
  assign t[197] = (t[251] & ~t[252]);
  assign t[198] = (t[253] & ~t[254]);
  assign t[199] = (t[255] & ~t[256]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[257] & ~t[258]);
  assign t[201] = (t[259] & ~t[260]);
  assign t[202] = (t[261] & ~t[262]);
  assign t[203] = (t[263] & ~t[264]);
  assign t[204] = (t[265] & ~t[266]);
  assign t[205] = (t[267] & ~t[268]);
  assign t[206] = (t[269] & ~t[270]);
  assign t[207] = (t[271] & ~t[272]);
  assign t[208] = (t[273] & ~t[274]);
  assign t[209] = (t[275] & ~t[276]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[277] & ~t[278]);
  assign t[211] = (t[279] & ~t[280]);
  assign t[212] = (t[281] & ~t[282]);
  assign t[213] = (t[283] & ~t[284]);
  assign t[214] = (t[285] & ~t[286]);
  assign t[215] = (t[287] & ~t[288]);
  assign t[216] = (t[289] & ~t[290]);
  assign t[217] = (t[291] & ~t[292]);
  assign t[218] = (t[293] & ~t[294]);
  assign t[219] = (t[295] & ~t[296]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[297] & ~t[298]);
  assign t[221] = (t[299] & ~t[300]);
  assign t[222] = (t[301] & ~t[302]);
  assign t[223] = (t[303] & ~t[304]);
  assign t[224] = (t[305] & ~t[306]);
  assign t[225] = t[307] ^ x[2];
  assign t[226] = t[308] ^ x[1];
  assign t[227] = t[309] ^ x[10];
  assign t[228] = t[310] ^ x[9];
  assign t[229] = t[311] ^ x[13];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[312] ^ x[12];
  assign t[231] = t[313] ^ x[16];
  assign t[232] = t[314] ^ x[15];
  assign t[233] = t[315] ^ x[19];
  assign t[234] = t[316] ^ x[18];
  assign t[235] = t[317] ^ x[22];
  assign t[236] = t[318] ^ x[21];
  assign t[237] = t[319] ^ x[27];
  assign t[238] = t[320] ^ x[26];
  assign t[239] = t[321] ^ x[32];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[31];
  assign t[241] = t[323] ^ x[35];
  assign t[242] = t[324] ^ x[34];
  assign t[243] = t[325] ^ x[38];
  assign t[244] = t[326] ^ x[37];
  assign t[245] = t[327] ^ x[43];
  assign t[246] = t[328] ^ x[42];
  assign t[247] = t[329] ^ x[48];
  assign t[248] = t[330] ^ x[47];
  assign t[249] = t[331] ^ x[51];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[50];
  assign t[251] = t[333] ^ x[54];
  assign t[252] = t[334] ^ x[53];
  assign t[253] = t[335] ^ x[57];
  assign t[254] = t[336] ^ x[56];
  assign t[255] = t[337] ^ x[62];
  assign t[256] = t[338] ^ x[61];
  assign t[257] = t[339] ^ x[67];
  assign t[258] = t[340] ^ x[66];
  assign t[259] = t[341] ^ x[70];
  assign t[25] = ~(t[105]);
  assign t[260] = t[342] ^ x[69];
  assign t[261] = t[343] ^ x[73];
  assign t[262] = t[344] ^ x[72];
  assign t[263] = t[345] ^ x[76];
  assign t[264] = t[346] ^ x[75];
  assign t[265] = t[347] ^ x[79];
  assign t[266] = t[348] ^ x[78];
  assign t[267] = t[349] ^ x[82];
  assign t[268] = t[350] ^ x[81];
  assign t[269] = t[351] ^ x[85];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[84];
  assign t[271] = t[353] ^ x[88];
  assign t[272] = t[354] ^ x[87];
  assign t[273] = t[355] ^ x[91];
  assign t[274] = t[356] ^ x[90];
  assign t[275] = t[357] ^ x[94];
  assign t[276] = t[358] ^ x[93];
  assign t[277] = t[359] ^ x[97];
  assign t[278] = t[360] ^ x[96];
  assign t[279] = t[361] ^ x[100];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[99];
  assign t[281] = t[363] ^ x[103];
  assign t[282] = t[364] ^ x[102];
  assign t[283] = t[365] ^ x[106];
  assign t[284] = t[366] ^ x[105];
  assign t[285] = t[367] ^ x[109];
  assign t[286] = t[368] ^ x[108];
  assign t[287] = t[369] ^ x[112];
  assign t[288] = t[370] ^ x[111];
  assign t[289] = t[371] ^ x[115];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[114];
  assign t[291] = t[373] ^ x[118];
  assign t[292] = t[374] ^ x[117];
  assign t[293] = t[375] ^ x[121];
  assign t[294] = t[376] ^ x[120];
  assign t[295] = t[377] ^ x[124];
  assign t[296] = t[378] ^ x[123];
  assign t[297] = t[379] ^ x[127];
  assign t[298] = t[380] ^ x[126];
  assign t[299] = t[381] ^ x[130];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[129];
  assign t[301] = t[383] ^ x[133];
  assign t[302] = t[384] ^ x[132];
  assign t[303] = t[385] ^ x[136];
  assign t[304] = t[386] ^ x[135];
  assign t[305] = t[387] ^ x[139];
  assign t[306] = t[388] ^ x[138];
  assign t[307] = (x[0]);
  assign t[308] = (x[0]);
  assign t[309] = (x[8]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[11]);
  assign t[312] = (x[11]);
  assign t[313] = (x[14]);
  assign t[314] = (x[14]);
  assign t[315] = (x[17]);
  assign t[316] = (x[17]);
  assign t[317] = (x[20]);
  assign t[318] = (x[20]);
  assign t[319] = (x[25]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[25]);
  assign t[321] = (x[30]);
  assign t[322] = (x[30]);
  assign t[323] = (x[33]);
  assign t[324] = (x[33]);
  assign t[325] = (x[36]);
  assign t[326] = (x[36]);
  assign t[327] = (x[41]);
  assign t[328] = (x[41]);
  assign t[329] = (x[46]);
  assign t[32] = t[105] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[49]);
  assign t[332] = (x[49]);
  assign t[333] = (x[52]);
  assign t[334] = (x[52]);
  assign t[335] = (x[55]);
  assign t[336] = (x[55]);
  assign t[337] = (x[60]);
  assign t[338] = (x[60]);
  assign t[339] = (x[65]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[68]);
  assign t[342] = (x[68]);
  assign t[343] = (x[71]);
  assign t[344] = (x[71]);
  assign t[345] = (x[74]);
  assign t[346] = (x[74]);
  assign t[347] = (x[77]);
  assign t[348] = (x[77]);
  assign t[349] = (x[80]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[80]);
  assign t[351] = (x[83]);
  assign t[352] = (x[83]);
  assign t[353] = (x[86]);
  assign t[354] = (x[86]);
  assign t[355] = (x[89]);
  assign t[356] = (x[89]);
  assign t[357] = (x[92]);
  assign t[358] = (x[92]);
  assign t[359] = (x[95]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[95]);
  assign t[361] = (x[98]);
  assign t[362] = (x[98]);
  assign t[363] = (x[101]);
  assign t[364] = (x[101]);
  assign t[365] = (x[104]);
  assign t[366] = (x[104]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[54] ^ t[41];
  assign t[370] = (x[110]);
  assign t[371] = (x[113]);
  assign t[372] = (x[113]);
  assign t[373] = (x[116]);
  assign t[374] = (x[116]);
  assign t[375] = (x[119]);
  assign t[376] = (x[119]);
  assign t[377] = (x[122]);
  assign t[378] = (x[122]);
  assign t[379] = (x[125]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[128]);
  assign t[382] = (x[128]);
  assign t[383] = (x[131]);
  assign t[384] = (x[131]);
  assign t[385] = (x[134]);
  assign t[386] = (x[134]);
  assign t[387] = (x[137]);
  assign t[388] = (x[137]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[18] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[67] | t[45]);
  assign t[48] = ~(t[68] & t[69]);
  assign t[49] = t[70] | t[111];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[105] ? x[40] : x[39];
  assign t[51] = ~(t[71] & t[72]);
  assign t[52] = ~(t[73] & t[74]);
  assign t[53] = t[75] | t[112];
  assign t[54] = t[76] ? x[45] : x[44];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = t[80] | t[115];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[116];
  assign t[62] = t[76] ? x[59] : x[58];
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = t[86] | t[117];
  assign t[65] = t[76] ? x[64] : x[63];
  assign t[66] = ~(t[87] & t[88]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = t[92] | t[121];
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[93] | t[73]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [151:0] x;
 output y;

 wire [520:0] t;
  assign t[0] = t[1] ? t[2] : t[206];
  assign t[100] = ~(t[228] | t[142]);
  assign t[101] = t[30] ? x[79] : x[78];
  assign t[102] = ~(t[143] & t[144]);
  assign t[103] = ~(t[229]);
  assign t[104] = ~(t[230]);
  assign t[105] = ~(t[145] | t[146]);
  assign t[106] = t[30] ? x[87] : x[86];
  assign t[107] = ~(t[147] & t[148]);
  assign t[108] = ~(t[231]);
  assign t[109] = ~(t[218] | t[219]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[232]);
  assign t[111] = ~(t[233]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[151] | t[152]);
  assign t[114] = ~(t[234]);
  assign t[115] = ~(t[235]);
  assign t[116] = ~(t[153] | t[154]);
  assign t[117] = t[155] ? x[104] : x[103];
  assign t[118] = t[156] | t[84];
  assign t[119] = ~(t[236]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[237]);
  assign t[121] = ~(t[157] | t[158]);
  assign t[122] = ~(t[159] | t[160]);
  assign t[123] = ~(t[238] | t[161]);
  assign t[124] = t[155] ? x[115] : x[114];
  assign t[125] = ~(t[162] & t[163]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(t[208] | t[166]);
  assign t[128] = t[129] & t[207];
  assign t[129] = ~(t[132]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[207] ? t[164] : t[167];
  assign t[131] = t[207] ? t[169] : t[168];
  assign t[132] = ~(t[209]);
  assign t[133] = ~(t[239]);
  assign t[134] = ~(t[224] | t[225]);
  assign t[135] = ~(t[132] | t[170]);
  assign t[136] = ~(t[129] | t[171]);
  assign t[137] = ~(t[172] & t[173]);
  assign t[138] = ~(t[240]);
  assign t[139] = ~(t[226] | t[227]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[241]);
  assign t[141] = ~(t[242]);
  assign t[142] = ~(t[174] | t[175]);
  assign t[143] = ~(t[151] | t[176]);
  assign t[144] = ~(t[118] | t[177]);
  assign t[145] = ~(t[243]);
  assign t[146] = ~(t[229] | t[230]);
  assign t[147] = ~(t[178] | t[85]);
  assign t[148] = ~(t[135] | t[156]);
  assign t[149] = ~(t[244]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[232] | t[233]);
  assign t[151] = ~(t[129] | t[179]);
  assign t[152] = ~(t[94] & t[180]);
  assign t[153] = ~(t[245]);
  assign t[154] = ~(t[234] | t[235]);
  assign t[155] = ~(t[49]);
  assign t[156] = ~(t[181] & t[83]);
  assign t[157] = ~(t[246]);
  assign t[158] = ~(t[236] | t[237]);
  assign t[159] = ~(t[247]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[248]);
  assign t[161] = ~(t[182] | t[183]);
  assign t[162] = ~(t[151]);
  assign t[163] = ~(t[184] | t[84]);
  assign t[164] = ~(t[210] & t[185]);
  assign t[165] = ~(x[4] & t[127]);
  assign t[166] = ~(t[210]);
  assign t[167] = ~(x[4] & t[186]);
  assign t[168] = ~(t[88] & t[166]);
  assign t[169] = ~(t[87] & t[210]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = t[207] ? t[187] : t[168];
  assign t[171] = t[207] ? t[188] : t[165];
  assign t[172] = ~(t[151] | t[189]);
  assign t[173] = t[132] | t[190];
  assign t[174] = ~(t[249]);
  assign t[175] = ~(t[241] | t[242]);
  assign t[176] = ~(t[129] | t[191]);
  assign t[177] = ~(t[192] & t[173]);
  assign t[178] = ~(t[129] | t[193]);
  assign t[179] = t[207] ? t[194] : t[187];
  assign t[17] = ~(t[209] & t[210]);
  assign t[180] = ~(t[132] & t[195]);
  assign t[181] = ~(t[196] | t[197]);
  assign t[182] = ~(t[250]);
  assign t[183] = ~(t[247] | t[248]);
  assign t[184] = ~(t[198]);
  assign t[185] = ~(x[4] | t[199]);
  assign t[186] = ~(t[208] | t[210]);
  assign t[187] = ~(t[87] & t[166]);
  assign t[188] = ~(t[185] & t[166]);
  assign t[189] = ~(t[129] | t[200]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[207] ? t[167] : t[188];
  assign t[191] = t[207] ? t[167] : t[164];
  assign t[192] = ~(t[201] | t[202]);
  assign t[193] = t[207] ? t[187] : t[194];
  assign t[194] = ~(t[88] & t[210]);
  assign t[195] = ~(t[167] & t[164]);
  assign t[196] = ~(t[132] | t[203]);
  assign t[197] = ~(t[132] | t[204]);
  assign t[198] = ~(t[202] | t[189]);
  assign t[199] = ~(t[208]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[207] ? t[168] : t[169];
  assign t[201] = ~(t[82]);
  assign t[202] = ~(t[129] | t[205]);
  assign t[203] = t[207] ? t[168] : t[187];
  assign t[204] = t[207] ? t[188] : t[167];
  assign t[205] = t[207] ? t[165] : t[188];
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = t[296] ^ x[2];
  assign t[252] = t[297] ^ x[10];
  assign t[253] = t[298] ^ x[13];
  assign t[254] = t[299] ^ x[16];
  assign t[255] = t[300] ^ x[19];
  assign t[256] = t[301] ^ x[22];
  assign t[257] = t[302] ^ x[25];
  assign t[258] = t[303] ^ x[28];
  assign t[259] = t[304] ^ x[31];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[34];
  assign t[261] = t[306] ^ x[39];
  assign t[262] = t[307] ^ x[42];
  assign t[263] = t[308] ^ x[45];
  assign t[264] = t[309] ^ x[48];
  assign t[265] = t[310] ^ x[51];
  assign t[266] = t[311] ^ x[56];
  assign t[267] = t[312] ^ x[59];
  assign t[268] = t[313] ^ x[62];
  assign t[269] = t[314] ^ x[65];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[68];
  assign t[271] = t[316] ^ x[71];
  assign t[272] = t[317] ^ x[74];
  assign t[273] = t[318] ^ x[77];
  assign t[274] = t[319] ^ x[82];
  assign t[275] = t[320] ^ x[85];
  assign t[276] = t[321] ^ x[90];
  assign t[277] = t[322] ^ x[93];
  assign t[278] = t[323] ^ x[96];
  assign t[279] = t[324] ^ x[99];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[102];
  assign t[281] = t[326] ^ x[107];
  assign t[282] = t[327] ^ x[110];
  assign t[283] = t[328] ^ x[113];
  assign t[284] = t[329] ^ x[118];
  assign t[285] = t[330] ^ x[121];
  assign t[286] = t[331] ^ x[124];
  assign t[287] = t[332] ^ x[127];
  assign t[288] = t[333] ^ x[130];
  assign t[289] = t[334] ^ x[133];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[136];
  assign t[291] = t[336] ^ x[139];
  assign t[292] = t[337] ^ x[142];
  assign t[293] = t[338] ^ x[145];
  assign t[294] = t[339] ^ x[148];
  assign t[295] = t[340] ^ x[151];
  assign t[296] = (t[341] & ~t[342]);
  assign t[297] = (t[343] & ~t[344]);
  assign t[298] = (t[345] & ~t[346]);
  assign t[299] = (t[347] & ~t[348]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[349] & ~t[350]);
  assign t[301] = (t[351] & ~t[352]);
  assign t[302] = (t[353] & ~t[354]);
  assign t[303] = (t[355] & ~t[356]);
  assign t[304] = (t[357] & ~t[358]);
  assign t[305] = (t[359] & ~t[360]);
  assign t[306] = (t[361] & ~t[362]);
  assign t[307] = (t[363] & ~t[364]);
  assign t[308] = (t[365] & ~t[366]);
  assign t[309] = (t[367] & ~t[368]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[369] & ~t[370]);
  assign t[311] = (t[371] & ~t[372]);
  assign t[312] = (t[373] & ~t[374]);
  assign t[313] = (t[375] & ~t[376]);
  assign t[314] = (t[377] & ~t[378]);
  assign t[315] = (t[379] & ~t[380]);
  assign t[316] = (t[381] & ~t[382]);
  assign t[317] = (t[383] & ~t[384]);
  assign t[318] = (t[385] & ~t[386]);
  assign t[319] = (t[387] & ~t[388]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[389] & ~t[390]);
  assign t[321] = (t[391] & ~t[392]);
  assign t[322] = (t[393] & ~t[394]);
  assign t[323] = (t[395] & ~t[396]);
  assign t[324] = (t[397] & ~t[398]);
  assign t[325] = (t[399] & ~t[400]);
  assign t[326] = (t[401] & ~t[402]);
  assign t[327] = (t[403] & ~t[404]);
  assign t[328] = (t[405] & ~t[406]);
  assign t[329] = (t[407] & ~t[408]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (t[409] & ~t[410]);
  assign t[331] = (t[411] & ~t[412]);
  assign t[332] = (t[413] & ~t[414]);
  assign t[333] = (t[415] & ~t[416]);
  assign t[334] = (t[417] & ~t[418]);
  assign t[335] = (t[419] & ~t[420]);
  assign t[336] = (t[421] & ~t[422]);
  assign t[337] = (t[423] & ~t[424]);
  assign t[338] = (t[425] & ~t[426]);
  assign t[339] = (t[427] & ~t[428]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (t[429] & ~t[430]);
  assign t[341] = t[431] ^ x[2];
  assign t[342] = t[432] ^ x[1];
  assign t[343] = t[433] ^ x[10];
  assign t[344] = t[434] ^ x[9];
  assign t[345] = t[435] ^ x[13];
  assign t[346] = t[436] ^ x[12];
  assign t[347] = t[437] ^ x[16];
  assign t[348] = t[438] ^ x[15];
  assign t[349] = t[439] ^ x[19];
  assign t[34] = ~(t[211] | t[56]);
  assign t[350] = t[440] ^ x[18];
  assign t[351] = t[441] ^ x[22];
  assign t[352] = t[442] ^ x[21];
  assign t[353] = t[443] ^ x[25];
  assign t[354] = t[444] ^ x[24];
  assign t[355] = t[445] ^ x[28];
  assign t[356] = t[446] ^ x[27];
  assign t[357] = t[447] ^ x[31];
  assign t[358] = t[448] ^ x[30];
  assign t[359] = t[449] ^ x[34];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[33];
  assign t[361] = t[451] ^ x[39];
  assign t[362] = t[452] ^ x[38];
  assign t[363] = t[453] ^ x[42];
  assign t[364] = t[454] ^ x[41];
  assign t[365] = t[455] ^ x[45];
  assign t[366] = t[456] ^ x[44];
  assign t[367] = t[457] ^ x[48];
  assign t[368] = t[458] ^ x[47];
  assign t[369] = t[459] ^ x[51];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[50];
  assign t[371] = t[461] ^ x[56];
  assign t[372] = t[462] ^ x[55];
  assign t[373] = t[463] ^ x[59];
  assign t[374] = t[464] ^ x[58];
  assign t[375] = t[465] ^ x[62];
  assign t[376] = t[466] ^ x[61];
  assign t[377] = t[467] ^ x[65];
  assign t[378] = t[468] ^ x[64];
  assign t[379] = t[469] ^ x[68];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[67];
  assign t[381] = t[471] ^ x[71];
  assign t[382] = t[472] ^ x[70];
  assign t[383] = t[473] ^ x[74];
  assign t[384] = t[474] ^ x[73];
  assign t[385] = t[475] ^ x[77];
  assign t[386] = t[476] ^ x[76];
  assign t[387] = t[477] ^ x[82];
  assign t[388] = t[478] ^ x[81];
  assign t[389] = t[479] ^ x[85];
  assign t[38] = ~(t[63] ^ t[64]);
  assign t[390] = t[480] ^ x[84];
  assign t[391] = t[481] ^ x[90];
  assign t[392] = t[482] ^ x[89];
  assign t[393] = t[483] ^ x[93];
  assign t[394] = t[484] ^ x[92];
  assign t[395] = t[485] ^ x[96];
  assign t[396] = t[486] ^ x[95];
  assign t[397] = t[487] ^ x[99];
  assign t[398] = t[488] ^ x[98];
  assign t[399] = t[489] ^ x[102];
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[101];
  assign t[401] = t[491] ^ x[107];
  assign t[402] = t[492] ^ x[106];
  assign t[403] = t[493] ^ x[110];
  assign t[404] = t[494] ^ x[109];
  assign t[405] = t[495] ^ x[113];
  assign t[406] = t[496] ^ x[112];
  assign t[407] = t[497] ^ x[118];
  assign t[408] = t[498] ^ x[117];
  assign t[409] = t[499] ^ x[121];
  assign t[40] = ~(t[37] ^ t[67]);
  assign t[410] = t[500] ^ x[120];
  assign t[411] = t[501] ^ x[124];
  assign t[412] = t[502] ^ x[123];
  assign t[413] = t[503] ^ x[127];
  assign t[414] = t[504] ^ x[126];
  assign t[415] = t[505] ^ x[130];
  assign t[416] = t[506] ^ x[129];
  assign t[417] = t[507] ^ x[133];
  assign t[418] = t[508] ^ x[132];
  assign t[419] = t[509] ^ x[136];
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = t[510] ^ x[135];
  assign t[421] = t[511] ^ x[139];
  assign t[422] = t[512] ^ x[138];
  assign t[423] = t[513] ^ x[142];
  assign t[424] = t[514] ^ x[141];
  assign t[425] = t[515] ^ x[145];
  assign t[426] = t[516] ^ x[144];
  assign t[427] = t[517] ^ x[148];
  assign t[428] = t[518] ^ x[147];
  assign t[429] = t[519] ^ x[151];
  assign t[42] = ~(t[212] | t[70]);
  assign t[430] = t[520] ^ x[150];
  assign t[431] = (x[0]);
  assign t[432] = (x[0]);
  assign t[433] = (x[8]);
  assign t[434] = (x[8]);
  assign t[435] = (x[11]);
  assign t[436] = (x[11]);
  assign t[437] = (x[14]);
  assign t[438] = (x[14]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[17]);
  assign t[441] = (x[20]);
  assign t[442] = (x[20]);
  assign t[443] = (x[23]);
  assign t[444] = (x[23]);
  assign t[445] = (x[26]);
  assign t[446] = (x[26]);
  assign t[447] = (x[29]);
  assign t[448] = (x[29]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[32]);
  assign t[451] = (x[37]);
  assign t[452] = (x[37]);
  assign t[453] = (x[40]);
  assign t[454] = (x[40]);
  assign t[455] = (x[43]);
  assign t[456] = (x[43]);
  assign t[457] = (x[46]);
  assign t[458] = (x[46]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = (x[49]);
  assign t[461] = (x[54]);
  assign t[462] = (x[54]);
  assign t[463] = (x[57]);
  assign t[464] = (x[57]);
  assign t[465] = (x[60]);
  assign t[466] = (x[60]);
  assign t[467] = (x[63]);
  assign t[468] = (x[63]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[47] ^ t[77]);
  assign t[470] = (x[66]);
  assign t[471] = (x[69]);
  assign t[472] = (x[69]);
  assign t[473] = (x[72]);
  assign t[474] = (x[72]);
  assign t[475] = (x[75]);
  assign t[476] = (x[75]);
  assign t[477] = (x[80]);
  assign t[478] = (x[80]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = (x[83]);
  assign t[481] = (x[88]);
  assign t[482] = (x[88]);
  assign t[483] = (x[91]);
  assign t[484] = (x[91]);
  assign t[485] = (x[94]);
  assign t[486] = (x[94]);
  assign t[487] = (x[97]);
  assign t[488] = (x[97]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = (x[100]);
  assign t[491] = (x[105]);
  assign t[492] = (x[105]);
  assign t[493] = (x[108]);
  assign t[494] = (x[108]);
  assign t[495] = (x[111]);
  assign t[496] = (x[111]);
  assign t[497] = (x[116]);
  assign t[498] = (x[116]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[209]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[119]);
  assign t[501] = (x[122]);
  assign t[502] = (x[122]);
  assign t[503] = (x[125]);
  assign t[504] = (x[125]);
  assign t[505] = (x[128]);
  assign t[506] = (x[128]);
  assign t[507] = (x[131]);
  assign t[508] = (x[131]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (x[134]);
  assign t[511] = (x[137]);
  assign t[512] = (x[137]);
  assign t[513] = (x[140]);
  assign t[514] = (x[140]);
  assign t[515] = (x[143]);
  assign t[516] = (x[143]);
  assign t[517] = (x[146]);
  assign t[518] = (x[146]);
  assign t[519] = (x[149]);
  assign t[51] = t[84] | t[85];
  assign t[520] = (x[149]);
  assign t[52] = t[210] & t[86];
  assign t[53] = t[87] | t[88];
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[214]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[215] | t[93]);
  assign t[59] = t[30] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[216] | t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[66] = ~(t[217] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[218]);
  assign t[69] = ~(t[219]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[220] | t[112]);
  assign t[73] = t[30] ? x[53] : x[52];
  assign t[74] = ~(t[113] & t[83]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[221] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119] | t[120]);
  assign t[79] = ~(t[222] | t[121]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[122] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[86] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = ~(t[129] | t[130]);
  assign t[85] = ~(t[129] | t[131]);
  assign t[86] = ~(t[132] | t[207]);
  assign t[87] = ~(x[4] | t[208]);
  assign t[88] = x[4] & t[208];
  assign t[89] = ~(t[223]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[213] | t[214]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[225]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[135] | t[136]);
  assign t[95] = ~(t[85] | t[137]);
  assign t[96] = ~(t[226]);
  assign t[97] = ~(t[227]);
  assign t[98] = ~(t[138] | t[139]);
  assign t[99] = ~(t[140] | t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [151:0] x;
 output y;

 wire [520:0] t;
  assign t[0] = t[1] ? t[2] : t[206];
  assign t[100] = ~(t[228] | t[142]);
  assign t[101] = t[30] ? x[79] : x[78];
  assign t[102] = ~(t[143] & t[144]);
  assign t[103] = ~(t[229]);
  assign t[104] = ~(t[230]);
  assign t[105] = ~(t[145] | t[146]);
  assign t[106] = t[30] ? x[87] : x[86];
  assign t[107] = ~(t[147] & t[148]);
  assign t[108] = ~(t[231]);
  assign t[109] = ~(t[218] | t[219]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[232]);
  assign t[111] = ~(t[233]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[151] | t[152]);
  assign t[114] = ~(t[234]);
  assign t[115] = ~(t[235]);
  assign t[116] = ~(t[153] | t[154]);
  assign t[117] = t[155] ? x[104] : x[103];
  assign t[118] = t[156] | t[84];
  assign t[119] = ~(t[236]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[237]);
  assign t[121] = ~(t[157] | t[158]);
  assign t[122] = ~(t[159] | t[160]);
  assign t[123] = ~(t[238] | t[161]);
  assign t[124] = t[155] ? x[115] : x[114];
  assign t[125] = ~(t[162] & t[163]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(t[208] | t[166]);
  assign t[128] = t[129] & t[207];
  assign t[129] = ~(t[132]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[207] ? t[164] : t[167];
  assign t[131] = t[207] ? t[169] : t[168];
  assign t[132] = ~(t[209]);
  assign t[133] = ~(t[239]);
  assign t[134] = ~(t[224] | t[225]);
  assign t[135] = ~(t[132] | t[170]);
  assign t[136] = ~(t[129] | t[171]);
  assign t[137] = ~(t[172] & t[173]);
  assign t[138] = ~(t[240]);
  assign t[139] = ~(t[226] | t[227]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[241]);
  assign t[141] = ~(t[242]);
  assign t[142] = ~(t[174] | t[175]);
  assign t[143] = ~(t[151] | t[176]);
  assign t[144] = ~(t[118] | t[177]);
  assign t[145] = ~(t[243]);
  assign t[146] = ~(t[229] | t[230]);
  assign t[147] = ~(t[178] | t[85]);
  assign t[148] = ~(t[135] | t[156]);
  assign t[149] = ~(t[244]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[232] | t[233]);
  assign t[151] = ~(t[129] | t[179]);
  assign t[152] = ~(t[94] & t[180]);
  assign t[153] = ~(t[245]);
  assign t[154] = ~(t[234] | t[235]);
  assign t[155] = ~(t[49]);
  assign t[156] = ~(t[181] & t[83]);
  assign t[157] = ~(t[246]);
  assign t[158] = ~(t[236] | t[237]);
  assign t[159] = ~(t[247]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[248]);
  assign t[161] = ~(t[182] | t[183]);
  assign t[162] = ~(t[151]);
  assign t[163] = ~(t[184] | t[84]);
  assign t[164] = ~(t[210] & t[185]);
  assign t[165] = ~(x[4] & t[127]);
  assign t[166] = ~(t[210]);
  assign t[167] = ~(x[4] & t[186]);
  assign t[168] = ~(t[88] & t[166]);
  assign t[169] = ~(t[87] & t[210]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = t[207] ? t[187] : t[168];
  assign t[171] = t[207] ? t[188] : t[165];
  assign t[172] = ~(t[151] | t[189]);
  assign t[173] = t[132] | t[190];
  assign t[174] = ~(t[249]);
  assign t[175] = ~(t[241] | t[242]);
  assign t[176] = ~(t[129] | t[191]);
  assign t[177] = ~(t[192] & t[173]);
  assign t[178] = ~(t[129] | t[193]);
  assign t[179] = t[207] ? t[194] : t[187];
  assign t[17] = ~(t[209] & t[210]);
  assign t[180] = ~(t[132] & t[195]);
  assign t[181] = ~(t[196] | t[197]);
  assign t[182] = ~(t[250]);
  assign t[183] = ~(t[247] | t[248]);
  assign t[184] = ~(t[198]);
  assign t[185] = ~(x[4] | t[199]);
  assign t[186] = ~(t[208] | t[210]);
  assign t[187] = ~(t[87] & t[166]);
  assign t[188] = ~(t[185] & t[166]);
  assign t[189] = ~(t[129] | t[200]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[207] ? t[167] : t[188];
  assign t[191] = t[207] ? t[167] : t[164];
  assign t[192] = ~(t[201] | t[202]);
  assign t[193] = t[207] ? t[187] : t[194];
  assign t[194] = ~(t[88] & t[210]);
  assign t[195] = ~(t[167] & t[164]);
  assign t[196] = ~(t[132] | t[203]);
  assign t[197] = ~(t[132] | t[204]);
  assign t[198] = ~(t[202] | t[189]);
  assign t[199] = ~(t[208]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[207] ? t[168] : t[169];
  assign t[201] = ~(t[82]);
  assign t[202] = ~(t[129] | t[205]);
  assign t[203] = t[207] ? t[168] : t[187];
  assign t[204] = t[207] ? t[188] : t[167];
  assign t[205] = t[207] ? t[165] : t[188];
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = t[296] ^ x[2];
  assign t[252] = t[297] ^ x[10];
  assign t[253] = t[298] ^ x[13];
  assign t[254] = t[299] ^ x[16];
  assign t[255] = t[300] ^ x[19];
  assign t[256] = t[301] ^ x[22];
  assign t[257] = t[302] ^ x[25];
  assign t[258] = t[303] ^ x[28];
  assign t[259] = t[304] ^ x[31];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[34];
  assign t[261] = t[306] ^ x[39];
  assign t[262] = t[307] ^ x[42];
  assign t[263] = t[308] ^ x[45];
  assign t[264] = t[309] ^ x[48];
  assign t[265] = t[310] ^ x[51];
  assign t[266] = t[311] ^ x[56];
  assign t[267] = t[312] ^ x[59];
  assign t[268] = t[313] ^ x[62];
  assign t[269] = t[314] ^ x[65];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[68];
  assign t[271] = t[316] ^ x[71];
  assign t[272] = t[317] ^ x[74];
  assign t[273] = t[318] ^ x[77];
  assign t[274] = t[319] ^ x[82];
  assign t[275] = t[320] ^ x[85];
  assign t[276] = t[321] ^ x[90];
  assign t[277] = t[322] ^ x[93];
  assign t[278] = t[323] ^ x[96];
  assign t[279] = t[324] ^ x[99];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[102];
  assign t[281] = t[326] ^ x[107];
  assign t[282] = t[327] ^ x[110];
  assign t[283] = t[328] ^ x[113];
  assign t[284] = t[329] ^ x[118];
  assign t[285] = t[330] ^ x[121];
  assign t[286] = t[331] ^ x[124];
  assign t[287] = t[332] ^ x[127];
  assign t[288] = t[333] ^ x[130];
  assign t[289] = t[334] ^ x[133];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[136];
  assign t[291] = t[336] ^ x[139];
  assign t[292] = t[337] ^ x[142];
  assign t[293] = t[338] ^ x[145];
  assign t[294] = t[339] ^ x[148];
  assign t[295] = t[340] ^ x[151];
  assign t[296] = (t[341] & ~t[342]);
  assign t[297] = (t[343] & ~t[344]);
  assign t[298] = (t[345] & ~t[346]);
  assign t[299] = (t[347] & ~t[348]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[349] & ~t[350]);
  assign t[301] = (t[351] & ~t[352]);
  assign t[302] = (t[353] & ~t[354]);
  assign t[303] = (t[355] & ~t[356]);
  assign t[304] = (t[357] & ~t[358]);
  assign t[305] = (t[359] & ~t[360]);
  assign t[306] = (t[361] & ~t[362]);
  assign t[307] = (t[363] & ~t[364]);
  assign t[308] = (t[365] & ~t[366]);
  assign t[309] = (t[367] & ~t[368]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[369] & ~t[370]);
  assign t[311] = (t[371] & ~t[372]);
  assign t[312] = (t[373] & ~t[374]);
  assign t[313] = (t[375] & ~t[376]);
  assign t[314] = (t[377] & ~t[378]);
  assign t[315] = (t[379] & ~t[380]);
  assign t[316] = (t[381] & ~t[382]);
  assign t[317] = (t[383] & ~t[384]);
  assign t[318] = (t[385] & ~t[386]);
  assign t[319] = (t[387] & ~t[388]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[389] & ~t[390]);
  assign t[321] = (t[391] & ~t[392]);
  assign t[322] = (t[393] & ~t[394]);
  assign t[323] = (t[395] & ~t[396]);
  assign t[324] = (t[397] & ~t[398]);
  assign t[325] = (t[399] & ~t[400]);
  assign t[326] = (t[401] & ~t[402]);
  assign t[327] = (t[403] & ~t[404]);
  assign t[328] = (t[405] & ~t[406]);
  assign t[329] = (t[407] & ~t[408]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (t[409] & ~t[410]);
  assign t[331] = (t[411] & ~t[412]);
  assign t[332] = (t[413] & ~t[414]);
  assign t[333] = (t[415] & ~t[416]);
  assign t[334] = (t[417] & ~t[418]);
  assign t[335] = (t[419] & ~t[420]);
  assign t[336] = (t[421] & ~t[422]);
  assign t[337] = (t[423] & ~t[424]);
  assign t[338] = (t[425] & ~t[426]);
  assign t[339] = (t[427] & ~t[428]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (t[429] & ~t[430]);
  assign t[341] = t[431] ^ x[2];
  assign t[342] = t[432] ^ x[1];
  assign t[343] = t[433] ^ x[10];
  assign t[344] = t[434] ^ x[9];
  assign t[345] = t[435] ^ x[13];
  assign t[346] = t[436] ^ x[12];
  assign t[347] = t[437] ^ x[16];
  assign t[348] = t[438] ^ x[15];
  assign t[349] = t[439] ^ x[19];
  assign t[34] = ~(t[211] | t[56]);
  assign t[350] = t[440] ^ x[18];
  assign t[351] = t[441] ^ x[22];
  assign t[352] = t[442] ^ x[21];
  assign t[353] = t[443] ^ x[25];
  assign t[354] = t[444] ^ x[24];
  assign t[355] = t[445] ^ x[28];
  assign t[356] = t[446] ^ x[27];
  assign t[357] = t[447] ^ x[31];
  assign t[358] = t[448] ^ x[30];
  assign t[359] = t[449] ^ x[34];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[450] ^ x[33];
  assign t[361] = t[451] ^ x[39];
  assign t[362] = t[452] ^ x[38];
  assign t[363] = t[453] ^ x[42];
  assign t[364] = t[454] ^ x[41];
  assign t[365] = t[455] ^ x[45];
  assign t[366] = t[456] ^ x[44];
  assign t[367] = t[457] ^ x[48];
  assign t[368] = t[458] ^ x[47];
  assign t[369] = t[459] ^ x[51];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[460] ^ x[50];
  assign t[371] = t[461] ^ x[56];
  assign t[372] = t[462] ^ x[55];
  assign t[373] = t[463] ^ x[59];
  assign t[374] = t[464] ^ x[58];
  assign t[375] = t[465] ^ x[62];
  assign t[376] = t[466] ^ x[61];
  assign t[377] = t[467] ^ x[65];
  assign t[378] = t[468] ^ x[64];
  assign t[379] = t[469] ^ x[68];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[470] ^ x[67];
  assign t[381] = t[471] ^ x[71];
  assign t[382] = t[472] ^ x[70];
  assign t[383] = t[473] ^ x[74];
  assign t[384] = t[474] ^ x[73];
  assign t[385] = t[475] ^ x[77];
  assign t[386] = t[476] ^ x[76];
  assign t[387] = t[477] ^ x[82];
  assign t[388] = t[478] ^ x[81];
  assign t[389] = t[479] ^ x[85];
  assign t[38] = ~(t[63] ^ t[64]);
  assign t[390] = t[480] ^ x[84];
  assign t[391] = t[481] ^ x[90];
  assign t[392] = t[482] ^ x[89];
  assign t[393] = t[483] ^ x[93];
  assign t[394] = t[484] ^ x[92];
  assign t[395] = t[485] ^ x[96];
  assign t[396] = t[486] ^ x[95];
  assign t[397] = t[487] ^ x[99];
  assign t[398] = t[488] ^ x[98];
  assign t[399] = t[489] ^ x[102];
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[101];
  assign t[401] = t[491] ^ x[107];
  assign t[402] = t[492] ^ x[106];
  assign t[403] = t[493] ^ x[110];
  assign t[404] = t[494] ^ x[109];
  assign t[405] = t[495] ^ x[113];
  assign t[406] = t[496] ^ x[112];
  assign t[407] = t[497] ^ x[118];
  assign t[408] = t[498] ^ x[117];
  assign t[409] = t[499] ^ x[121];
  assign t[40] = ~(t[37] ^ t[67]);
  assign t[410] = t[500] ^ x[120];
  assign t[411] = t[501] ^ x[124];
  assign t[412] = t[502] ^ x[123];
  assign t[413] = t[503] ^ x[127];
  assign t[414] = t[504] ^ x[126];
  assign t[415] = t[505] ^ x[130];
  assign t[416] = t[506] ^ x[129];
  assign t[417] = t[507] ^ x[133];
  assign t[418] = t[508] ^ x[132];
  assign t[419] = t[509] ^ x[136];
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = t[510] ^ x[135];
  assign t[421] = t[511] ^ x[139];
  assign t[422] = t[512] ^ x[138];
  assign t[423] = t[513] ^ x[142];
  assign t[424] = t[514] ^ x[141];
  assign t[425] = t[515] ^ x[145];
  assign t[426] = t[516] ^ x[144];
  assign t[427] = t[517] ^ x[148];
  assign t[428] = t[518] ^ x[147];
  assign t[429] = t[519] ^ x[151];
  assign t[42] = ~(t[212] | t[70]);
  assign t[430] = t[520] ^ x[150];
  assign t[431] = (x[0]);
  assign t[432] = (x[0]);
  assign t[433] = (x[8]);
  assign t[434] = (x[8]);
  assign t[435] = (x[11]);
  assign t[436] = (x[11]);
  assign t[437] = (x[14]);
  assign t[438] = (x[14]);
  assign t[439] = (x[17]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[17]);
  assign t[441] = (x[20]);
  assign t[442] = (x[20]);
  assign t[443] = (x[23]);
  assign t[444] = (x[23]);
  assign t[445] = (x[26]);
  assign t[446] = (x[26]);
  assign t[447] = (x[29]);
  assign t[448] = (x[29]);
  assign t[449] = (x[32]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[32]);
  assign t[451] = (x[37]);
  assign t[452] = (x[37]);
  assign t[453] = (x[40]);
  assign t[454] = (x[40]);
  assign t[455] = (x[43]);
  assign t[456] = (x[43]);
  assign t[457] = (x[46]);
  assign t[458] = (x[46]);
  assign t[459] = (x[49]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = (x[49]);
  assign t[461] = (x[54]);
  assign t[462] = (x[54]);
  assign t[463] = (x[57]);
  assign t[464] = (x[57]);
  assign t[465] = (x[60]);
  assign t[466] = (x[60]);
  assign t[467] = (x[63]);
  assign t[468] = (x[63]);
  assign t[469] = (x[66]);
  assign t[46] = ~(t[47] ^ t[77]);
  assign t[470] = (x[66]);
  assign t[471] = (x[69]);
  assign t[472] = (x[69]);
  assign t[473] = (x[72]);
  assign t[474] = (x[72]);
  assign t[475] = (x[75]);
  assign t[476] = (x[75]);
  assign t[477] = (x[80]);
  assign t[478] = (x[80]);
  assign t[479] = (x[83]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = (x[83]);
  assign t[481] = (x[88]);
  assign t[482] = (x[88]);
  assign t[483] = (x[91]);
  assign t[484] = (x[91]);
  assign t[485] = (x[94]);
  assign t[486] = (x[94]);
  assign t[487] = (x[97]);
  assign t[488] = (x[97]);
  assign t[489] = (x[100]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = (x[100]);
  assign t[491] = (x[105]);
  assign t[492] = (x[105]);
  assign t[493] = (x[108]);
  assign t[494] = (x[108]);
  assign t[495] = (x[111]);
  assign t[496] = (x[111]);
  assign t[497] = (x[116]);
  assign t[498] = (x[116]);
  assign t[499] = (x[119]);
  assign t[49] = ~(t[209]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[119]);
  assign t[501] = (x[122]);
  assign t[502] = (x[122]);
  assign t[503] = (x[125]);
  assign t[504] = (x[125]);
  assign t[505] = (x[128]);
  assign t[506] = (x[128]);
  assign t[507] = (x[131]);
  assign t[508] = (x[131]);
  assign t[509] = (x[134]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (x[134]);
  assign t[511] = (x[137]);
  assign t[512] = (x[137]);
  assign t[513] = (x[140]);
  assign t[514] = (x[140]);
  assign t[515] = (x[143]);
  assign t[516] = (x[143]);
  assign t[517] = (x[146]);
  assign t[518] = (x[146]);
  assign t[519] = (x[149]);
  assign t[51] = t[84] | t[85];
  assign t[520] = (x[149]);
  assign t[52] = t[210] & t[86];
  assign t[53] = t[87] | t[88];
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[214]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[215] | t[93]);
  assign t[59] = t[30] ? x[36] : x[35];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[216] | t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[66] = ~(t[217] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[218]);
  assign t[69] = ~(t[219]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[220] | t[112]);
  assign t[73] = t[30] ? x[53] : x[52];
  assign t[74] = ~(t[113] & t[83]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[221] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119] | t[120]);
  assign t[79] = ~(t[222] | t[121]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[122] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[86] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = ~(t[129] | t[130]);
  assign t[85] = ~(t[129] | t[131]);
  assign t[86] = ~(t[132] | t[207]);
  assign t[87] = ~(x[4] | t[208]);
  assign t[88] = x[4] & t[208];
  assign t[89] = ~(t[223]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[213] | t[214]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[225]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[135] | t[136]);
  assign t[95] = ~(t[85] | t[137]);
  assign t[96] = ~(t[226]);
  assign t[97] = ~(t[227]);
  assign t[98] = ~(t[138] | t[139]);
  assign t[99] = ~(t[140] | t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [121:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[99];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = t[169] ^ x[2];
  assign t[135] = t[170] ^ x[10];
  assign t[136] = t[171] ^ x[13];
  assign t[137] = t[172] ^ x[16];
  assign t[138] = t[173] ^ x[19];
  assign t[139] = t[174] ^ x[22];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[25];
  assign t[141] = t[176] ^ x[30];
  assign t[142] = t[177] ^ x[33];
  assign t[143] = t[178] ^ x[38];
  assign t[144] = t[179] ^ x[41];
  assign t[145] = t[180] ^ x[44];
  assign t[146] = t[181] ^ x[47];
  assign t[147] = t[182] ^ x[50];
  assign t[148] = t[183] ^ x[55];
  assign t[149] = t[184] ^ x[58];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[63];
  assign t[151] = t[186] ^ x[66];
  assign t[152] = t[187] ^ x[69];
  assign t[153] = t[188] ^ x[72];
  assign t[154] = t[189] ^ x[75];
  assign t[155] = t[190] ^ x[80];
  assign t[156] = t[191] ^ x[83];
  assign t[157] = t[192] ^ x[88];
  assign t[158] = t[193] ^ x[91];
  assign t[159] = t[194] ^ x[94];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[97];
  assign t[161] = t[196] ^ x[100];
  assign t[162] = t[197] ^ x[103];
  assign t[163] = t[198] ^ x[106];
  assign t[164] = t[199] ^ x[109];
  assign t[165] = t[200] ^ x[112];
  assign t[166] = t[201] ^ x[115];
  assign t[167] = t[202] ^ x[118];
  assign t[168] = t[203] ^ x[121];
  assign t[169] = (t[204] & ~t[205]);
  assign t[16] = ~(t[100] & t[101]);
  assign t[170] = (t[206] & ~t[207]);
  assign t[171] = (t[208] & ~t[209]);
  assign t[172] = (t[210] & ~t[211]);
  assign t[173] = (t[212] & ~t[213]);
  assign t[174] = (t[214] & ~t[215]);
  assign t[175] = (t[216] & ~t[217]);
  assign t[176] = (t[218] & ~t[219]);
  assign t[177] = (t[220] & ~t[221]);
  assign t[178] = (t[222] & ~t[223]);
  assign t[179] = (t[224] & ~t[225]);
  assign t[17] = ~(t[102] & t[103]);
  assign t[180] = (t[226] & ~t[227]);
  assign t[181] = (t[228] & ~t[229]);
  assign t[182] = (t[230] & ~t[231]);
  assign t[183] = (t[232] & ~t[233]);
  assign t[184] = (t[234] & ~t[235]);
  assign t[185] = (t[236] & ~t[237]);
  assign t[186] = (t[238] & ~t[239]);
  assign t[187] = (t[240] & ~t[241]);
  assign t[188] = (t[242] & ~t[243]);
  assign t[189] = (t[244] & ~t[245]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[246] & ~t[247]);
  assign t[191] = (t[248] & ~t[249]);
  assign t[192] = (t[250] & ~t[251]);
  assign t[193] = (t[252] & ~t[253]);
  assign t[194] = (t[254] & ~t[255]);
  assign t[195] = (t[256] & ~t[257]);
  assign t[196] = (t[258] & ~t[259]);
  assign t[197] = (t[260] & ~t[261]);
  assign t[198] = (t[262] & ~t[263]);
  assign t[199] = (t[264] & ~t[265]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[266] & ~t[267]);
  assign t[201] = (t[268] & ~t[269]);
  assign t[202] = (t[270] & ~t[271]);
  assign t[203] = (t[272] & ~t[273]);
  assign t[204] = t[274] ^ x[2];
  assign t[205] = t[275] ^ x[1];
  assign t[206] = t[276] ^ x[10];
  assign t[207] = t[277] ^ x[9];
  assign t[208] = t[278] ^ x[13];
  assign t[209] = t[279] ^ x[12];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[16];
  assign t[211] = t[281] ^ x[15];
  assign t[212] = t[282] ^ x[19];
  assign t[213] = t[283] ^ x[18];
  assign t[214] = t[284] ^ x[22];
  assign t[215] = t[285] ^ x[21];
  assign t[216] = t[286] ^ x[25];
  assign t[217] = t[287] ^ x[24];
  assign t[218] = t[288] ^ x[30];
  assign t[219] = t[289] ^ x[29];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[33];
  assign t[221] = t[291] ^ x[32];
  assign t[222] = t[292] ^ x[38];
  assign t[223] = t[293] ^ x[37];
  assign t[224] = t[294] ^ x[41];
  assign t[225] = t[295] ^ x[40];
  assign t[226] = t[296] ^ x[44];
  assign t[227] = t[297] ^ x[43];
  assign t[228] = t[298] ^ x[47];
  assign t[229] = t[299] ^ x[46];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[50];
  assign t[231] = t[301] ^ x[49];
  assign t[232] = t[302] ^ x[55];
  assign t[233] = t[303] ^ x[54];
  assign t[234] = t[304] ^ x[58];
  assign t[235] = t[305] ^ x[57];
  assign t[236] = t[306] ^ x[63];
  assign t[237] = t[307] ^ x[62];
  assign t[238] = t[308] ^ x[66];
  assign t[239] = t[309] ^ x[65];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[69];
  assign t[241] = t[311] ^ x[68];
  assign t[242] = t[312] ^ x[72];
  assign t[243] = t[313] ^ x[71];
  assign t[244] = t[314] ^ x[75];
  assign t[245] = t[315] ^ x[74];
  assign t[246] = t[316] ^ x[80];
  assign t[247] = t[317] ^ x[79];
  assign t[248] = t[318] ^ x[83];
  assign t[249] = t[319] ^ x[82];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[88];
  assign t[251] = t[321] ^ x[87];
  assign t[252] = t[322] ^ x[91];
  assign t[253] = t[323] ^ x[90];
  assign t[254] = t[324] ^ x[94];
  assign t[255] = t[325] ^ x[93];
  assign t[256] = t[326] ^ x[97];
  assign t[257] = t[327] ^ x[96];
  assign t[258] = t[328] ^ x[100];
  assign t[259] = t[329] ^ x[99];
  assign t[25] = ~(t[102]);
  assign t[260] = t[330] ^ x[103];
  assign t[261] = t[331] ^ x[102];
  assign t[262] = t[332] ^ x[106];
  assign t[263] = t[333] ^ x[105];
  assign t[264] = t[334] ^ x[109];
  assign t[265] = t[335] ^ x[108];
  assign t[266] = t[336] ^ x[112];
  assign t[267] = t[337] ^ x[111];
  assign t[268] = t[338] ^ x[115];
  assign t[269] = t[339] ^ x[114];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[118];
  assign t[271] = t[341] ^ x[117];
  assign t[272] = t[342] ^ x[121];
  assign t[273] = t[343] ^ x[120];
  assign t[274] = (x[0]);
  assign t[275] = (x[0]);
  assign t[276] = (x[8]);
  assign t[277] = (x[8]);
  assign t[278] = (x[11]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[14]);
  assign t[281] = (x[14]);
  assign t[282] = (x[17]);
  assign t[283] = (x[17]);
  assign t[284] = (x[20]);
  assign t[285] = (x[20]);
  assign t[286] = (x[23]);
  assign t[287] = (x[23]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[36]);
  assign t[293] = (x[36]);
  assign t[294] = (x[39]);
  assign t[295] = (x[39]);
  assign t[296] = (x[42]);
  assign t[297] = (x[42]);
  assign t[298] = (x[45]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[53]);
  assign t[303] = (x[53]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[61]);
  assign t[307] = (x[61]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[104] & t[46]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[70]);
  assign t[313] = (x[70]);
  assign t[314] = (x[73]);
  assign t[315] = (x[73]);
  assign t[316] = (x[78]);
  assign t[317] = (x[78]);
  assign t[318] = (x[81]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[105] & t[47]);
  assign t[320] = (x[86]);
  assign t[321] = (x[86]);
  assign t[322] = (x[89]);
  assign t[323] = (x[89]);
  assign t[324] = (x[92]);
  assign t[325] = (x[92]);
  assign t[326] = (x[95]);
  assign t[327] = (x[95]);
  assign t[328] = (x[98]);
  assign t[329] = (x[98]);
  assign t[32] = t[18] ? x[27] : x[26];
  assign t[330] = (x[101]);
  assign t[331] = (x[101]);
  assign t[332] = (x[104]);
  assign t[333] = (x[104]);
  assign t[334] = (x[107]);
  assign t[335] = (x[107]);
  assign t[336] = (x[110]);
  assign t[337] = (x[110]);
  assign t[338] = (x[113]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[116]);
  assign t[341] = (x[116]);
  assign t[342] = (x[119]);
  assign t[343] = (x[119]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[36];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[56];
  assign t[38] = ~(t[106] & t[57]);
  assign t[39] = ~(t[107] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[35] : x[34];
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[42];
  assign t[46] = ~(t[108]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[73] ? x[52] : x[51];
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = t[18] ? x[60] : x[59];
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[73] ? x[77] : x[76];
  assign t[64] = ~(t[83] & t[84]);
  assign t[65] = ~(t[120] & t[85]);
  assign t[66] = ~(t[121] & t[86]);
  assign t[67] = t[73] ? x[85] : x[84];
  assign t[68] = ~(t[104]);
  assign t[69] = ~(t[122]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[25]);
  assign t[74] = ~(t[124]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[132]);
  assign t[91] = ~(t[132] & t[97]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[133]);
  assign t[95] = ~(t[133] & t[98]);
  assign t[96] = ~(t[120]);
  assign t[97] = ~(t[125]);
  assign t[98] = ~(t[129]);
  assign t[99] = (t[134]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [121:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[99];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = t[169] ^ x[2];
  assign t[135] = t[170] ^ x[10];
  assign t[136] = t[171] ^ x[13];
  assign t[137] = t[172] ^ x[16];
  assign t[138] = t[173] ^ x[19];
  assign t[139] = t[174] ^ x[22];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[25];
  assign t[141] = t[176] ^ x[30];
  assign t[142] = t[177] ^ x[33];
  assign t[143] = t[178] ^ x[38];
  assign t[144] = t[179] ^ x[41];
  assign t[145] = t[180] ^ x[44];
  assign t[146] = t[181] ^ x[47];
  assign t[147] = t[182] ^ x[50];
  assign t[148] = t[183] ^ x[55];
  assign t[149] = t[184] ^ x[58];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[63];
  assign t[151] = t[186] ^ x[66];
  assign t[152] = t[187] ^ x[69];
  assign t[153] = t[188] ^ x[72];
  assign t[154] = t[189] ^ x[75];
  assign t[155] = t[190] ^ x[80];
  assign t[156] = t[191] ^ x[83];
  assign t[157] = t[192] ^ x[88];
  assign t[158] = t[193] ^ x[91];
  assign t[159] = t[194] ^ x[94];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[97];
  assign t[161] = t[196] ^ x[100];
  assign t[162] = t[197] ^ x[103];
  assign t[163] = t[198] ^ x[106];
  assign t[164] = t[199] ^ x[109];
  assign t[165] = t[200] ^ x[112];
  assign t[166] = t[201] ^ x[115];
  assign t[167] = t[202] ^ x[118];
  assign t[168] = t[203] ^ x[121];
  assign t[169] = (t[204] & ~t[205]);
  assign t[16] = ~(t[100] & t[101]);
  assign t[170] = (t[206] & ~t[207]);
  assign t[171] = (t[208] & ~t[209]);
  assign t[172] = (t[210] & ~t[211]);
  assign t[173] = (t[212] & ~t[213]);
  assign t[174] = (t[214] & ~t[215]);
  assign t[175] = (t[216] & ~t[217]);
  assign t[176] = (t[218] & ~t[219]);
  assign t[177] = (t[220] & ~t[221]);
  assign t[178] = (t[222] & ~t[223]);
  assign t[179] = (t[224] & ~t[225]);
  assign t[17] = ~(t[102] & t[103]);
  assign t[180] = (t[226] & ~t[227]);
  assign t[181] = (t[228] & ~t[229]);
  assign t[182] = (t[230] & ~t[231]);
  assign t[183] = (t[232] & ~t[233]);
  assign t[184] = (t[234] & ~t[235]);
  assign t[185] = (t[236] & ~t[237]);
  assign t[186] = (t[238] & ~t[239]);
  assign t[187] = (t[240] & ~t[241]);
  assign t[188] = (t[242] & ~t[243]);
  assign t[189] = (t[244] & ~t[245]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[246] & ~t[247]);
  assign t[191] = (t[248] & ~t[249]);
  assign t[192] = (t[250] & ~t[251]);
  assign t[193] = (t[252] & ~t[253]);
  assign t[194] = (t[254] & ~t[255]);
  assign t[195] = (t[256] & ~t[257]);
  assign t[196] = (t[258] & ~t[259]);
  assign t[197] = (t[260] & ~t[261]);
  assign t[198] = (t[262] & ~t[263]);
  assign t[199] = (t[264] & ~t[265]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[266] & ~t[267]);
  assign t[201] = (t[268] & ~t[269]);
  assign t[202] = (t[270] & ~t[271]);
  assign t[203] = (t[272] & ~t[273]);
  assign t[204] = t[274] ^ x[2];
  assign t[205] = t[275] ^ x[1];
  assign t[206] = t[276] ^ x[10];
  assign t[207] = t[277] ^ x[9];
  assign t[208] = t[278] ^ x[13];
  assign t[209] = t[279] ^ x[12];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[16];
  assign t[211] = t[281] ^ x[15];
  assign t[212] = t[282] ^ x[19];
  assign t[213] = t[283] ^ x[18];
  assign t[214] = t[284] ^ x[22];
  assign t[215] = t[285] ^ x[21];
  assign t[216] = t[286] ^ x[25];
  assign t[217] = t[287] ^ x[24];
  assign t[218] = t[288] ^ x[30];
  assign t[219] = t[289] ^ x[29];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[33];
  assign t[221] = t[291] ^ x[32];
  assign t[222] = t[292] ^ x[38];
  assign t[223] = t[293] ^ x[37];
  assign t[224] = t[294] ^ x[41];
  assign t[225] = t[295] ^ x[40];
  assign t[226] = t[296] ^ x[44];
  assign t[227] = t[297] ^ x[43];
  assign t[228] = t[298] ^ x[47];
  assign t[229] = t[299] ^ x[46];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[50];
  assign t[231] = t[301] ^ x[49];
  assign t[232] = t[302] ^ x[55];
  assign t[233] = t[303] ^ x[54];
  assign t[234] = t[304] ^ x[58];
  assign t[235] = t[305] ^ x[57];
  assign t[236] = t[306] ^ x[63];
  assign t[237] = t[307] ^ x[62];
  assign t[238] = t[308] ^ x[66];
  assign t[239] = t[309] ^ x[65];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[69];
  assign t[241] = t[311] ^ x[68];
  assign t[242] = t[312] ^ x[72];
  assign t[243] = t[313] ^ x[71];
  assign t[244] = t[314] ^ x[75];
  assign t[245] = t[315] ^ x[74];
  assign t[246] = t[316] ^ x[80];
  assign t[247] = t[317] ^ x[79];
  assign t[248] = t[318] ^ x[83];
  assign t[249] = t[319] ^ x[82];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[88];
  assign t[251] = t[321] ^ x[87];
  assign t[252] = t[322] ^ x[91];
  assign t[253] = t[323] ^ x[90];
  assign t[254] = t[324] ^ x[94];
  assign t[255] = t[325] ^ x[93];
  assign t[256] = t[326] ^ x[97];
  assign t[257] = t[327] ^ x[96];
  assign t[258] = t[328] ^ x[100];
  assign t[259] = t[329] ^ x[99];
  assign t[25] = ~(t[102]);
  assign t[260] = t[330] ^ x[103];
  assign t[261] = t[331] ^ x[102];
  assign t[262] = t[332] ^ x[106];
  assign t[263] = t[333] ^ x[105];
  assign t[264] = t[334] ^ x[109];
  assign t[265] = t[335] ^ x[108];
  assign t[266] = t[336] ^ x[112];
  assign t[267] = t[337] ^ x[111];
  assign t[268] = t[338] ^ x[115];
  assign t[269] = t[339] ^ x[114];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[118];
  assign t[271] = t[341] ^ x[117];
  assign t[272] = t[342] ^ x[121];
  assign t[273] = t[343] ^ x[120];
  assign t[274] = (x[0]);
  assign t[275] = (x[0]);
  assign t[276] = (x[8]);
  assign t[277] = (x[8]);
  assign t[278] = (x[11]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[14]);
  assign t[281] = (x[14]);
  assign t[282] = (x[17]);
  assign t[283] = (x[17]);
  assign t[284] = (x[20]);
  assign t[285] = (x[20]);
  assign t[286] = (x[23]);
  assign t[287] = (x[23]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[36]);
  assign t[293] = (x[36]);
  assign t[294] = (x[39]);
  assign t[295] = (x[39]);
  assign t[296] = (x[42]);
  assign t[297] = (x[42]);
  assign t[298] = (x[45]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[53]);
  assign t[303] = (x[53]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[61]);
  assign t[307] = (x[61]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[104] & t[46]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[70]);
  assign t[313] = (x[70]);
  assign t[314] = (x[73]);
  assign t[315] = (x[73]);
  assign t[316] = (x[78]);
  assign t[317] = (x[78]);
  assign t[318] = (x[81]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[105] & t[47]);
  assign t[320] = (x[86]);
  assign t[321] = (x[86]);
  assign t[322] = (x[89]);
  assign t[323] = (x[89]);
  assign t[324] = (x[92]);
  assign t[325] = (x[92]);
  assign t[326] = (x[95]);
  assign t[327] = (x[95]);
  assign t[328] = (x[98]);
  assign t[329] = (x[98]);
  assign t[32] = t[18] ? x[27] : x[26];
  assign t[330] = (x[101]);
  assign t[331] = (x[101]);
  assign t[332] = (x[104]);
  assign t[333] = (x[104]);
  assign t[334] = (x[107]);
  assign t[335] = (x[107]);
  assign t[336] = (x[110]);
  assign t[337] = (x[110]);
  assign t[338] = (x[113]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[116]);
  assign t[341] = (x[116]);
  assign t[342] = (x[119]);
  assign t[343] = (x[119]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[36];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[56];
  assign t[38] = ~(t[106] & t[57]);
  assign t[39] = ~(t[107] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[35] : x[34];
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[42];
  assign t[46] = ~(t[108]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[73] ? x[52] : x[51];
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = t[18] ? x[60] : x[59];
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[73] ? x[77] : x[76];
  assign t[64] = ~(t[83] & t[84]);
  assign t[65] = ~(t[120] & t[85]);
  assign t[66] = ~(t[121] & t[86]);
  assign t[67] = t[73] ? x[85] : x[84];
  assign t[68] = ~(t[104]);
  assign t[69] = ~(t[122]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[25]);
  assign t[74] = ~(t[124]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[132]);
  assign t[91] = ~(t[132] & t[97]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[133]);
  assign t[95] = ~(t[133] & t[98]);
  assign t[96] = ~(t[120]);
  assign t[97] = ~(t[125]);
  assign t[98] = ~(t[129]);
  assign t[99] = (t[134]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind216(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[115] & t[116]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[156]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[155] & t[154]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[58] ^ t[34];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[61] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[128]);
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = ~(t[78] & t[129]);
  assign t[54] = t[18] ? x[43] : x[42];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[83] & t[130]);
  assign t[58] = t[122] ? x[48] : x[47];
  assign t[59] = ~(t[131]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[132]);
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[49] ? x[62] : x[61];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[135]);
  assign t[69] = t[49] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] & t[96]);
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[101] & t[102]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[103] & t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[104] & t[105]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[110] & t[111]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [151:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[115] & t[116]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[156]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[155] & t[154]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[2];
  assign t[165] = t[210] ^ x[10];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[27];
  assign t[171] = t[216] ^ x[32];
  assign t[172] = t[217] ^ x[35];
  assign t[173] = t[218] ^ x[38];
  assign t[174] = t[219] ^ x[41];
  assign t[175] = t[220] ^ x[46];
  assign t[176] = t[221] ^ x[51];
  assign t[177] = t[222] ^ x[54];
  assign t[178] = t[223] ^ x[57];
  assign t[179] = t[224] ^ x[60];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[65];
  assign t[181] = t[226] ^ x[70];
  assign t[182] = t[227] ^ x[73];
  assign t[183] = t[228] ^ x[76];
  assign t[184] = t[229] ^ x[79];
  assign t[185] = t[230] ^ x[82];
  assign t[186] = t[231] ^ x[85];
  assign t[187] = t[232] ^ x[88];
  assign t[188] = t[233] ^ x[91];
  assign t[189] = t[234] ^ x[94];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[100];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[106];
  assign t[194] = t[239] ^ x[109];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[115];
  assign t[197] = t[242] ^ x[118];
  assign t[198] = t[243] ^ x[121];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[127];
  assign t[201] = t[246] ^ x[130];
  assign t[202] = t[247] ^ x[133];
  assign t[203] = t[248] ^ x[136];
  assign t[204] = t[249] ^ x[139];
  assign t[205] = t[250] ^ x[142];
  assign t[206] = t[251] ^ x[145];
  assign t[207] = t[252] ^ x[148];
  assign t[208] = t[253] ^ x[151];
  assign t[209] = (t[254] & ~t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[256] & ~t[257]);
  assign t[211] = (t[258] & ~t[259]);
  assign t[212] = (t[260] & ~t[261]);
  assign t[213] = (t[262] & ~t[263]);
  assign t[214] = (t[264] & ~t[265]);
  assign t[215] = (t[266] & ~t[267]);
  assign t[216] = (t[268] & ~t[269]);
  assign t[217] = (t[270] & ~t[271]);
  assign t[218] = (t[272] & ~t[273]);
  assign t[219] = (t[274] & ~t[275]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[276] & ~t[277]);
  assign t[221] = (t[278] & ~t[279]);
  assign t[222] = (t[280] & ~t[281]);
  assign t[223] = (t[282] & ~t[283]);
  assign t[224] = (t[284] & ~t[285]);
  assign t[225] = (t[286] & ~t[287]);
  assign t[226] = (t[288] & ~t[289]);
  assign t[227] = (t[290] & ~t[291]);
  assign t[228] = (t[292] & ~t[293]);
  assign t[229] = (t[294] & ~t[295]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[296] & ~t[297]);
  assign t[231] = (t[298] & ~t[299]);
  assign t[232] = (t[300] & ~t[301]);
  assign t[233] = (t[302] & ~t[303]);
  assign t[234] = (t[304] & ~t[305]);
  assign t[235] = (t[306] & ~t[307]);
  assign t[236] = (t[308] & ~t[309]);
  assign t[237] = (t[310] & ~t[311]);
  assign t[238] = (t[312] & ~t[313]);
  assign t[239] = (t[314] & ~t[315]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[316] & ~t[317]);
  assign t[241] = (t[318] & ~t[319]);
  assign t[242] = (t[320] & ~t[321]);
  assign t[243] = (t[322] & ~t[323]);
  assign t[244] = (t[324] & ~t[325]);
  assign t[245] = (t[326] & ~t[327]);
  assign t[246] = (t[328] & ~t[329]);
  assign t[247] = (t[330] & ~t[331]);
  assign t[248] = (t[332] & ~t[333]);
  assign t[249] = (t[334] & ~t[335]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[336] & ~t[337]);
  assign t[251] = (t[338] & ~t[339]);
  assign t[252] = (t[340] & ~t[341]);
  assign t[253] = (t[342] & ~t[343]);
  assign t[254] = t[344] ^ x[2];
  assign t[255] = t[345] ^ x[1];
  assign t[256] = t[346] ^ x[10];
  assign t[257] = t[347] ^ x[9];
  assign t[258] = t[348] ^ x[13];
  assign t[259] = t[349] ^ x[12];
  assign t[25] = ~(t[122]);
  assign t[260] = t[350] ^ x[16];
  assign t[261] = t[351] ^ x[15];
  assign t[262] = t[352] ^ x[19];
  assign t[263] = t[353] ^ x[18];
  assign t[264] = t[354] ^ x[22];
  assign t[265] = t[355] ^ x[21];
  assign t[266] = t[356] ^ x[27];
  assign t[267] = t[357] ^ x[26];
  assign t[268] = t[358] ^ x[32];
  assign t[269] = t[359] ^ x[31];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[35];
  assign t[271] = t[361] ^ x[34];
  assign t[272] = t[362] ^ x[38];
  assign t[273] = t[363] ^ x[37];
  assign t[274] = t[364] ^ x[41];
  assign t[275] = t[365] ^ x[40];
  assign t[276] = t[366] ^ x[46];
  assign t[277] = t[367] ^ x[45];
  assign t[278] = t[368] ^ x[51];
  assign t[279] = t[369] ^ x[50];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[54];
  assign t[281] = t[371] ^ x[53];
  assign t[282] = t[372] ^ x[57];
  assign t[283] = t[373] ^ x[56];
  assign t[284] = t[374] ^ x[60];
  assign t[285] = t[375] ^ x[59];
  assign t[286] = t[376] ^ x[65];
  assign t[287] = t[377] ^ x[64];
  assign t[288] = t[378] ^ x[70];
  assign t[289] = t[379] ^ x[69];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[73];
  assign t[291] = t[381] ^ x[72];
  assign t[292] = t[382] ^ x[76];
  assign t[293] = t[383] ^ x[75];
  assign t[294] = t[384] ^ x[79];
  assign t[295] = t[385] ^ x[78];
  assign t[296] = t[386] ^ x[82];
  assign t[297] = t[387] ^ x[81];
  assign t[298] = t[388] ^ x[85];
  assign t[299] = t[389] ^ x[84];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[88];
  assign t[301] = t[391] ^ x[87];
  assign t[302] = t[392] ^ x[91];
  assign t[303] = t[393] ^ x[90];
  assign t[304] = t[394] ^ x[94];
  assign t[305] = t[395] ^ x[93];
  assign t[306] = t[396] ^ x[97];
  assign t[307] = t[397] ^ x[96];
  assign t[308] = t[398] ^ x[100];
  assign t[309] = t[399] ^ x[99];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[103];
  assign t[311] = t[401] ^ x[102];
  assign t[312] = t[402] ^ x[106];
  assign t[313] = t[403] ^ x[105];
  assign t[314] = t[404] ^ x[109];
  assign t[315] = t[405] ^ x[108];
  assign t[316] = t[406] ^ x[112];
  assign t[317] = t[407] ^ x[111];
  assign t[318] = t[408] ^ x[115];
  assign t[319] = t[409] ^ x[114];
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = t[410] ^ x[118];
  assign t[321] = t[411] ^ x[117];
  assign t[322] = t[412] ^ x[121];
  assign t[323] = t[413] ^ x[120];
  assign t[324] = t[414] ^ x[124];
  assign t[325] = t[415] ^ x[123];
  assign t[326] = t[416] ^ x[127];
  assign t[327] = t[417] ^ x[126];
  assign t[328] = t[418] ^ x[130];
  assign t[329] = t[419] ^ x[129];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[133];
  assign t[331] = t[421] ^ x[132];
  assign t[332] = t[422] ^ x[136];
  assign t[333] = t[423] ^ x[135];
  assign t[334] = t[424] ^ x[139];
  assign t[335] = t[425] ^ x[138];
  assign t[336] = t[426] ^ x[142];
  assign t[337] = t[427] ^ x[141];
  assign t[338] = t[428] ^ x[145];
  assign t[339] = t[429] ^ x[144];
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = t[430] ^ x[148];
  assign t[341] = t[431] ^ x[147];
  assign t[342] = t[432] ^ x[151];
  assign t[343] = t[433] ^ x[150];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[8]);
  assign t[347] = (x[8]);
  assign t[348] = (x[11]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[14]);
  assign t[351] = (x[14]);
  assign t[352] = (x[17]);
  assign t[353] = (x[17]);
  assign t[354] = (x[20]);
  assign t[355] = (x[20]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[30]);
  assign t[359] = (x[30]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[33]);
  assign t[361] = (x[33]);
  assign t[362] = (x[36]);
  assign t[363] = (x[36]);
  assign t[364] = (x[39]);
  assign t[365] = (x[39]);
  assign t[366] = (x[44]);
  assign t[367] = (x[44]);
  assign t[368] = (x[49]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[52]);
  assign t[371] = (x[52]);
  assign t[372] = (x[55]);
  assign t[373] = (x[55]);
  assign t[374] = (x[58]);
  assign t[375] = (x[58]);
  assign t[376] = (x[63]);
  assign t[377] = (x[63]);
  assign t[378] = (x[68]);
  assign t[379] = (x[68]);
  assign t[37] = t[58] ^ t[34];
  assign t[380] = (x[71]);
  assign t[381] = (x[71]);
  assign t[382] = (x[74]);
  assign t[383] = (x[74]);
  assign t[384] = (x[77]);
  assign t[385] = (x[77]);
  assign t[386] = (x[80]);
  assign t[387] = (x[80]);
  assign t[388] = (x[83]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[86]);
  assign t[391] = (x[86]);
  assign t[392] = (x[89]);
  assign t[393] = (x[89]);
  assign t[394] = (x[92]);
  assign t[395] = (x[92]);
  assign t[396] = (x[95]);
  assign t[397] = (x[95]);
  assign t[398] = (x[98]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[61] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[101]);
  assign t[401] = (x[101]);
  assign t[402] = (x[104]);
  assign t[403] = (x[104]);
  assign t[404] = (x[107]);
  assign t[405] = (x[107]);
  assign t[406] = (x[110]);
  assign t[407] = (x[110]);
  assign t[408] = (x[113]);
  assign t[409] = (x[113]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[116]);
  assign t[411] = (x[116]);
  assign t[412] = (x[119]);
  assign t[413] = (x[119]);
  assign t[414] = (x[122]);
  assign t[415] = (x[122]);
  assign t[416] = (x[125]);
  assign t[417] = (x[125]);
  assign t[418] = (x[128]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[131]);
  assign t[421] = (x[131]);
  assign t[422] = (x[134]);
  assign t[423] = (x[134]);
  assign t[424] = (x[137]);
  assign t[425] = (x[137]);
  assign t[426] = (x[140]);
  assign t[427] = (x[140]);
  assign t[428] = (x[143]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[146]);
  assign t[432] = (x[149]);
  assign t[433] = (x[149]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[128]);
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = ~(t[78] & t[129]);
  assign t[54] = t[18] ? x[43] : x[42];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[83] & t[130]);
  assign t[58] = t[122] ? x[48] : x[47];
  assign t[59] = ~(t[131]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[132]);
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[49] ? x[62] : x[61];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[135]);
  assign t[69] = t[49] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] & t[96]);
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[101] & t[102]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[103] & t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[104] & t[105]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[110] & t[111]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[58] ^ t[34];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[18] ? x[43] : x[42];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = t[82] | t[121];
  assign t[58] = t[18] ? x[48] : x[47];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[83] | t[59]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[124];
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = t[89] | t[125];
  assign t[66] = t[90] ? x[62] : x[61];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = t[93] | t[126];
  assign t[69] = t[90] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[98] & t[99]);
  assign t[79] = t[100] | t[132];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[101] | t[80]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[102] | t[84]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[103] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[25]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[58] ^ t[34];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[18] ? x[43] : x[42];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = t[82] | t[121];
  assign t[58] = t[18] ? x[48] : x[47];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[83] | t[59]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[124];
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = t[89] | t[125];
  assign t[66] = t[90] ? x[62] : x[61];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = t[93] | t[126];
  assign t[69] = t[90] ? x[67] : x[66];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[98] & t[99]);
  assign t[79] = t[100] | t[132];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[101] | t[80]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[102] | t[84]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[103] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[25]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [151:0] x;
 output y;

 wire [515:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = t[135] ? x[84] : x[83];
  assign t[101] = ~(t[139] & t[140]);
  assign t[102] = ~(t[225]);
  assign t[103] = ~(t[213] | t[214]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[227]);
  assign t[106] = ~(t[141] | t[142]);
  assign t[107] = ~(t[139] & t[143]);
  assign t[108] = ~(t[228]);
  assign t[109] = ~(t[229]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[144] | t[145]);
  assign t[111] = ~(t[146] | t[147]);
  assign t[112] = ~(t[230] | t[148]);
  assign t[113] = t[149] ? x[104] : x[103];
  assign t[114] = ~(t[150] & t[151]);
  assign t[115] = ~(t[231]);
  assign t[116] = ~(t[232]);
  assign t[117] = ~(t[152] | t[153]);
  assign t[118] = ~(t[154] | t[155]);
  assign t[119] = ~(t[233] | t[156]);
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ? x[115] : x[114];
  assign t[121] = ~(t[157] & t[143]);
  assign t[122] = ~(t[204]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[81] | t[161]);
  assign t[126] = ~(t[81] | t[162]);
  assign t[127] = ~(x[4] & t[163]);
  assign t[128] = ~(t[205] & t[164]);
  assign t[129] = ~(t[234]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[219] | t[220]);
  assign t[131] = ~(t[157] & t[139]);
  assign t[132] = ~(t[81] | t[165]);
  assign t[133] = ~(t[235]);
  assign t[134] = ~(t[221] | t[222]);
  assign t[135] = ~(t[49]);
  assign t[136] = ~(t[166] | t[167]);
  assign t[137] = ~(t[236]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[168] | t[167]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[169] | t[170]);
  assign t[141] = ~(t[237]);
  assign t[142] = ~(t[226] | t[227]);
  assign t[143] = ~(t[171] & t[172]);
  assign t[144] = ~(t[238]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[239]);
  assign t[147] = ~(t[240]);
  assign t[148] = ~(t[173] | t[174]);
  assign t[149] = ~(t[49]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[175] | t[176]);
  assign t[151] = ~(t[177] & t[178]);
  assign t[152] = ~(t[241]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[179] | t[180]);
  assign t[157] = ~(t[50] | t[169]);
  assign t[158] = ~(x[4] | t[203]);
  assign t[159] = ~(t[205]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[4] & t[203];
  assign t[161] = t[202] ? t[182] : t[181];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[203] | t[205]);
  assign t[164] = ~(x[4] | t[185]);
  assign t[165] = t[202] ? t[123] : t[124];
  assign t[166] = ~(t[122] | t[186]);
  assign t[167] = ~(t[122] | t[187]);
  assign t[168] = ~(t[122] | t[188]);
  assign t[169] = ~(t[189] & t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[151] & t[191]);
  assign t[171] = ~(t[203] | t[159]);
  assign t[172] = t[81] & t[202];
  assign t[173] = ~(t[244]);
  assign t[174] = ~(t[239] | t[240]);
  assign t[175] = ~(t[192] & t[143]);
  assign t[176] = t[52] | t[193];
  assign t[177] = t[205] & t[194];
  assign t[178] = t[158] | t[160];
  assign t[179] = ~(t[245]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[242] | t[243]);
  assign t[181] = ~(t[164] & t[159]);
  assign t[182] = ~(x[4] & t[171]);
  assign t[183] = ~(t[158] & t[205]);
  assign t[184] = ~(t[160] & t[159]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[123] : t[184];
  assign t[187] = t[202] ? t[181] : t[127];
  assign t[188] = t[202] ? t[184] : t[123];
  assign t[189] = ~(t[166] | t[195]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[122] & t[196]);
  assign t[191] = t[122] | t[197];
  assign t[192] = ~(t[194] & t[198]);
  assign t[193] = ~(t[81] | t[199]);
  assign t[194] = ~(t[122] | t[202]);
  assign t[195] = ~(t[81] | t[200]);
  assign t[196] = ~(t[127] & t[128]);
  assign t[197] = t[202] ? t[127] : t[181];
  assign t[198] = ~(t[128] & t[182]);
  assign t[199] = t[202] ? t[183] : t[184];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[181] : t[182];
  assign t[201] = (t[246]);
  assign t[202] = (t[247]);
  assign t[203] = (t[248]);
  assign t[204] = (t[249]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = t[291] ^ x[2];
  assign t[247] = t[292] ^ x[10];
  assign t[248] = t[293] ^ x[13];
  assign t[249] = t[294] ^ x[16];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[19];
  assign t[251] = t[296] ^ x[22];
  assign t[252] = t[297] ^ x[25];
  assign t[253] = t[298] ^ x[28];
  assign t[254] = t[299] ^ x[31];
  assign t[255] = t[300] ^ x[34];
  assign t[256] = t[301] ^ x[39];
  assign t[257] = t[302] ^ x[42];
  assign t[258] = t[303] ^ x[45];
  assign t[259] = t[304] ^ x[48];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[51];
  assign t[261] = t[306] ^ x[56];
  assign t[262] = t[307] ^ x[59];
  assign t[263] = t[308] ^ x[62];
  assign t[264] = t[309] ^ x[65];
  assign t[265] = t[310] ^ x[68];
  assign t[266] = t[311] ^ x[71];
  assign t[267] = t[312] ^ x[74];
  assign t[268] = t[313] ^ x[79];
  assign t[269] = t[314] ^ x[82];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[87];
  assign t[271] = t[316] ^ x[90];
  assign t[272] = t[317] ^ x[93];
  assign t[273] = t[318] ^ x[96];
  assign t[274] = t[319] ^ x[99];
  assign t[275] = t[320] ^ x[102];
  assign t[276] = t[321] ^ x[107];
  assign t[277] = t[322] ^ x[110];
  assign t[278] = t[323] ^ x[113];
  assign t[279] = t[324] ^ x[118];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[121];
  assign t[281] = t[326] ^ x[124];
  assign t[282] = t[327] ^ x[127];
  assign t[283] = t[328] ^ x[130];
  assign t[284] = t[329] ^ x[133];
  assign t[285] = t[330] ^ x[136];
  assign t[286] = t[331] ^ x[139];
  assign t[287] = t[332] ^ x[142];
  assign t[288] = t[333] ^ x[145];
  assign t[289] = t[334] ^ x[148];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[151];
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[354] & ~t[355]);
  assign t[301] = (t[356] & ~t[357]);
  assign t[302] = (t[358] & ~t[359]);
  assign t[303] = (t[360] & ~t[361]);
  assign t[304] = (t[362] & ~t[363]);
  assign t[305] = (t[364] & ~t[365]);
  assign t[306] = (t[366] & ~t[367]);
  assign t[307] = (t[368] & ~t[369]);
  assign t[308] = (t[370] & ~t[371]);
  assign t[309] = (t[372] & ~t[373]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[374] & ~t[375]);
  assign t[311] = (t[376] & ~t[377]);
  assign t[312] = (t[378] & ~t[379]);
  assign t[313] = (t[380] & ~t[381]);
  assign t[314] = (t[382] & ~t[383]);
  assign t[315] = (t[384] & ~t[385]);
  assign t[316] = (t[386] & ~t[387]);
  assign t[317] = (t[388] & ~t[389]);
  assign t[318] = (t[390] & ~t[391]);
  assign t[319] = (t[392] & ~t[393]);
  assign t[31] = ~(t[50]);
  assign t[320] = (t[394] & ~t[395]);
  assign t[321] = (t[396] & ~t[397]);
  assign t[322] = (t[398] & ~t[399]);
  assign t[323] = (t[400] & ~t[401]);
  assign t[324] = (t[402] & ~t[403]);
  assign t[325] = (t[404] & ~t[405]);
  assign t[326] = (t[406] & ~t[407]);
  assign t[327] = (t[408] & ~t[409]);
  assign t[328] = (t[410] & ~t[411]);
  assign t[329] = (t[412] & ~t[413]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (t[414] & ~t[415]);
  assign t[331] = (t[416] & ~t[417]);
  assign t[332] = (t[418] & ~t[419]);
  assign t[333] = (t[420] & ~t[421]);
  assign t[334] = (t[422] & ~t[423]);
  assign t[335] = (t[424] & ~t[425]);
  assign t[336] = t[426] ^ x[2];
  assign t[337] = t[427] ^ x[1];
  assign t[338] = t[428] ^ x[10];
  assign t[339] = t[429] ^ x[9];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[430] ^ x[13];
  assign t[341] = t[431] ^ x[12];
  assign t[342] = t[432] ^ x[16];
  assign t[343] = t[433] ^ x[15];
  assign t[344] = t[434] ^ x[19];
  assign t[345] = t[435] ^ x[18];
  assign t[346] = t[436] ^ x[22];
  assign t[347] = t[437] ^ x[21];
  assign t[348] = t[438] ^ x[25];
  assign t[349] = t[439] ^ x[24];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[440] ^ x[28];
  assign t[351] = t[441] ^ x[27];
  assign t[352] = t[442] ^ x[31];
  assign t[353] = t[443] ^ x[30];
  assign t[354] = t[444] ^ x[34];
  assign t[355] = t[445] ^ x[33];
  assign t[356] = t[446] ^ x[39];
  assign t[357] = t[447] ^ x[38];
  assign t[358] = t[448] ^ x[42];
  assign t[359] = t[449] ^ x[41];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[450] ^ x[45];
  assign t[361] = t[451] ^ x[44];
  assign t[362] = t[452] ^ x[48];
  assign t[363] = t[453] ^ x[47];
  assign t[364] = t[454] ^ x[51];
  assign t[365] = t[455] ^ x[50];
  assign t[366] = t[456] ^ x[56];
  assign t[367] = t[457] ^ x[55];
  assign t[368] = t[458] ^ x[59];
  assign t[369] = t[459] ^ x[58];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[460] ^ x[62];
  assign t[371] = t[461] ^ x[61];
  assign t[372] = t[462] ^ x[65];
  assign t[373] = t[463] ^ x[64];
  assign t[374] = t[464] ^ x[68];
  assign t[375] = t[465] ^ x[67];
  assign t[376] = t[466] ^ x[71];
  assign t[377] = t[467] ^ x[70];
  assign t[378] = t[468] ^ x[74];
  assign t[379] = t[469] ^ x[73];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[470] ^ x[79];
  assign t[381] = t[471] ^ x[78];
  assign t[382] = t[472] ^ x[82];
  assign t[383] = t[473] ^ x[81];
  assign t[384] = t[474] ^ x[87];
  assign t[385] = t[475] ^ x[86];
  assign t[386] = t[476] ^ x[90];
  assign t[387] = t[477] ^ x[89];
  assign t[388] = t[478] ^ x[93];
  assign t[389] = t[479] ^ x[92];
  assign t[38] = ~(t[37] ^ t[62]);
  assign t[390] = t[480] ^ x[96];
  assign t[391] = t[481] ^ x[95];
  assign t[392] = t[482] ^ x[99];
  assign t[393] = t[483] ^ x[98];
  assign t[394] = t[484] ^ x[102];
  assign t[395] = t[485] ^ x[101];
  assign t[396] = t[486] ^ x[107];
  assign t[397] = t[487] ^ x[106];
  assign t[398] = t[488] ^ x[110];
  assign t[399] = t[489] ^ x[109];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[113];
  assign t[401] = t[491] ^ x[112];
  assign t[402] = t[492] ^ x[118];
  assign t[403] = t[493] ^ x[117];
  assign t[404] = t[494] ^ x[121];
  assign t[405] = t[495] ^ x[120];
  assign t[406] = t[496] ^ x[124];
  assign t[407] = t[497] ^ x[123];
  assign t[408] = t[498] ^ x[127];
  assign t[409] = t[499] ^ x[126];
  assign t[40] = ~(t[47] ^ t[65]);
  assign t[410] = t[500] ^ x[130];
  assign t[411] = t[501] ^ x[129];
  assign t[412] = t[502] ^ x[133];
  assign t[413] = t[503] ^ x[132];
  assign t[414] = t[504] ^ x[136];
  assign t[415] = t[505] ^ x[135];
  assign t[416] = t[506] ^ x[139];
  assign t[417] = t[507] ^ x[138];
  assign t[418] = t[508] ^ x[142];
  assign t[419] = t[509] ^ x[141];
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = t[510] ^ x[145];
  assign t[421] = t[511] ^ x[144];
  assign t[422] = t[512] ^ x[148];
  assign t[423] = t[513] ^ x[147];
  assign t[424] = t[514] ^ x[151];
  assign t[425] = t[515] ^ x[150];
  assign t[426] = (x[0]);
  assign t[427] = (x[0]);
  assign t[428] = (x[8]);
  assign t[429] = (x[8]);
  assign t[42] = ~(t[207] | t[68]);
  assign t[430] = (x[11]);
  assign t[431] = (x[11]);
  assign t[432] = (x[14]);
  assign t[433] = (x[14]);
  assign t[434] = (x[17]);
  assign t[435] = (x[17]);
  assign t[436] = (x[20]);
  assign t[437] = (x[20]);
  assign t[438] = (x[23]);
  assign t[439] = (x[23]);
  assign t[43] = ~(t[69] | t[70]);
  assign t[440] = (x[26]);
  assign t[441] = (x[26]);
  assign t[442] = (x[29]);
  assign t[443] = (x[29]);
  assign t[444] = (x[32]);
  assign t[445] = (x[32]);
  assign t[446] = (x[37]);
  assign t[447] = (x[37]);
  assign t[448] = (x[40]);
  assign t[449] = (x[40]);
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[450] = (x[43]);
  assign t[451] = (x[43]);
  assign t[452] = (x[46]);
  assign t[453] = (x[46]);
  assign t[454] = (x[49]);
  assign t[455] = (x[49]);
  assign t[456] = (x[54]);
  assign t[457] = (x[54]);
  assign t[458] = (x[57]);
  assign t[459] = (x[57]);
  assign t[45] = ~(t[73] | t[74]);
  assign t[460] = (x[60]);
  assign t[461] = (x[60]);
  assign t[462] = (x[63]);
  assign t[463] = (x[63]);
  assign t[464] = (x[66]);
  assign t[465] = (x[66]);
  assign t[466] = (x[69]);
  assign t[467] = (x[69]);
  assign t[468] = (x[72]);
  assign t[469] = (x[72]);
  assign t[46] = ~(t[75] ^ t[76]);
  assign t[470] = (x[77]);
  assign t[471] = (x[77]);
  assign t[472] = (x[80]);
  assign t[473] = (x[80]);
  assign t[474] = (x[85]);
  assign t[475] = (x[85]);
  assign t[476] = (x[88]);
  assign t[477] = (x[88]);
  assign t[478] = (x[91]);
  assign t[479] = (x[91]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[94]);
  assign t[481] = (x[94]);
  assign t[482] = (x[97]);
  assign t[483] = (x[97]);
  assign t[484] = (x[100]);
  assign t[485] = (x[100]);
  assign t[486] = (x[105]);
  assign t[487] = (x[105]);
  assign t[488] = (x[108]);
  assign t[489] = (x[108]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = (x[111]);
  assign t[491] = (x[111]);
  assign t[492] = (x[116]);
  assign t[493] = (x[116]);
  assign t[494] = (x[119]);
  assign t[495] = (x[119]);
  assign t[496] = (x[122]);
  assign t[497] = (x[122]);
  assign t[498] = (x[125]);
  assign t[499] = (x[125]);
  assign t[49] = ~(t[204]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[128]);
  assign t[501] = (x[128]);
  assign t[502] = (x[131]);
  assign t[503] = (x[131]);
  assign t[504] = (x[134]);
  assign t[505] = (x[134]);
  assign t[506] = (x[137]);
  assign t[507] = (x[137]);
  assign t[508] = (x[140]);
  assign t[509] = (x[140]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (x[143]);
  assign t[511] = (x[143]);
  assign t[512] = (x[146]);
  assign t[513] = (x[146]);
  assign t[514] = (x[149]);
  assign t[515] = (x[149]);
  assign t[51] = ~(t[83]);
  assign t[52] = ~(t[81] | t[84]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[85] | t[86]);
  assign t[56] = ~(t[87] | t[88]);
  assign t[57] = ~(t[210] | t[89]);
  assign t[58] = t[30] ? x[36] : x[35];
  assign t[59] = ~(t[90] & t[91]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[92] | t[93]);
  assign t[61] = ~(t[211] | t[94]);
  assign t[62] = ~(t[95] ^ t[96]);
  assign t[63] = ~(t[97] | t[98]);
  assign t[64] = ~(t[212] | t[99]);
  assign t[65] = ~(t[100] ^ t[101]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[214]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[104] | t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[215] | t[106]);
  assign t[71] = t[30] ? x[53] : x[52];
  assign t[72] = t[107] | t[52];
  assign t[73] = ~(t[108] | t[109]);
  assign t[74] = ~(t[216] | t[110]);
  assign t[75] = ~(t[111] | t[112]);
  assign t[76] = ~(t[113] ^ t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[217] | t[117]);
  assign t[79] = ~(t[118] | t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[120] ^ t[121]);
  assign t[81] = ~(t[122]);
  assign t[82] = t[202] ? t[124] : t[123];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[202] ? t[128] : t[127];
  assign t[85] = ~(t[218]);
  assign t[86] = ~(t[208] | t[209]);
  assign t[87] = ~(t[219]);
  assign t[88] = ~(t[220]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] | t[131]);
  assign t[91] = ~(t[132]);
  assign t[92] = ~(t[221]);
  assign t[93] = ~(t[222]);
  assign t[94] = ~(t[133] | t[134]);
  assign t[95] = t[135] ? x[76] : x[75];
  assign t[96] = ~(t[136] & t[32]);
  assign t[97] = ~(t[223]);
  assign t[98] = ~(t[224]);
  assign t[99] = ~(t[137] | t[138]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind221(x, y);
 input [151:0] x;
 output y;

 wire [515:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = t[135] ? x[84] : x[83];
  assign t[101] = ~(t[139] & t[140]);
  assign t[102] = ~(t[225]);
  assign t[103] = ~(t[213] | t[214]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[227]);
  assign t[106] = ~(t[141] | t[142]);
  assign t[107] = ~(t[139] & t[143]);
  assign t[108] = ~(t[228]);
  assign t[109] = ~(t[229]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[144] | t[145]);
  assign t[111] = ~(t[146] | t[147]);
  assign t[112] = ~(t[230] | t[148]);
  assign t[113] = t[149] ? x[104] : x[103];
  assign t[114] = ~(t[150] & t[151]);
  assign t[115] = ~(t[231]);
  assign t[116] = ~(t[232]);
  assign t[117] = ~(t[152] | t[153]);
  assign t[118] = ~(t[154] | t[155]);
  assign t[119] = ~(t[233] | t[156]);
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ? x[115] : x[114];
  assign t[121] = ~(t[157] & t[143]);
  assign t[122] = ~(t[204]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[81] | t[161]);
  assign t[126] = ~(t[81] | t[162]);
  assign t[127] = ~(x[4] & t[163]);
  assign t[128] = ~(t[205] & t[164]);
  assign t[129] = ~(t[234]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[219] | t[220]);
  assign t[131] = ~(t[157] & t[139]);
  assign t[132] = ~(t[81] | t[165]);
  assign t[133] = ~(t[235]);
  assign t[134] = ~(t[221] | t[222]);
  assign t[135] = ~(t[49]);
  assign t[136] = ~(t[166] | t[167]);
  assign t[137] = ~(t[236]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[168] | t[167]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[169] | t[170]);
  assign t[141] = ~(t[237]);
  assign t[142] = ~(t[226] | t[227]);
  assign t[143] = ~(t[171] & t[172]);
  assign t[144] = ~(t[238]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[239]);
  assign t[147] = ~(t[240]);
  assign t[148] = ~(t[173] | t[174]);
  assign t[149] = ~(t[49]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[175] | t[176]);
  assign t[151] = ~(t[177] & t[178]);
  assign t[152] = ~(t[241]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[179] | t[180]);
  assign t[157] = ~(t[50] | t[169]);
  assign t[158] = ~(x[4] | t[203]);
  assign t[159] = ~(t[205]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[4] & t[203];
  assign t[161] = t[202] ? t[182] : t[181];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[203] | t[205]);
  assign t[164] = ~(x[4] | t[185]);
  assign t[165] = t[202] ? t[123] : t[124];
  assign t[166] = ~(t[122] | t[186]);
  assign t[167] = ~(t[122] | t[187]);
  assign t[168] = ~(t[122] | t[188]);
  assign t[169] = ~(t[189] & t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[151] & t[191]);
  assign t[171] = ~(t[203] | t[159]);
  assign t[172] = t[81] & t[202];
  assign t[173] = ~(t[244]);
  assign t[174] = ~(t[239] | t[240]);
  assign t[175] = ~(t[192] & t[143]);
  assign t[176] = t[52] | t[193];
  assign t[177] = t[205] & t[194];
  assign t[178] = t[158] | t[160];
  assign t[179] = ~(t[245]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[242] | t[243]);
  assign t[181] = ~(t[164] & t[159]);
  assign t[182] = ~(x[4] & t[171]);
  assign t[183] = ~(t[158] & t[205]);
  assign t[184] = ~(t[160] & t[159]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[123] : t[184];
  assign t[187] = t[202] ? t[181] : t[127];
  assign t[188] = t[202] ? t[184] : t[123];
  assign t[189] = ~(t[166] | t[195]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[122] & t[196]);
  assign t[191] = t[122] | t[197];
  assign t[192] = ~(t[194] & t[198]);
  assign t[193] = ~(t[81] | t[199]);
  assign t[194] = ~(t[122] | t[202]);
  assign t[195] = ~(t[81] | t[200]);
  assign t[196] = ~(t[127] & t[128]);
  assign t[197] = t[202] ? t[127] : t[181];
  assign t[198] = ~(t[128] & t[182]);
  assign t[199] = t[202] ? t[183] : t[184];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[181] : t[182];
  assign t[201] = (t[246]);
  assign t[202] = (t[247]);
  assign t[203] = (t[248]);
  assign t[204] = (t[249]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = t[291] ^ x[2];
  assign t[247] = t[292] ^ x[10];
  assign t[248] = t[293] ^ x[13];
  assign t[249] = t[294] ^ x[16];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[19];
  assign t[251] = t[296] ^ x[22];
  assign t[252] = t[297] ^ x[25];
  assign t[253] = t[298] ^ x[28];
  assign t[254] = t[299] ^ x[31];
  assign t[255] = t[300] ^ x[34];
  assign t[256] = t[301] ^ x[39];
  assign t[257] = t[302] ^ x[42];
  assign t[258] = t[303] ^ x[45];
  assign t[259] = t[304] ^ x[48];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[51];
  assign t[261] = t[306] ^ x[56];
  assign t[262] = t[307] ^ x[59];
  assign t[263] = t[308] ^ x[62];
  assign t[264] = t[309] ^ x[65];
  assign t[265] = t[310] ^ x[68];
  assign t[266] = t[311] ^ x[71];
  assign t[267] = t[312] ^ x[74];
  assign t[268] = t[313] ^ x[79];
  assign t[269] = t[314] ^ x[82];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[87];
  assign t[271] = t[316] ^ x[90];
  assign t[272] = t[317] ^ x[93];
  assign t[273] = t[318] ^ x[96];
  assign t[274] = t[319] ^ x[99];
  assign t[275] = t[320] ^ x[102];
  assign t[276] = t[321] ^ x[107];
  assign t[277] = t[322] ^ x[110];
  assign t[278] = t[323] ^ x[113];
  assign t[279] = t[324] ^ x[118];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[121];
  assign t[281] = t[326] ^ x[124];
  assign t[282] = t[327] ^ x[127];
  assign t[283] = t[328] ^ x[130];
  assign t[284] = t[329] ^ x[133];
  assign t[285] = t[330] ^ x[136];
  assign t[286] = t[331] ^ x[139];
  assign t[287] = t[332] ^ x[142];
  assign t[288] = t[333] ^ x[145];
  assign t[289] = t[334] ^ x[148];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[151];
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[354] & ~t[355]);
  assign t[301] = (t[356] & ~t[357]);
  assign t[302] = (t[358] & ~t[359]);
  assign t[303] = (t[360] & ~t[361]);
  assign t[304] = (t[362] & ~t[363]);
  assign t[305] = (t[364] & ~t[365]);
  assign t[306] = (t[366] & ~t[367]);
  assign t[307] = (t[368] & ~t[369]);
  assign t[308] = (t[370] & ~t[371]);
  assign t[309] = (t[372] & ~t[373]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[374] & ~t[375]);
  assign t[311] = (t[376] & ~t[377]);
  assign t[312] = (t[378] & ~t[379]);
  assign t[313] = (t[380] & ~t[381]);
  assign t[314] = (t[382] & ~t[383]);
  assign t[315] = (t[384] & ~t[385]);
  assign t[316] = (t[386] & ~t[387]);
  assign t[317] = (t[388] & ~t[389]);
  assign t[318] = (t[390] & ~t[391]);
  assign t[319] = (t[392] & ~t[393]);
  assign t[31] = ~(t[50]);
  assign t[320] = (t[394] & ~t[395]);
  assign t[321] = (t[396] & ~t[397]);
  assign t[322] = (t[398] & ~t[399]);
  assign t[323] = (t[400] & ~t[401]);
  assign t[324] = (t[402] & ~t[403]);
  assign t[325] = (t[404] & ~t[405]);
  assign t[326] = (t[406] & ~t[407]);
  assign t[327] = (t[408] & ~t[409]);
  assign t[328] = (t[410] & ~t[411]);
  assign t[329] = (t[412] & ~t[413]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (t[414] & ~t[415]);
  assign t[331] = (t[416] & ~t[417]);
  assign t[332] = (t[418] & ~t[419]);
  assign t[333] = (t[420] & ~t[421]);
  assign t[334] = (t[422] & ~t[423]);
  assign t[335] = (t[424] & ~t[425]);
  assign t[336] = t[426] ^ x[2];
  assign t[337] = t[427] ^ x[1];
  assign t[338] = t[428] ^ x[10];
  assign t[339] = t[429] ^ x[9];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[430] ^ x[13];
  assign t[341] = t[431] ^ x[12];
  assign t[342] = t[432] ^ x[16];
  assign t[343] = t[433] ^ x[15];
  assign t[344] = t[434] ^ x[19];
  assign t[345] = t[435] ^ x[18];
  assign t[346] = t[436] ^ x[22];
  assign t[347] = t[437] ^ x[21];
  assign t[348] = t[438] ^ x[25];
  assign t[349] = t[439] ^ x[24];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[440] ^ x[28];
  assign t[351] = t[441] ^ x[27];
  assign t[352] = t[442] ^ x[31];
  assign t[353] = t[443] ^ x[30];
  assign t[354] = t[444] ^ x[34];
  assign t[355] = t[445] ^ x[33];
  assign t[356] = t[446] ^ x[39];
  assign t[357] = t[447] ^ x[38];
  assign t[358] = t[448] ^ x[42];
  assign t[359] = t[449] ^ x[41];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[450] ^ x[45];
  assign t[361] = t[451] ^ x[44];
  assign t[362] = t[452] ^ x[48];
  assign t[363] = t[453] ^ x[47];
  assign t[364] = t[454] ^ x[51];
  assign t[365] = t[455] ^ x[50];
  assign t[366] = t[456] ^ x[56];
  assign t[367] = t[457] ^ x[55];
  assign t[368] = t[458] ^ x[59];
  assign t[369] = t[459] ^ x[58];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[460] ^ x[62];
  assign t[371] = t[461] ^ x[61];
  assign t[372] = t[462] ^ x[65];
  assign t[373] = t[463] ^ x[64];
  assign t[374] = t[464] ^ x[68];
  assign t[375] = t[465] ^ x[67];
  assign t[376] = t[466] ^ x[71];
  assign t[377] = t[467] ^ x[70];
  assign t[378] = t[468] ^ x[74];
  assign t[379] = t[469] ^ x[73];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[470] ^ x[79];
  assign t[381] = t[471] ^ x[78];
  assign t[382] = t[472] ^ x[82];
  assign t[383] = t[473] ^ x[81];
  assign t[384] = t[474] ^ x[87];
  assign t[385] = t[475] ^ x[86];
  assign t[386] = t[476] ^ x[90];
  assign t[387] = t[477] ^ x[89];
  assign t[388] = t[478] ^ x[93];
  assign t[389] = t[479] ^ x[92];
  assign t[38] = ~(t[37] ^ t[62]);
  assign t[390] = t[480] ^ x[96];
  assign t[391] = t[481] ^ x[95];
  assign t[392] = t[482] ^ x[99];
  assign t[393] = t[483] ^ x[98];
  assign t[394] = t[484] ^ x[102];
  assign t[395] = t[485] ^ x[101];
  assign t[396] = t[486] ^ x[107];
  assign t[397] = t[487] ^ x[106];
  assign t[398] = t[488] ^ x[110];
  assign t[399] = t[489] ^ x[109];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[113];
  assign t[401] = t[491] ^ x[112];
  assign t[402] = t[492] ^ x[118];
  assign t[403] = t[493] ^ x[117];
  assign t[404] = t[494] ^ x[121];
  assign t[405] = t[495] ^ x[120];
  assign t[406] = t[496] ^ x[124];
  assign t[407] = t[497] ^ x[123];
  assign t[408] = t[498] ^ x[127];
  assign t[409] = t[499] ^ x[126];
  assign t[40] = ~(t[47] ^ t[65]);
  assign t[410] = t[500] ^ x[130];
  assign t[411] = t[501] ^ x[129];
  assign t[412] = t[502] ^ x[133];
  assign t[413] = t[503] ^ x[132];
  assign t[414] = t[504] ^ x[136];
  assign t[415] = t[505] ^ x[135];
  assign t[416] = t[506] ^ x[139];
  assign t[417] = t[507] ^ x[138];
  assign t[418] = t[508] ^ x[142];
  assign t[419] = t[509] ^ x[141];
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = t[510] ^ x[145];
  assign t[421] = t[511] ^ x[144];
  assign t[422] = t[512] ^ x[148];
  assign t[423] = t[513] ^ x[147];
  assign t[424] = t[514] ^ x[151];
  assign t[425] = t[515] ^ x[150];
  assign t[426] = (x[0]);
  assign t[427] = (x[0]);
  assign t[428] = (x[8]);
  assign t[429] = (x[8]);
  assign t[42] = ~(t[207] | t[68]);
  assign t[430] = (x[11]);
  assign t[431] = (x[11]);
  assign t[432] = (x[14]);
  assign t[433] = (x[14]);
  assign t[434] = (x[17]);
  assign t[435] = (x[17]);
  assign t[436] = (x[20]);
  assign t[437] = (x[20]);
  assign t[438] = (x[23]);
  assign t[439] = (x[23]);
  assign t[43] = ~(t[69] | t[70]);
  assign t[440] = (x[26]);
  assign t[441] = (x[26]);
  assign t[442] = (x[29]);
  assign t[443] = (x[29]);
  assign t[444] = (x[32]);
  assign t[445] = (x[32]);
  assign t[446] = (x[37]);
  assign t[447] = (x[37]);
  assign t[448] = (x[40]);
  assign t[449] = (x[40]);
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[450] = (x[43]);
  assign t[451] = (x[43]);
  assign t[452] = (x[46]);
  assign t[453] = (x[46]);
  assign t[454] = (x[49]);
  assign t[455] = (x[49]);
  assign t[456] = (x[54]);
  assign t[457] = (x[54]);
  assign t[458] = (x[57]);
  assign t[459] = (x[57]);
  assign t[45] = ~(t[73] | t[74]);
  assign t[460] = (x[60]);
  assign t[461] = (x[60]);
  assign t[462] = (x[63]);
  assign t[463] = (x[63]);
  assign t[464] = (x[66]);
  assign t[465] = (x[66]);
  assign t[466] = (x[69]);
  assign t[467] = (x[69]);
  assign t[468] = (x[72]);
  assign t[469] = (x[72]);
  assign t[46] = ~(t[75] ^ t[76]);
  assign t[470] = (x[77]);
  assign t[471] = (x[77]);
  assign t[472] = (x[80]);
  assign t[473] = (x[80]);
  assign t[474] = (x[85]);
  assign t[475] = (x[85]);
  assign t[476] = (x[88]);
  assign t[477] = (x[88]);
  assign t[478] = (x[91]);
  assign t[479] = (x[91]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[94]);
  assign t[481] = (x[94]);
  assign t[482] = (x[97]);
  assign t[483] = (x[97]);
  assign t[484] = (x[100]);
  assign t[485] = (x[100]);
  assign t[486] = (x[105]);
  assign t[487] = (x[105]);
  assign t[488] = (x[108]);
  assign t[489] = (x[108]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = (x[111]);
  assign t[491] = (x[111]);
  assign t[492] = (x[116]);
  assign t[493] = (x[116]);
  assign t[494] = (x[119]);
  assign t[495] = (x[119]);
  assign t[496] = (x[122]);
  assign t[497] = (x[122]);
  assign t[498] = (x[125]);
  assign t[499] = (x[125]);
  assign t[49] = ~(t[204]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[128]);
  assign t[501] = (x[128]);
  assign t[502] = (x[131]);
  assign t[503] = (x[131]);
  assign t[504] = (x[134]);
  assign t[505] = (x[134]);
  assign t[506] = (x[137]);
  assign t[507] = (x[137]);
  assign t[508] = (x[140]);
  assign t[509] = (x[140]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (x[143]);
  assign t[511] = (x[143]);
  assign t[512] = (x[146]);
  assign t[513] = (x[146]);
  assign t[514] = (x[149]);
  assign t[515] = (x[149]);
  assign t[51] = ~(t[83]);
  assign t[52] = ~(t[81] | t[84]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[85] | t[86]);
  assign t[56] = ~(t[87] | t[88]);
  assign t[57] = ~(t[210] | t[89]);
  assign t[58] = t[30] ? x[36] : x[35];
  assign t[59] = ~(t[90] & t[91]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[92] | t[93]);
  assign t[61] = ~(t[211] | t[94]);
  assign t[62] = ~(t[95] ^ t[96]);
  assign t[63] = ~(t[97] | t[98]);
  assign t[64] = ~(t[212] | t[99]);
  assign t[65] = ~(t[100] ^ t[101]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[214]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[104] | t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[215] | t[106]);
  assign t[71] = t[30] ? x[53] : x[52];
  assign t[72] = t[107] | t[52];
  assign t[73] = ~(t[108] | t[109]);
  assign t[74] = ~(t[216] | t[110]);
  assign t[75] = ~(t[111] | t[112]);
  assign t[76] = ~(t[113] ^ t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[217] | t[117]);
  assign t[79] = ~(t[118] | t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[120] ^ t[121]);
  assign t[81] = ~(t[122]);
  assign t[82] = t[202] ? t[124] : t[123];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[202] ? t[128] : t[127];
  assign t[85] = ~(t[218]);
  assign t[86] = ~(t[208] | t[209]);
  assign t[87] = ~(t[219]);
  assign t[88] = ~(t[220]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] | t[131]);
  assign t[91] = ~(t[132]);
  assign t[92] = ~(t[221]);
  assign t[93] = ~(t[222]);
  assign t[94] = ~(t[133] | t[134]);
  assign t[95] = t[135] ? x[76] : x[75];
  assign t[96] = ~(t[136] & t[32]);
  assign t[97] = ~(t[223]);
  assign t[98] = ~(t[224]);
  assign t[99] = ~(t[137] | t[138]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [121:0] x;
 output y;

 wire [342:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[2];
  assign t[134] = t[169] ^ x[8];
  assign t[135] = t[170] ^ x[11];
  assign t[136] = t[171] ^ x[14];
  assign t[137] = t[172] ^ x[17];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[25];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[30];
  assign t[141] = t[176] ^ x[33];
  assign t[142] = t[177] ^ x[38];
  assign t[143] = t[178] ^ x[41];
  assign t[144] = t[179] ^ x[44];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[50];
  assign t[147] = t[182] ^ x[55];
  assign t[148] = t[183] ^ x[58];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[66];
  assign t[151] = t[186] ^ x[69];
  assign t[152] = t[187] ^ x[72];
  assign t[153] = t[188] ^ x[75];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[83];
  assign t[156] = t[191] ^ x[88];
  assign t[157] = t[192] ^ x[91];
  assign t[158] = t[193] ^ x[94];
  assign t[159] = t[194] ^ x[97];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[106];
  assign t[163] = t[198] ^ x[109];
  assign t[164] = t[199] ^ x[112];
  assign t[165] = t[200] ^ x[115];
  assign t[166] = t[201] ^ x[118];
  assign t[167] = t[202] ^ x[121];
  assign t[168] = (t[203] & ~t[204]);
  assign t[169] = (t[205] & ~t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (t[207] & ~t[208]);
  assign t[171] = (t[209] & ~t[210]);
  assign t[172] = (t[211] & ~t[212]);
  assign t[173] = (t[213] & ~t[214]);
  assign t[174] = (t[215] & ~t[216]);
  assign t[175] = (t[217] & ~t[218]);
  assign t[176] = (t[219] & ~t[220]);
  assign t[177] = (t[221] & ~t[222]);
  assign t[178] = (t[223] & ~t[224]);
  assign t[179] = (t[225] & ~t[226]);
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = (t[227] & ~t[228]);
  assign t[181] = (t[229] & ~t[230]);
  assign t[182] = (t[231] & ~t[232]);
  assign t[183] = (t[233] & ~t[234]);
  assign t[184] = (t[235] & ~t[236]);
  assign t[185] = (t[237] & ~t[238]);
  assign t[186] = (t[239] & ~t[240]);
  assign t[187] = (t[241] & ~t[242]);
  assign t[188] = (t[243] & ~t[244]);
  assign t[189] = (t[245] & ~t[246]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (t[247] & ~t[248]);
  assign t[191] = (t[249] & ~t[250]);
  assign t[192] = (t[251] & ~t[252]);
  assign t[193] = (t[253] & ~t[254]);
  assign t[194] = (t[255] & ~t[256]);
  assign t[195] = (t[257] & ~t[258]);
  assign t[196] = (t[259] & ~t[260]);
  assign t[197] = (t[261] & ~t[262]);
  assign t[198] = (t[263] & ~t[264]);
  assign t[199] = (t[265] & ~t[266]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[267] & ~t[268]);
  assign t[201] = (t[269] & ~t[270]);
  assign t[202] = (t[271] & ~t[272]);
  assign t[203] = t[273] ^ x[2];
  assign t[204] = t[274] ^ x[1];
  assign t[205] = t[275] ^ x[8];
  assign t[206] = t[276] ^ x[7];
  assign t[207] = t[277] ^ x[11];
  assign t[208] = t[278] ^ x[10];
  assign t[209] = t[279] ^ x[14];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[280] ^ x[13];
  assign t[211] = t[281] ^ x[17];
  assign t[212] = t[282] ^ x[16];
  assign t[213] = t[283] ^ x[22];
  assign t[214] = t[284] ^ x[21];
  assign t[215] = t[285] ^ x[25];
  assign t[216] = t[286] ^ x[24];
  assign t[217] = t[287] ^ x[30];
  assign t[218] = t[288] ^ x[29];
  assign t[219] = t[289] ^ x[33];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[290] ^ x[32];
  assign t[221] = t[291] ^ x[38];
  assign t[222] = t[292] ^ x[37];
  assign t[223] = t[293] ^ x[41];
  assign t[224] = t[294] ^ x[40];
  assign t[225] = t[295] ^ x[44];
  assign t[226] = t[296] ^ x[43];
  assign t[227] = t[297] ^ x[47];
  assign t[228] = t[298] ^ x[46];
  assign t[229] = t[299] ^ x[50];
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = t[300] ^ x[49];
  assign t[231] = t[301] ^ x[55];
  assign t[232] = t[302] ^ x[54];
  assign t[233] = t[303] ^ x[58];
  assign t[234] = t[304] ^ x[57];
  assign t[235] = t[305] ^ x[63];
  assign t[236] = t[306] ^ x[62];
  assign t[237] = t[307] ^ x[66];
  assign t[238] = t[308] ^ x[65];
  assign t[239] = t[309] ^ x[69];
  assign t[23] = ~(t[101]);
  assign t[240] = t[310] ^ x[68];
  assign t[241] = t[311] ^ x[72];
  assign t[242] = t[312] ^ x[71];
  assign t[243] = t[313] ^ x[75];
  assign t[244] = t[314] ^ x[74];
  assign t[245] = t[315] ^ x[80];
  assign t[246] = t[316] ^ x[79];
  assign t[247] = t[317] ^ x[83];
  assign t[248] = t[318] ^ x[82];
  assign t[249] = t[319] ^ x[88];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[320] ^ x[87];
  assign t[251] = t[321] ^ x[91];
  assign t[252] = t[322] ^ x[90];
  assign t[253] = t[323] ^ x[94];
  assign t[254] = t[324] ^ x[93];
  assign t[255] = t[325] ^ x[97];
  assign t[256] = t[326] ^ x[96];
  assign t[257] = t[327] ^ x[100];
  assign t[258] = t[328] ^ x[99];
  assign t[259] = t[329] ^ x[103];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[330] ^ x[102];
  assign t[261] = t[331] ^ x[106];
  assign t[262] = t[332] ^ x[105];
  assign t[263] = t[333] ^ x[109];
  assign t[264] = t[334] ^ x[108];
  assign t[265] = t[335] ^ x[112];
  assign t[266] = t[336] ^ x[111];
  assign t[267] = t[337] ^ x[115];
  assign t[268] = t[338] ^ x[114];
  assign t[269] = t[339] ^ x[118];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[340] ^ x[117];
  assign t[271] = t[341] ^ x[121];
  assign t[272] = t[342] ^ x[120];
  assign t[273] = (x[0]);
  assign t[274] = (x[0]);
  assign t[275] = (x[6]);
  assign t[276] = (x[6]);
  assign t[277] = (x[9]);
  assign t[278] = (x[9]);
  assign t[279] = (x[12]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[12]);
  assign t[281] = (x[15]);
  assign t[282] = (x[15]);
  assign t[283] = (x[20]);
  assign t[284] = (x[20]);
  assign t[285] = (x[23]);
  assign t[286] = (x[23]);
  assign t[287] = (x[28]);
  assign t[288] = (x[28]);
  assign t[289] = (x[31]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[31]);
  assign t[291] = (x[36]);
  assign t[292] = (x[36]);
  assign t[293] = (x[39]);
  assign t[294] = (x[39]);
  assign t[295] = (x[42]);
  assign t[296] = (x[42]);
  assign t[297] = (x[45]);
  assign t[298] = (x[45]);
  assign t[299] = (x[48]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[48]);
  assign t[301] = (x[53]);
  assign t[302] = (x[53]);
  assign t[303] = (x[56]);
  assign t[304] = (x[56]);
  assign t[305] = (x[61]);
  assign t[306] = (x[61]);
  assign t[307] = (x[64]);
  assign t[308] = (x[64]);
  assign t[309] = (x[67]);
  assign t[30] = t[16] ? x[27] : x[26];
  assign t[310] = (x[67]);
  assign t[311] = (x[70]);
  assign t[312] = (x[70]);
  assign t[313] = (x[73]);
  assign t[314] = (x[73]);
  assign t[315] = (x[78]);
  assign t[316] = (x[78]);
  assign t[317] = (x[81]);
  assign t[318] = (x[81]);
  assign t[319] = (x[86]);
  assign t[31] = ~(t[46] & t[47]);
  assign t[320] = (x[86]);
  assign t[321] = (x[89]);
  assign t[322] = (x[89]);
  assign t[323] = (x[92]);
  assign t[324] = (x[92]);
  assign t[325] = (x[95]);
  assign t[326] = (x[95]);
  assign t[327] = (x[98]);
  assign t[328] = (x[98]);
  assign t[329] = (x[101]);
  assign t[32] = ~(t[48] & t[49]);
  assign t[330] = (x[101]);
  assign t[331] = (x[104]);
  assign t[332] = (x[104]);
  assign t[333] = (x[107]);
  assign t[334] = (x[107]);
  assign t[335] = (x[110]);
  assign t[336] = (x[110]);
  assign t[337] = (x[113]);
  assign t[338] = (x[113]);
  assign t[339] = (x[116]);
  assign t[33] = t[50] ^ t[40];
  assign t[340] = (x[116]);
  assign t[341] = (x[119]);
  assign t[342] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[105] & t[54]);
  assign t[37] = ~(t[106] & t[55]);
  assign t[38] = t[16] ? x[35] : x[34];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[61];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[66]);
  assign t[46] = ~(t[108] & t[67]);
  assign t[47] = ~(t[109] & t[68]);
  assign t[48] = ~(t[110] & t[69]);
  assign t[49] = ~(t[111] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[71] ? x[52] : x[51];
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[71] ? x[60] : x[59];
  assign t[54] = ~(t[114]);
  assign t[55] = ~(t[114] & t[74]);
  assign t[56] = ~(t[115] & t[75]);
  assign t[57] = ~(t[116] & t[76]);
  assign t[58] = ~(t[117] & t[77]);
  assign t[59] = ~(t[118] & t[78]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[79] ? x[77] : x[76];
  assign t[61] = ~(t[80] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[79] ? x[85] : x[84];
  assign t[65] = ~(t[84] & t[85]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[121]);
  assign t[68] = ~(t[121] & t[86]);
  assign t[69] = ~(t[122]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[23]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[105]);
  assign t[75] = ~(t[124]);
  assign t[76] = ~(t[124] & t[89]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[23]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[115]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[131]);
  assign t[92] = ~(t[131] & t[96]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[126]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [121:0] x;
 output y;

 wire [342:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[2];
  assign t[134] = t[169] ^ x[8];
  assign t[135] = t[170] ^ x[11];
  assign t[136] = t[171] ^ x[14];
  assign t[137] = t[172] ^ x[17];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[25];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[30];
  assign t[141] = t[176] ^ x[33];
  assign t[142] = t[177] ^ x[38];
  assign t[143] = t[178] ^ x[41];
  assign t[144] = t[179] ^ x[44];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[50];
  assign t[147] = t[182] ^ x[55];
  assign t[148] = t[183] ^ x[58];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[66];
  assign t[151] = t[186] ^ x[69];
  assign t[152] = t[187] ^ x[72];
  assign t[153] = t[188] ^ x[75];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[83];
  assign t[156] = t[191] ^ x[88];
  assign t[157] = t[192] ^ x[91];
  assign t[158] = t[193] ^ x[94];
  assign t[159] = t[194] ^ x[97];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[106];
  assign t[163] = t[198] ^ x[109];
  assign t[164] = t[199] ^ x[112];
  assign t[165] = t[200] ^ x[115];
  assign t[166] = t[201] ^ x[118];
  assign t[167] = t[202] ^ x[121];
  assign t[168] = (t[203] & ~t[204]);
  assign t[169] = (t[205] & ~t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (t[207] & ~t[208]);
  assign t[171] = (t[209] & ~t[210]);
  assign t[172] = (t[211] & ~t[212]);
  assign t[173] = (t[213] & ~t[214]);
  assign t[174] = (t[215] & ~t[216]);
  assign t[175] = (t[217] & ~t[218]);
  assign t[176] = (t[219] & ~t[220]);
  assign t[177] = (t[221] & ~t[222]);
  assign t[178] = (t[223] & ~t[224]);
  assign t[179] = (t[225] & ~t[226]);
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = (t[227] & ~t[228]);
  assign t[181] = (t[229] & ~t[230]);
  assign t[182] = (t[231] & ~t[232]);
  assign t[183] = (t[233] & ~t[234]);
  assign t[184] = (t[235] & ~t[236]);
  assign t[185] = (t[237] & ~t[238]);
  assign t[186] = (t[239] & ~t[240]);
  assign t[187] = (t[241] & ~t[242]);
  assign t[188] = (t[243] & ~t[244]);
  assign t[189] = (t[245] & ~t[246]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (t[247] & ~t[248]);
  assign t[191] = (t[249] & ~t[250]);
  assign t[192] = (t[251] & ~t[252]);
  assign t[193] = (t[253] & ~t[254]);
  assign t[194] = (t[255] & ~t[256]);
  assign t[195] = (t[257] & ~t[258]);
  assign t[196] = (t[259] & ~t[260]);
  assign t[197] = (t[261] & ~t[262]);
  assign t[198] = (t[263] & ~t[264]);
  assign t[199] = (t[265] & ~t[266]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (t[267] & ~t[268]);
  assign t[201] = (t[269] & ~t[270]);
  assign t[202] = (t[271] & ~t[272]);
  assign t[203] = t[273] ^ x[2];
  assign t[204] = t[274] ^ x[1];
  assign t[205] = t[275] ^ x[8];
  assign t[206] = t[276] ^ x[7];
  assign t[207] = t[277] ^ x[11];
  assign t[208] = t[278] ^ x[10];
  assign t[209] = t[279] ^ x[14];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[280] ^ x[13];
  assign t[211] = t[281] ^ x[17];
  assign t[212] = t[282] ^ x[16];
  assign t[213] = t[283] ^ x[22];
  assign t[214] = t[284] ^ x[21];
  assign t[215] = t[285] ^ x[25];
  assign t[216] = t[286] ^ x[24];
  assign t[217] = t[287] ^ x[30];
  assign t[218] = t[288] ^ x[29];
  assign t[219] = t[289] ^ x[33];
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = t[290] ^ x[32];
  assign t[221] = t[291] ^ x[38];
  assign t[222] = t[292] ^ x[37];
  assign t[223] = t[293] ^ x[41];
  assign t[224] = t[294] ^ x[40];
  assign t[225] = t[295] ^ x[44];
  assign t[226] = t[296] ^ x[43];
  assign t[227] = t[297] ^ x[47];
  assign t[228] = t[298] ^ x[46];
  assign t[229] = t[299] ^ x[50];
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = t[300] ^ x[49];
  assign t[231] = t[301] ^ x[55];
  assign t[232] = t[302] ^ x[54];
  assign t[233] = t[303] ^ x[58];
  assign t[234] = t[304] ^ x[57];
  assign t[235] = t[305] ^ x[63];
  assign t[236] = t[306] ^ x[62];
  assign t[237] = t[307] ^ x[66];
  assign t[238] = t[308] ^ x[65];
  assign t[239] = t[309] ^ x[69];
  assign t[23] = ~(t[101]);
  assign t[240] = t[310] ^ x[68];
  assign t[241] = t[311] ^ x[72];
  assign t[242] = t[312] ^ x[71];
  assign t[243] = t[313] ^ x[75];
  assign t[244] = t[314] ^ x[74];
  assign t[245] = t[315] ^ x[80];
  assign t[246] = t[316] ^ x[79];
  assign t[247] = t[317] ^ x[83];
  assign t[248] = t[318] ^ x[82];
  assign t[249] = t[319] ^ x[88];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[320] ^ x[87];
  assign t[251] = t[321] ^ x[91];
  assign t[252] = t[322] ^ x[90];
  assign t[253] = t[323] ^ x[94];
  assign t[254] = t[324] ^ x[93];
  assign t[255] = t[325] ^ x[97];
  assign t[256] = t[326] ^ x[96];
  assign t[257] = t[327] ^ x[100];
  assign t[258] = t[328] ^ x[99];
  assign t[259] = t[329] ^ x[103];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[330] ^ x[102];
  assign t[261] = t[331] ^ x[106];
  assign t[262] = t[332] ^ x[105];
  assign t[263] = t[333] ^ x[109];
  assign t[264] = t[334] ^ x[108];
  assign t[265] = t[335] ^ x[112];
  assign t[266] = t[336] ^ x[111];
  assign t[267] = t[337] ^ x[115];
  assign t[268] = t[338] ^ x[114];
  assign t[269] = t[339] ^ x[118];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[340] ^ x[117];
  assign t[271] = t[341] ^ x[121];
  assign t[272] = t[342] ^ x[120];
  assign t[273] = (x[0]);
  assign t[274] = (x[0]);
  assign t[275] = (x[6]);
  assign t[276] = (x[6]);
  assign t[277] = (x[9]);
  assign t[278] = (x[9]);
  assign t[279] = (x[12]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[12]);
  assign t[281] = (x[15]);
  assign t[282] = (x[15]);
  assign t[283] = (x[20]);
  assign t[284] = (x[20]);
  assign t[285] = (x[23]);
  assign t[286] = (x[23]);
  assign t[287] = (x[28]);
  assign t[288] = (x[28]);
  assign t[289] = (x[31]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[31]);
  assign t[291] = (x[36]);
  assign t[292] = (x[36]);
  assign t[293] = (x[39]);
  assign t[294] = (x[39]);
  assign t[295] = (x[42]);
  assign t[296] = (x[42]);
  assign t[297] = (x[45]);
  assign t[298] = (x[45]);
  assign t[299] = (x[48]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = (x[48]);
  assign t[301] = (x[53]);
  assign t[302] = (x[53]);
  assign t[303] = (x[56]);
  assign t[304] = (x[56]);
  assign t[305] = (x[61]);
  assign t[306] = (x[61]);
  assign t[307] = (x[64]);
  assign t[308] = (x[64]);
  assign t[309] = (x[67]);
  assign t[30] = t[16] ? x[27] : x[26];
  assign t[310] = (x[67]);
  assign t[311] = (x[70]);
  assign t[312] = (x[70]);
  assign t[313] = (x[73]);
  assign t[314] = (x[73]);
  assign t[315] = (x[78]);
  assign t[316] = (x[78]);
  assign t[317] = (x[81]);
  assign t[318] = (x[81]);
  assign t[319] = (x[86]);
  assign t[31] = ~(t[46] & t[47]);
  assign t[320] = (x[86]);
  assign t[321] = (x[89]);
  assign t[322] = (x[89]);
  assign t[323] = (x[92]);
  assign t[324] = (x[92]);
  assign t[325] = (x[95]);
  assign t[326] = (x[95]);
  assign t[327] = (x[98]);
  assign t[328] = (x[98]);
  assign t[329] = (x[101]);
  assign t[32] = ~(t[48] & t[49]);
  assign t[330] = (x[101]);
  assign t[331] = (x[104]);
  assign t[332] = (x[104]);
  assign t[333] = (x[107]);
  assign t[334] = (x[107]);
  assign t[335] = (x[110]);
  assign t[336] = (x[110]);
  assign t[337] = (x[113]);
  assign t[338] = (x[113]);
  assign t[339] = (x[116]);
  assign t[33] = t[50] ^ t[40];
  assign t[340] = (x[116]);
  assign t[341] = (x[119]);
  assign t[342] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[105] & t[54]);
  assign t[37] = ~(t[106] & t[55]);
  assign t[38] = t[16] ? x[35] : x[34];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[61];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[66]);
  assign t[46] = ~(t[108] & t[67]);
  assign t[47] = ~(t[109] & t[68]);
  assign t[48] = ~(t[110] & t[69]);
  assign t[49] = ~(t[111] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = t[71] ? x[52] : x[51];
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[71] ? x[60] : x[59];
  assign t[54] = ~(t[114]);
  assign t[55] = ~(t[114] & t[74]);
  assign t[56] = ~(t[115] & t[75]);
  assign t[57] = ~(t[116] & t[76]);
  assign t[58] = ~(t[117] & t[77]);
  assign t[59] = ~(t[118] & t[78]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = t[79] ? x[77] : x[76];
  assign t[61] = ~(t[80] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[79] ? x[85] : x[84];
  assign t[65] = ~(t[84] & t[85]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[121]);
  assign t[68] = ~(t[121] & t[86]);
  assign t[69] = ~(t[122]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[23]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[105]);
  assign t[75] = ~(t[124]);
  assign t[76] = ~(t[124] & t[89]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[23]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[115]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[131]);
  assign t[92] = ~(t[131] & t[96]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[126]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [151:0] x;
 output y;

 wire [432:0] t;
  assign t[0] = t[1] ? t[2] : t[118];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[144] & t[143]);
  assign t[103] = ~(t[154]);
  assign t[104] = ~(t[146] & t[145]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[114] & t[115]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = t[208] ^ x[2];
  assign t[164] = t[209] ^ x[8];
  assign t[165] = t[210] ^ x[11];
  assign t[166] = t[211] ^ x[14];
  assign t[167] = t[212] ^ x[17];
  assign t[168] = t[213] ^ x[22];
  assign t[169] = t[214] ^ x[27];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[32];
  assign t[171] = t[216] ^ x[35];
  assign t[172] = t[217] ^ x[38];
  assign t[173] = t[218] ^ x[41];
  assign t[174] = t[219] ^ x[46];
  assign t[175] = t[220] ^ x[51];
  assign t[176] = t[221] ^ x[54];
  assign t[177] = t[222] ^ x[57];
  assign t[178] = t[223] ^ x[60];
  assign t[179] = t[224] ^ x[65];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[70];
  assign t[181] = t[226] ^ x[73];
  assign t[182] = t[227] ^ x[76];
  assign t[183] = t[228] ^ x[79];
  assign t[184] = t[229] ^ x[82];
  assign t[185] = t[230] ^ x[85];
  assign t[186] = t[231] ^ x[88];
  assign t[187] = t[232] ^ x[91];
  assign t[188] = t[233] ^ x[94];
  assign t[189] = t[234] ^ x[97];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[100];
  assign t[191] = t[236] ^ x[103];
  assign t[192] = t[237] ^ x[106];
  assign t[193] = t[238] ^ x[109];
  assign t[194] = t[239] ^ x[112];
  assign t[195] = t[240] ^ x[115];
  assign t[196] = t[241] ^ x[118];
  assign t[197] = t[242] ^ x[121];
  assign t[198] = t[243] ^ x[124];
  assign t[199] = t[244] ^ x[127];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[130];
  assign t[201] = t[246] ^ x[133];
  assign t[202] = t[247] ^ x[136];
  assign t[203] = t[248] ^ x[139];
  assign t[204] = t[249] ^ x[142];
  assign t[205] = t[250] ^ x[145];
  assign t[206] = t[251] ^ x[148];
  assign t[207] = t[252] ^ x[151];
  assign t[208] = (t[253] & ~t[254]);
  assign t[209] = (t[255] & ~t[256]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[257] & ~t[258]);
  assign t[211] = (t[259] & ~t[260]);
  assign t[212] = (t[261] & ~t[262]);
  assign t[213] = (t[263] & ~t[264]);
  assign t[214] = (t[265] & ~t[266]);
  assign t[215] = (t[267] & ~t[268]);
  assign t[216] = (t[269] & ~t[270]);
  assign t[217] = (t[271] & ~t[272]);
  assign t[218] = (t[273] & ~t[274]);
  assign t[219] = (t[275] & ~t[276]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[277] & ~t[278]);
  assign t[221] = (t[279] & ~t[280]);
  assign t[222] = (t[281] & ~t[282]);
  assign t[223] = (t[283] & ~t[284]);
  assign t[224] = (t[285] & ~t[286]);
  assign t[225] = (t[287] & ~t[288]);
  assign t[226] = (t[289] & ~t[290]);
  assign t[227] = (t[291] & ~t[292]);
  assign t[228] = (t[293] & ~t[294]);
  assign t[229] = (t[295] & ~t[296]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[297] & ~t[298]);
  assign t[231] = (t[299] & ~t[300]);
  assign t[232] = (t[301] & ~t[302]);
  assign t[233] = (t[303] & ~t[304]);
  assign t[234] = (t[305] & ~t[306]);
  assign t[235] = (t[307] & ~t[308]);
  assign t[236] = (t[309] & ~t[310]);
  assign t[237] = (t[311] & ~t[312]);
  assign t[238] = (t[313] & ~t[314]);
  assign t[239] = (t[315] & ~t[316]);
  assign t[23] = ~(t[121]);
  assign t[240] = (t[317] & ~t[318]);
  assign t[241] = (t[319] & ~t[320]);
  assign t[242] = (t[321] & ~t[322]);
  assign t[243] = (t[323] & ~t[324]);
  assign t[244] = (t[325] & ~t[326]);
  assign t[245] = (t[327] & ~t[328]);
  assign t[246] = (t[329] & ~t[330]);
  assign t[247] = (t[331] & ~t[332]);
  assign t[248] = (t[333] & ~t[334]);
  assign t[249] = (t[335] & ~t[336]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (t[337] & ~t[338]);
  assign t[251] = (t[339] & ~t[340]);
  assign t[252] = (t[341] & ~t[342]);
  assign t[253] = t[343] ^ x[2];
  assign t[254] = t[344] ^ x[1];
  assign t[255] = t[345] ^ x[8];
  assign t[256] = t[346] ^ x[7];
  assign t[257] = t[347] ^ x[11];
  assign t[258] = t[348] ^ x[10];
  assign t[259] = t[349] ^ x[14];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[13];
  assign t[261] = t[351] ^ x[17];
  assign t[262] = t[352] ^ x[16];
  assign t[263] = t[353] ^ x[22];
  assign t[264] = t[354] ^ x[21];
  assign t[265] = t[355] ^ x[27];
  assign t[266] = t[356] ^ x[26];
  assign t[267] = t[357] ^ x[32];
  assign t[268] = t[358] ^ x[31];
  assign t[269] = t[359] ^ x[35];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[34];
  assign t[271] = t[361] ^ x[38];
  assign t[272] = t[362] ^ x[37];
  assign t[273] = t[363] ^ x[41];
  assign t[274] = t[364] ^ x[40];
  assign t[275] = t[365] ^ x[46];
  assign t[276] = t[366] ^ x[45];
  assign t[277] = t[367] ^ x[51];
  assign t[278] = t[368] ^ x[50];
  assign t[279] = t[369] ^ x[54];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[53];
  assign t[281] = t[371] ^ x[57];
  assign t[282] = t[372] ^ x[56];
  assign t[283] = t[373] ^ x[60];
  assign t[284] = t[374] ^ x[59];
  assign t[285] = t[375] ^ x[65];
  assign t[286] = t[376] ^ x[64];
  assign t[287] = t[377] ^ x[70];
  assign t[288] = t[378] ^ x[69];
  assign t[289] = t[379] ^ x[73];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[72];
  assign t[291] = t[381] ^ x[76];
  assign t[292] = t[382] ^ x[75];
  assign t[293] = t[383] ^ x[79];
  assign t[294] = t[384] ^ x[78];
  assign t[295] = t[385] ^ x[82];
  assign t[296] = t[386] ^ x[81];
  assign t[297] = t[387] ^ x[85];
  assign t[298] = t[388] ^ x[84];
  assign t[299] = t[389] ^ x[88];
  assign t[29] = ~(t[46] & t[123]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[87];
  assign t[301] = t[391] ^ x[91];
  assign t[302] = t[392] ^ x[90];
  assign t[303] = t[393] ^ x[94];
  assign t[304] = t[394] ^ x[93];
  assign t[305] = t[395] ^ x[97];
  assign t[306] = t[396] ^ x[96];
  assign t[307] = t[397] ^ x[100];
  assign t[308] = t[398] ^ x[99];
  assign t[309] = t[399] ^ x[103];
  assign t[30] = t[16] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[102];
  assign t[311] = t[401] ^ x[106];
  assign t[312] = t[402] ^ x[105];
  assign t[313] = t[403] ^ x[109];
  assign t[314] = t[404] ^ x[108];
  assign t[315] = t[405] ^ x[112];
  assign t[316] = t[406] ^ x[111];
  assign t[317] = t[407] ^ x[115];
  assign t[318] = t[408] ^ x[114];
  assign t[319] = t[409] ^ x[118];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[410] ^ x[117];
  assign t[321] = t[411] ^ x[121];
  assign t[322] = t[412] ^ x[120];
  assign t[323] = t[413] ^ x[124];
  assign t[324] = t[414] ^ x[123];
  assign t[325] = t[415] ^ x[127];
  assign t[326] = t[416] ^ x[126];
  assign t[327] = t[417] ^ x[130];
  assign t[328] = t[418] ^ x[129];
  assign t[329] = t[419] ^ x[133];
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = t[420] ^ x[132];
  assign t[331] = t[421] ^ x[136];
  assign t[332] = t[422] ^ x[135];
  assign t[333] = t[423] ^ x[139];
  assign t[334] = t[424] ^ x[138];
  assign t[335] = t[425] ^ x[142];
  assign t[336] = t[426] ^ x[141];
  assign t[337] = t[427] ^ x[145];
  assign t[338] = t[428] ^ x[144];
  assign t[339] = t[429] ^ x[148];
  assign t[33] = t[51] ^ t[32];
  assign t[340] = t[430] ^ x[147];
  assign t[341] = t[431] ^ x[151];
  assign t[342] = t[432] ^ x[150];
  assign t[343] = (x[0]);
  assign t[344] = (x[0]);
  assign t[345] = (x[6]);
  assign t[346] = (x[6]);
  assign t[347] = (x[9]);
  assign t[348] = (x[9]);
  assign t[349] = (x[12]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[12]);
  assign t[351] = (x[15]);
  assign t[352] = (x[15]);
  assign t[353] = (x[20]);
  assign t[354] = (x[20]);
  assign t[355] = (x[25]);
  assign t[356] = (x[25]);
  assign t[357] = (x[30]);
  assign t[358] = (x[30]);
  assign t[359] = (x[33]);
  assign t[35] = t[54] ^ t[40];
  assign t[360] = (x[33]);
  assign t[361] = (x[36]);
  assign t[362] = (x[36]);
  assign t[363] = (x[39]);
  assign t[364] = (x[39]);
  assign t[365] = (x[44]);
  assign t[366] = (x[44]);
  assign t[367] = (x[49]);
  assign t[368] = (x[49]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[370] = (x[52]);
  assign t[371] = (x[55]);
  assign t[372] = (x[55]);
  assign t[373] = (x[58]);
  assign t[374] = (x[58]);
  assign t[375] = (x[63]);
  assign t[376] = (x[63]);
  assign t[377] = (x[68]);
  assign t[378] = (x[68]);
  assign t[379] = (x[71]);
  assign t[37] = ~(t[57] & t[124]);
  assign t[380] = (x[71]);
  assign t[381] = (x[74]);
  assign t[382] = (x[74]);
  assign t[383] = (x[77]);
  assign t[384] = (x[77]);
  assign t[385] = (x[80]);
  assign t[386] = (x[80]);
  assign t[387] = (x[83]);
  assign t[388] = (x[83]);
  assign t[389] = (x[86]);
  assign t[38] = t[16] ? x[29] : x[28];
  assign t[390] = (x[86]);
  assign t[391] = (x[89]);
  assign t[392] = (x[89]);
  assign t[393] = (x[92]);
  assign t[394] = (x[92]);
  assign t[395] = (x[95]);
  assign t[396] = (x[95]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[399] = (x[101]);
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[101]);
  assign t[401] = (x[104]);
  assign t[402] = (x[104]);
  assign t[403] = (x[107]);
  assign t[404] = (x[107]);
  assign t[405] = (x[110]);
  assign t[406] = (x[110]);
  assign t[407] = (x[113]);
  assign t[408] = (x[113]);
  assign t[409] = (x[116]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[410] = (x[116]);
  assign t[411] = (x[119]);
  assign t[412] = (x[119]);
  assign t[413] = (x[122]);
  assign t[414] = (x[122]);
  assign t[415] = (x[125]);
  assign t[416] = (x[125]);
  assign t[417] = (x[128]);
  assign t[418] = (x[128]);
  assign t[419] = (x[131]);
  assign t[41] = t[62] ^ t[63];
  assign t[420] = (x[131]);
  assign t[421] = (x[134]);
  assign t[422] = (x[134]);
  assign t[423] = (x[137]);
  assign t[424] = (x[137]);
  assign t[425] = (x[140]);
  assign t[426] = (x[140]);
  assign t[427] = (x[143]);
  assign t[428] = (x[143]);
  assign t[429] = (x[146]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[149]);
  assign t[432] = (x[149]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[125]);
  assign t[45] = ~(t[126]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[127]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = t[76] ? x[43] : x[42];
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[129]);
  assign t[54] = t[76] ? x[48] : x[47];
  assign t[55] = ~(t[130]);
  assign t[56] = ~(t[131]);
  assign t[57] = ~(t[80] & t[81]);
  assign t[58] = ~(t[82] & t[83]);
  assign t[59] = ~(t[84] & t[132]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[85] & t[86]);
  assign t[61] = ~(t[87] & t[133]);
  assign t[62] = t[88] ? x[62] : x[61];
  assign t[63] = ~(t[89] & t[90]);
  assign t[64] = ~(t[91] & t[92]);
  assign t[65] = ~(t[93] & t[134]);
  assign t[66] = t[88] ? x[67] : x[66];
  assign t[67] = ~(t[94] & t[95]);
  assign t[68] = ~(t[126] & t[125]);
  assign t[69] = ~(t[135]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[136]);
  assign t[71] = ~(t[137]);
  assign t[72] = ~(t[96] & t[97]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[139]);
  assign t[75] = ~(t[98] & t[99]);
  assign t[76] = ~(t[23]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[119] & t[120]);
  assign t[80] = ~(t[131] & t[130]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[102] & t[103]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[104] & t[105]);
  assign t[88] = ~(t[23]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[121] & t[122]);
  assign t[90] = ~(t[108] & t[147]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[109] & t[110]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [151:0] x;
 output y;

 wire [432:0] t;
  assign t[0] = t[1] ? t[2] : t[118];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[144] & t[143]);
  assign t[103] = ~(t[154]);
  assign t[104] = ~(t[146] & t[145]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[114] & t[115]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[18] ^ x[19];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[19] : x[18];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = t[208] ^ x[2];
  assign t[164] = t[209] ^ x[8];
  assign t[165] = t[210] ^ x[11];
  assign t[166] = t[211] ^ x[14];
  assign t[167] = t[212] ^ x[17];
  assign t[168] = t[213] ^ x[22];
  assign t[169] = t[214] ^ x[27];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[32];
  assign t[171] = t[216] ^ x[35];
  assign t[172] = t[217] ^ x[38];
  assign t[173] = t[218] ^ x[41];
  assign t[174] = t[219] ^ x[46];
  assign t[175] = t[220] ^ x[51];
  assign t[176] = t[221] ^ x[54];
  assign t[177] = t[222] ^ x[57];
  assign t[178] = t[223] ^ x[60];
  assign t[179] = t[224] ^ x[65];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[70];
  assign t[181] = t[226] ^ x[73];
  assign t[182] = t[227] ^ x[76];
  assign t[183] = t[228] ^ x[79];
  assign t[184] = t[229] ^ x[82];
  assign t[185] = t[230] ^ x[85];
  assign t[186] = t[231] ^ x[88];
  assign t[187] = t[232] ^ x[91];
  assign t[188] = t[233] ^ x[94];
  assign t[189] = t[234] ^ x[97];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[100];
  assign t[191] = t[236] ^ x[103];
  assign t[192] = t[237] ^ x[106];
  assign t[193] = t[238] ^ x[109];
  assign t[194] = t[239] ^ x[112];
  assign t[195] = t[240] ^ x[115];
  assign t[196] = t[241] ^ x[118];
  assign t[197] = t[242] ^ x[121];
  assign t[198] = t[243] ^ x[124];
  assign t[199] = t[244] ^ x[127];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[130];
  assign t[201] = t[246] ^ x[133];
  assign t[202] = t[247] ^ x[136];
  assign t[203] = t[248] ^ x[139];
  assign t[204] = t[249] ^ x[142];
  assign t[205] = t[250] ^ x[145];
  assign t[206] = t[251] ^ x[148];
  assign t[207] = t[252] ^ x[151];
  assign t[208] = (t[253] & ~t[254]);
  assign t[209] = (t[255] & ~t[256]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (t[257] & ~t[258]);
  assign t[211] = (t[259] & ~t[260]);
  assign t[212] = (t[261] & ~t[262]);
  assign t[213] = (t[263] & ~t[264]);
  assign t[214] = (t[265] & ~t[266]);
  assign t[215] = (t[267] & ~t[268]);
  assign t[216] = (t[269] & ~t[270]);
  assign t[217] = (t[271] & ~t[272]);
  assign t[218] = (t[273] & ~t[274]);
  assign t[219] = (t[275] & ~t[276]);
  assign t[21] = x[4] ? t[33] : t[32];
  assign t[220] = (t[277] & ~t[278]);
  assign t[221] = (t[279] & ~t[280]);
  assign t[222] = (t[281] & ~t[282]);
  assign t[223] = (t[283] & ~t[284]);
  assign t[224] = (t[285] & ~t[286]);
  assign t[225] = (t[287] & ~t[288]);
  assign t[226] = (t[289] & ~t[290]);
  assign t[227] = (t[291] & ~t[292]);
  assign t[228] = (t[293] & ~t[294]);
  assign t[229] = (t[295] & ~t[296]);
  assign t[22] = x[4] ? t[35] : t[34];
  assign t[230] = (t[297] & ~t[298]);
  assign t[231] = (t[299] & ~t[300]);
  assign t[232] = (t[301] & ~t[302]);
  assign t[233] = (t[303] & ~t[304]);
  assign t[234] = (t[305] & ~t[306]);
  assign t[235] = (t[307] & ~t[308]);
  assign t[236] = (t[309] & ~t[310]);
  assign t[237] = (t[311] & ~t[312]);
  assign t[238] = (t[313] & ~t[314]);
  assign t[239] = (t[315] & ~t[316]);
  assign t[23] = ~(t[121]);
  assign t[240] = (t[317] & ~t[318]);
  assign t[241] = (t[319] & ~t[320]);
  assign t[242] = (t[321] & ~t[322]);
  assign t[243] = (t[323] & ~t[324]);
  assign t[244] = (t[325] & ~t[326]);
  assign t[245] = (t[327] & ~t[328]);
  assign t[246] = (t[329] & ~t[330]);
  assign t[247] = (t[331] & ~t[332]);
  assign t[248] = (t[333] & ~t[334]);
  assign t[249] = (t[335] & ~t[336]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (t[337] & ~t[338]);
  assign t[251] = (t[339] & ~t[340]);
  assign t[252] = (t[341] & ~t[342]);
  assign t[253] = t[343] ^ x[2];
  assign t[254] = t[344] ^ x[1];
  assign t[255] = t[345] ^ x[8];
  assign t[256] = t[346] ^ x[7];
  assign t[257] = t[347] ^ x[11];
  assign t[258] = t[348] ^ x[10];
  assign t[259] = t[349] ^ x[14];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[350] ^ x[13];
  assign t[261] = t[351] ^ x[17];
  assign t[262] = t[352] ^ x[16];
  assign t[263] = t[353] ^ x[22];
  assign t[264] = t[354] ^ x[21];
  assign t[265] = t[355] ^ x[27];
  assign t[266] = t[356] ^ x[26];
  assign t[267] = t[357] ^ x[32];
  assign t[268] = t[358] ^ x[31];
  assign t[269] = t[359] ^ x[35];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[270] = t[360] ^ x[34];
  assign t[271] = t[361] ^ x[38];
  assign t[272] = t[362] ^ x[37];
  assign t[273] = t[363] ^ x[41];
  assign t[274] = t[364] ^ x[40];
  assign t[275] = t[365] ^ x[46];
  assign t[276] = t[366] ^ x[45];
  assign t[277] = t[367] ^ x[51];
  assign t[278] = t[368] ^ x[50];
  assign t[279] = t[369] ^ x[54];
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = t[370] ^ x[53];
  assign t[281] = t[371] ^ x[57];
  assign t[282] = t[372] ^ x[56];
  assign t[283] = t[373] ^ x[60];
  assign t[284] = t[374] ^ x[59];
  assign t[285] = t[375] ^ x[65];
  assign t[286] = t[376] ^ x[64];
  assign t[287] = t[377] ^ x[70];
  assign t[288] = t[378] ^ x[69];
  assign t[289] = t[379] ^ x[73];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[380] ^ x[72];
  assign t[291] = t[381] ^ x[76];
  assign t[292] = t[382] ^ x[75];
  assign t[293] = t[383] ^ x[79];
  assign t[294] = t[384] ^ x[78];
  assign t[295] = t[385] ^ x[82];
  assign t[296] = t[386] ^ x[81];
  assign t[297] = t[387] ^ x[85];
  assign t[298] = t[388] ^ x[84];
  assign t[299] = t[389] ^ x[88];
  assign t[29] = ~(t[46] & t[123]);
  assign t[2] = x[3] ? t[6] : t[5];
  assign t[300] = t[390] ^ x[87];
  assign t[301] = t[391] ^ x[91];
  assign t[302] = t[392] ^ x[90];
  assign t[303] = t[393] ^ x[94];
  assign t[304] = t[394] ^ x[93];
  assign t[305] = t[395] ^ x[97];
  assign t[306] = t[396] ^ x[96];
  assign t[307] = t[397] ^ x[100];
  assign t[308] = t[398] ^ x[99];
  assign t[309] = t[399] ^ x[103];
  assign t[30] = t[16] ? x[24] : x[23];
  assign t[310] = t[400] ^ x[102];
  assign t[311] = t[401] ^ x[106];
  assign t[312] = t[402] ^ x[105];
  assign t[313] = t[403] ^ x[109];
  assign t[314] = t[404] ^ x[108];
  assign t[315] = t[405] ^ x[112];
  assign t[316] = t[406] ^ x[111];
  assign t[317] = t[407] ^ x[115];
  assign t[318] = t[408] ^ x[114];
  assign t[319] = t[409] ^ x[118];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[410] ^ x[117];
  assign t[321] = t[411] ^ x[121];
  assign t[322] = t[412] ^ x[120];
  assign t[323] = t[413] ^ x[124];
  assign t[324] = t[414] ^ x[123];
  assign t[325] = t[415] ^ x[127];
  assign t[326] = t[416] ^ x[126];
  assign t[327] = t[417] ^ x[130];
  assign t[328] = t[418] ^ x[129];
  assign t[329] = t[419] ^ x[133];
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = t[420] ^ x[132];
  assign t[331] = t[421] ^ x[136];
  assign t[332] = t[422] ^ x[135];
  assign t[333] = t[423] ^ x[139];
  assign t[334] = t[424] ^ x[138];
  assign t[335] = t[425] ^ x[142];
  assign t[336] = t[426] ^ x[141];
  assign t[337] = t[427] ^ x[145];
  assign t[338] = t[428] ^ x[144];
  assign t[339] = t[429] ^ x[148];
  assign t[33] = t[51] ^ t[32];
  assign t[340] = t[430] ^ x[147];
  assign t[341] = t[431] ^ x[151];
  assign t[342] = t[432] ^ x[150];
  assign t[343] = (x[0]);
  assign t[344] = (x[0]);
  assign t[345] = (x[6]);
  assign t[346] = (x[6]);
  assign t[347] = (x[9]);
  assign t[348] = (x[9]);
  assign t[349] = (x[12]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[12]);
  assign t[351] = (x[15]);
  assign t[352] = (x[15]);
  assign t[353] = (x[20]);
  assign t[354] = (x[20]);
  assign t[355] = (x[25]);
  assign t[356] = (x[25]);
  assign t[357] = (x[30]);
  assign t[358] = (x[30]);
  assign t[359] = (x[33]);
  assign t[35] = t[54] ^ t[40];
  assign t[360] = (x[33]);
  assign t[361] = (x[36]);
  assign t[362] = (x[36]);
  assign t[363] = (x[39]);
  assign t[364] = (x[39]);
  assign t[365] = (x[44]);
  assign t[366] = (x[44]);
  assign t[367] = (x[49]);
  assign t[368] = (x[49]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[370] = (x[52]);
  assign t[371] = (x[55]);
  assign t[372] = (x[55]);
  assign t[373] = (x[58]);
  assign t[374] = (x[58]);
  assign t[375] = (x[63]);
  assign t[376] = (x[63]);
  assign t[377] = (x[68]);
  assign t[378] = (x[68]);
  assign t[379] = (x[71]);
  assign t[37] = ~(t[57] & t[124]);
  assign t[380] = (x[71]);
  assign t[381] = (x[74]);
  assign t[382] = (x[74]);
  assign t[383] = (x[77]);
  assign t[384] = (x[77]);
  assign t[385] = (x[80]);
  assign t[386] = (x[80]);
  assign t[387] = (x[83]);
  assign t[388] = (x[83]);
  assign t[389] = (x[86]);
  assign t[38] = t[16] ? x[29] : x[28];
  assign t[390] = (x[86]);
  assign t[391] = (x[89]);
  assign t[392] = (x[89]);
  assign t[393] = (x[92]);
  assign t[394] = (x[92]);
  assign t[395] = (x[95]);
  assign t[396] = (x[95]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[399] = (x[101]);
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[101]);
  assign t[401] = (x[104]);
  assign t[402] = (x[104]);
  assign t[403] = (x[107]);
  assign t[404] = (x[107]);
  assign t[405] = (x[110]);
  assign t[406] = (x[110]);
  assign t[407] = (x[113]);
  assign t[408] = (x[113]);
  assign t[409] = (x[116]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[410] = (x[116]);
  assign t[411] = (x[119]);
  assign t[412] = (x[119]);
  assign t[413] = (x[122]);
  assign t[414] = (x[122]);
  assign t[415] = (x[125]);
  assign t[416] = (x[125]);
  assign t[417] = (x[128]);
  assign t[418] = (x[128]);
  assign t[419] = (x[131]);
  assign t[41] = t[62] ^ t[63];
  assign t[420] = (x[131]);
  assign t[421] = (x[134]);
  assign t[422] = (x[134]);
  assign t[423] = (x[137]);
  assign t[424] = (x[137]);
  assign t[425] = (x[140]);
  assign t[426] = (x[140]);
  assign t[427] = (x[143]);
  assign t[428] = (x[143]);
  assign t[429] = (x[146]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[430] = (x[146]);
  assign t[431] = (x[149]);
  assign t[432] = (x[149]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[125]);
  assign t[45] = ~(t[126]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[127]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = ~(x[3]);
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = t[76] ? x[43] : x[42];
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[129]);
  assign t[54] = t[76] ? x[48] : x[47];
  assign t[55] = ~(t[130]);
  assign t[56] = ~(t[131]);
  assign t[57] = ~(t[80] & t[81]);
  assign t[58] = ~(t[82] & t[83]);
  assign t[59] = ~(t[84] & t[132]);
  assign t[5] = x[4] ? t[10] : t[9];
  assign t[60] = ~(t[85] & t[86]);
  assign t[61] = ~(t[87] & t[133]);
  assign t[62] = t[88] ? x[62] : x[61];
  assign t[63] = ~(t[89] & t[90]);
  assign t[64] = ~(t[91] & t[92]);
  assign t[65] = ~(t[93] & t[134]);
  assign t[66] = t[88] ? x[67] : x[66];
  assign t[67] = ~(t[94] & t[95]);
  assign t[68] = ~(t[126] & t[125]);
  assign t[69] = ~(t[135]);
  assign t[6] = t[11] ^ x[5];
  assign t[70] = ~(t[136]);
  assign t[71] = ~(t[137]);
  assign t[72] = ~(t[96] & t[97]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[139]);
  assign t[75] = ~(t[98] & t[99]);
  assign t[76] = ~(t[23]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[119] & t[120]);
  assign t[80] = ~(t[131] & t[130]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[102] & t[103]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[104] & t[105]);
  assign t[88] = ~(t[23]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[121] & t[122]);
  assign t[90] = ~(t[108] & t[147]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[109] & t[110]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind226(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[53] ^ t[34];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[56] ^ t[42];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[59] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[70] | t[46]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[73] | t[119];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[120];
  assign t[53] = t[77] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = t[80] | t[121];
  assign t[56] = t[77] ? x[48] : x[47];
  assign t[57] = ~(t[122]);
  assign t[58] = ~(t[123]);
  assign t[59] = ~(t[81] | t[57]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = t[84] | t[124];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[125];
  assign t[64] = t[88] ? x[62] : x[61];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = t[93] | t[126];
  assign t[68] = t[88] ? x[67] : x[66];
  assign t[69] = ~(t[94] & t[95]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[129]);
  assign t[73] = ~(t[96] | t[71]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[97] | t[74]);
  assign t[77] = ~(t[25]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[25]);
  assign t[89] = ~(t[101] & t[102]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = t[103] | t[139];
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[18] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[53] ^ t[34];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[56] ^ t[42];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[59] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[70] | t[46]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[73] | t[119];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[120];
  assign t[53] = t[77] ? x[43] : x[42];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = t[80] | t[121];
  assign t[56] = t[77] ? x[48] : x[47];
  assign t[57] = ~(t[122]);
  assign t[58] = ~(t[123]);
  assign t[59] = ~(t[81] | t[57]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = t[84] | t[124];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[125];
  assign t[64] = t[88] ? x[62] : x[61];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = t[93] | t[126];
  assign t[68] = t[88] ? x[67] : x[66];
  assign t[69] = ~(t[94] & t[95]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[129]);
  assign t[73] = ~(t[96] | t[71]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[97] | t[74]);
  assign t[77] = ~(t[25]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[25]);
  assign t[89] = ~(t[101] & t[102]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = t[103] | t[139];
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [106:0] x;
 output y;

 wire [375:0] t;
  assign t[0] = t[1] ? t[2] : t[152];
  assign t[100] = ~(t[176]);
  assign t[101] = ~(t[177]);
  assign t[102] = ~(t[120] | t[121]);
  assign t[103] = ~(t[40]);
  assign t[104] = ~(t[122] | t[123]);
  assign t[105] = ~(t[124] & t[125]);
  assign t[106] = ~(t[178]);
  assign t[107] = ~(t[170] | t[171]);
  assign t[108] = ~(t[179]);
  assign t[109] = ~(t[180]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[126] | t[127]);
  assign t[111] = ~(t[114] | t[128]);
  assign t[112] = ~(t[181]);
  assign t[113] = ~(t[173] | t[174]);
  assign t[114] = ~(t[43] | t[129]);
  assign t[115] = ~(t[130]);
  assign t[116] = ~(t[131] & t[95]);
  assign t[117] = ~(t[132] & t[95]);
  assign t[118] = ~(t[97] & t[95]);
  assign t[119] = ~(t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[182]);
  assign t[121] = ~(t[176] | t[177]);
  assign t[122] = ~(t[133] & t[42]);
  assign t[123] = t[29] | t[134];
  assign t[124] = t[156] & t[135];
  assign t[125] = t[131] | t[132];
  assign t[126] = ~(t[183]);
  assign t[127] = ~(t[179] | t[180]);
  assign t[128] = ~(t[136] & t[137]);
  assign t[129] = t[153] ? t[138] : t[116];
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[139] | t[140]);
  assign t[131] = ~(x[4] | t[154]);
  assign t[132] = x[4] & t[154];
  assign t[133] = ~(t[135] & t[141]);
  assign t[134] = ~(t[43] | t[142]);
  assign t[135] = ~(t[67] | t[153]);
  assign t[136] = ~(t[143] | t[144]);
  assign t[137] = ~(t[67] & t[145]);
  assign t[138] = ~(t[132] & t[156]);
  assign t[139] = ~(t[43] | t[146]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(t[43] | t[147]);
  assign t[141] = ~(t[69] & t[148]);
  assign t[142] = t[153] ? t[149] : t[117];
  assign t[143] = ~(t[67] | t[150]);
  assign t[144] = ~(t[43] | t[151]);
  assign t[145] = ~(t[68] & t[69]);
  assign t[146] = t[153] ? t[148] : t[118];
  assign t[147] = t[153] ? t[117] : t[149];
  assign t[148] = ~(x[4] & t[65]);
  assign t[149] = ~(t[131] & t[156]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[153] ? t[116] : t[117];
  assign t[151] = t[153] ? t[118] : t[148];
  assign t[152] = (t[184]);
  assign t[153] = (t[185]);
  assign t[154] = (t[186]);
  assign t[155] = (t[187]);
  assign t[156] = (t[188]);
  assign t[157] = (t[189]);
  assign t[158] = (t[190]);
  assign t[159] = (t[191]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[192]);
  assign t[161] = (t[193]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[153] & t[154]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[155] & t[156]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = t[216] ^ x[2];
  assign t[185] = t[217] ^ x[10];
  assign t[186] = t[218] ^ x[13];
  assign t[187] = t[219] ^ x[16];
  assign t[188] = t[220] ^ x[19];
  assign t[189] = t[221] ^ x[22];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[222] ^ x[25];
  assign t[191] = t[223] ^ x[28];
  assign t[192] = t[224] ^ x[31];
  assign t[193] = t[225] ^ x[34];
  assign t[194] = t[226] ^ x[37];
  assign t[195] = t[227] ^ x[40];
  assign t[196] = t[228] ^ x[43];
  assign t[197] = t[229] ^ x[46];
  assign t[198] = t[230] ^ x[51];
  assign t[199] = t[231] ^ x[54];
  assign t[19] = t[27] ? x[7] : x[6];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[57];
  assign t[201] = t[233] ^ x[60];
  assign t[202] = t[234] ^ x[65];
  assign t[203] = t[235] ^ x[68];
  assign t[204] = t[236] ^ x[71];
  assign t[205] = t[237] ^ x[76];
  assign t[206] = t[238] ^ x[79];
  assign t[207] = t[239] ^ x[82];
  assign t[208] = t[240] ^ x[85];
  assign t[209] = t[241] ^ x[88];
  assign t[20] = t[28] | t[29];
  assign t[210] = t[242] ^ x[91];
  assign t[211] = t[243] ^ x[94];
  assign t[212] = t[244] ^ x[97];
  assign t[213] = t[245] ^ x[100];
  assign t[214] = t[246] ^ x[103];
  assign t[215] = t[247] ^ x[106];
  assign t[216] = (t[248] & ~t[249]);
  assign t[217] = (t[250] & ~t[251]);
  assign t[218] = (t[252] & ~t[253]);
  assign t[219] = (t[254] & ~t[255]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = (t[256] & ~t[257]);
  assign t[221] = (t[258] & ~t[259]);
  assign t[222] = (t[260] & ~t[261]);
  assign t[223] = (t[262] & ~t[263]);
  assign t[224] = (t[264] & ~t[265]);
  assign t[225] = (t[266] & ~t[267]);
  assign t[226] = (t[268] & ~t[269]);
  assign t[227] = (t[270] & ~t[271]);
  assign t[228] = (t[272] & ~t[273]);
  assign t[229] = (t[274] & ~t[275]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (t[276] & ~t[277]);
  assign t[231] = (t[278] & ~t[279]);
  assign t[232] = (t[280] & ~t[281]);
  assign t[233] = (t[282] & ~t[283]);
  assign t[234] = (t[284] & ~t[285]);
  assign t[235] = (t[286] & ~t[287]);
  assign t[236] = (t[288] & ~t[289]);
  assign t[237] = (t[290] & ~t[291]);
  assign t[238] = (t[292] & ~t[293]);
  assign t[239] = (t[294] & ~t[295]);
  assign t[23] = x[4] ? t[33] : t[32];
  assign t[240] = (t[296] & ~t[297]);
  assign t[241] = (t[298] & ~t[299]);
  assign t[242] = (t[300] & ~t[301]);
  assign t[243] = (t[302] & ~t[303]);
  assign t[244] = (t[304] & ~t[305]);
  assign t[245] = (t[306] & ~t[307]);
  assign t[246] = (t[308] & ~t[309]);
  assign t[247] = (t[310] & ~t[311]);
  assign t[248] = t[312] ^ x[2];
  assign t[249] = t[313] ^ x[1];
  assign t[24] = x[4] ? t[35] : t[34];
  assign t[250] = t[314] ^ x[10];
  assign t[251] = t[315] ^ x[9];
  assign t[252] = t[316] ^ x[13];
  assign t[253] = t[317] ^ x[12];
  assign t[254] = t[318] ^ x[16];
  assign t[255] = t[319] ^ x[15];
  assign t[256] = t[320] ^ x[19];
  assign t[257] = t[321] ^ x[18];
  assign t[258] = t[322] ^ x[22];
  assign t[259] = t[323] ^ x[21];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[324] ^ x[25];
  assign t[261] = t[325] ^ x[24];
  assign t[262] = t[326] ^ x[28];
  assign t[263] = t[327] ^ x[27];
  assign t[264] = t[328] ^ x[31];
  assign t[265] = t[329] ^ x[30];
  assign t[266] = t[330] ^ x[34];
  assign t[267] = t[331] ^ x[33];
  assign t[268] = t[332] ^ x[37];
  assign t[269] = t[333] ^ x[36];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[334] ^ x[40];
  assign t[271] = t[335] ^ x[39];
  assign t[272] = t[336] ^ x[43];
  assign t[273] = t[337] ^ x[42];
  assign t[274] = t[338] ^ x[46];
  assign t[275] = t[339] ^ x[45];
  assign t[276] = t[340] ^ x[51];
  assign t[277] = t[341] ^ x[50];
  assign t[278] = t[342] ^ x[54];
  assign t[279] = t[343] ^ x[53];
  assign t[27] = ~(t[40]);
  assign t[280] = t[344] ^ x[57];
  assign t[281] = t[345] ^ x[56];
  assign t[282] = t[346] ^ x[60];
  assign t[283] = t[347] ^ x[59];
  assign t[284] = t[348] ^ x[65];
  assign t[285] = t[349] ^ x[64];
  assign t[286] = t[350] ^ x[68];
  assign t[287] = t[351] ^ x[67];
  assign t[288] = t[352] ^ x[71];
  assign t[289] = t[353] ^ x[70];
  assign t[28] = ~(t[41] & t[42]);
  assign t[290] = t[354] ^ x[76];
  assign t[291] = t[355] ^ x[75];
  assign t[292] = t[356] ^ x[79];
  assign t[293] = t[357] ^ x[78];
  assign t[294] = t[358] ^ x[82];
  assign t[295] = t[359] ^ x[81];
  assign t[296] = t[360] ^ x[85];
  assign t[297] = t[361] ^ x[84];
  assign t[298] = t[362] ^ x[88];
  assign t[299] = t[363] ^ x[87];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[364] ^ x[91];
  assign t[301] = t[365] ^ x[90];
  assign t[302] = t[366] ^ x[94];
  assign t[303] = t[367] ^ x[93];
  assign t[304] = t[368] ^ x[97];
  assign t[305] = t[369] ^ x[96];
  assign t[306] = t[370] ^ x[100];
  assign t[307] = t[371] ^ x[99];
  assign t[308] = t[372] ^ x[103];
  assign t[309] = t[373] ^ x[102];
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = t[374] ^ x[106];
  assign t[311] = t[375] ^ x[105];
  assign t[312] = (x[0]);
  assign t[313] = (x[0]);
  assign t[314] = (x[8]);
  assign t[315] = (x[8]);
  assign t[316] = (x[11]);
  assign t[317] = (x[11]);
  assign t[318] = (x[14]);
  assign t[319] = (x[14]);
  assign t[31] = ~(t[157] | t[47]);
  assign t[320] = (x[17]);
  assign t[321] = (x[17]);
  assign t[322] = (x[20]);
  assign t[323] = (x[20]);
  assign t[324] = (x[23]);
  assign t[325] = (x[23]);
  assign t[326] = (x[26]);
  assign t[327] = (x[26]);
  assign t[328] = (x[29]);
  assign t[329] = (x[29]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[32]);
  assign t[331] = (x[32]);
  assign t[332] = (x[35]);
  assign t[333] = (x[35]);
  assign t[334] = (x[38]);
  assign t[335] = (x[38]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[44]);
  assign t[339] = (x[44]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[58]);
  assign t[347] = (x[58]);
  assign t[348] = (x[63]);
  assign t[349] = (x[63]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = (x[66]);
  assign t[351] = (x[66]);
  assign t[352] = (x[69]);
  assign t[353] = (x[69]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[37] = ~(t[158] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[155]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = ~(t[67]);
  assign t[44] = t[153] ? t[69] : t[68];
  assign t[45] = ~(t[159]);
  assign t[46] = ~(t[160]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[161] | t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[162] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[163]);
  assign t[57] = ~(t[164]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[165] | t[90]);
  assign t[61] = t[27] ? x[48] : x[47];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[67] | t[93]);
  assign t[64] = ~(t[67] | t[94]);
  assign t[65] = ~(t[154] | t[95]);
  assign t[66] = t[43] & t[153];
  assign t[67] = ~(t[155]);
  assign t[68] = ~(x[4] & t[96]);
  assign t[69] = ~(t[156] & t[97]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[166]);
  assign t[71] = ~(t[159] | t[160]);
  assign t[72] = ~(t[167]);
  assign t[73] = ~(t[168]);
  assign t[74] = ~(t[98] | t[99]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[169] | t[102]);
  assign t[77] = t[103] ? x[62] : x[61];
  assign t[78] = ~(t[104] & t[105]);
  assign t[79] = ~(t[170]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[171]);
  assign t[81] = ~(t[106] | t[107]);
  assign t[82] = ~(t[108] | t[109]);
  assign t[83] = ~(t[172] | t[110]);
  assign t[84] = t[103] ? x[73] : x[72];
  assign t[85] = ~(t[111] & t[42]);
  assign t[86] = ~(t[152]);
  assign t[87] = ~(t[163] | t[164]);
  assign t[88] = ~(t[173]);
  assign t[89] = ~(t[174]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112] | t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = ~(t[115] | t[29]);
  assign t[93] = t[153] ? t[117] : t[116];
  assign t[94] = t[153] ? t[118] : t[68];
  assign t[95] = ~(t[156]);
  assign t[96] = ~(t[154] | t[156]);
  assign t[97] = ~(x[4] | t[119]);
  assign t[98] = ~(t[175]);
  assign t[99] = ~(t[167] | t[168]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [106:0] x;
 output y;

 wire [375:0] t;
  assign t[0] = t[1] ? t[2] : t[152];
  assign t[100] = ~(t[176]);
  assign t[101] = ~(t[177]);
  assign t[102] = ~(t[120] | t[121]);
  assign t[103] = ~(t[40]);
  assign t[104] = ~(t[122] | t[123]);
  assign t[105] = ~(t[124] & t[125]);
  assign t[106] = ~(t[178]);
  assign t[107] = ~(t[170] | t[171]);
  assign t[108] = ~(t[179]);
  assign t[109] = ~(t[180]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[126] | t[127]);
  assign t[111] = ~(t[114] | t[128]);
  assign t[112] = ~(t[181]);
  assign t[113] = ~(t[173] | t[174]);
  assign t[114] = ~(t[43] | t[129]);
  assign t[115] = ~(t[130]);
  assign t[116] = ~(t[131] & t[95]);
  assign t[117] = ~(t[132] & t[95]);
  assign t[118] = ~(t[97] & t[95]);
  assign t[119] = ~(t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[182]);
  assign t[121] = ~(t[176] | t[177]);
  assign t[122] = ~(t[133] & t[42]);
  assign t[123] = t[29] | t[134];
  assign t[124] = t[156] & t[135];
  assign t[125] = t[131] | t[132];
  assign t[126] = ~(t[183]);
  assign t[127] = ~(t[179] | t[180]);
  assign t[128] = ~(t[136] & t[137]);
  assign t[129] = t[153] ? t[138] : t[116];
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[139] | t[140]);
  assign t[131] = ~(x[4] | t[154]);
  assign t[132] = x[4] & t[154];
  assign t[133] = ~(t[135] & t[141]);
  assign t[134] = ~(t[43] | t[142]);
  assign t[135] = ~(t[67] | t[153]);
  assign t[136] = ~(t[143] | t[144]);
  assign t[137] = ~(t[67] & t[145]);
  assign t[138] = ~(t[132] & t[156]);
  assign t[139] = ~(t[43] | t[146]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(t[43] | t[147]);
  assign t[141] = ~(t[69] & t[148]);
  assign t[142] = t[153] ? t[149] : t[117];
  assign t[143] = ~(t[67] | t[150]);
  assign t[144] = ~(t[43] | t[151]);
  assign t[145] = ~(t[68] & t[69]);
  assign t[146] = t[153] ? t[148] : t[118];
  assign t[147] = t[153] ? t[117] : t[149];
  assign t[148] = ~(x[4] & t[65]);
  assign t[149] = ~(t[131] & t[156]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[153] ? t[116] : t[117];
  assign t[151] = t[153] ? t[118] : t[148];
  assign t[152] = (t[184]);
  assign t[153] = (t[185]);
  assign t[154] = (t[186]);
  assign t[155] = (t[187]);
  assign t[156] = (t[188]);
  assign t[157] = (t[189]);
  assign t[158] = (t[190]);
  assign t[159] = (t[191]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[192]);
  assign t[161] = (t[193]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[153] & t[154]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[155] & t[156]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = t[216] ^ x[2];
  assign t[185] = t[217] ^ x[10];
  assign t[186] = t[218] ^ x[13];
  assign t[187] = t[219] ^ x[16];
  assign t[188] = t[220] ^ x[19];
  assign t[189] = t[221] ^ x[22];
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = t[222] ^ x[25];
  assign t[191] = t[223] ^ x[28];
  assign t[192] = t[224] ^ x[31];
  assign t[193] = t[225] ^ x[34];
  assign t[194] = t[226] ^ x[37];
  assign t[195] = t[227] ^ x[40];
  assign t[196] = t[228] ^ x[43];
  assign t[197] = t[229] ^ x[46];
  assign t[198] = t[230] ^ x[51];
  assign t[199] = t[231] ^ x[54];
  assign t[19] = t[27] ? x[7] : x[6];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[57];
  assign t[201] = t[233] ^ x[60];
  assign t[202] = t[234] ^ x[65];
  assign t[203] = t[235] ^ x[68];
  assign t[204] = t[236] ^ x[71];
  assign t[205] = t[237] ^ x[76];
  assign t[206] = t[238] ^ x[79];
  assign t[207] = t[239] ^ x[82];
  assign t[208] = t[240] ^ x[85];
  assign t[209] = t[241] ^ x[88];
  assign t[20] = t[28] | t[29];
  assign t[210] = t[242] ^ x[91];
  assign t[211] = t[243] ^ x[94];
  assign t[212] = t[244] ^ x[97];
  assign t[213] = t[245] ^ x[100];
  assign t[214] = t[246] ^ x[103];
  assign t[215] = t[247] ^ x[106];
  assign t[216] = (t[248] & ~t[249]);
  assign t[217] = (t[250] & ~t[251]);
  assign t[218] = (t[252] & ~t[253]);
  assign t[219] = (t[254] & ~t[255]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = (t[256] & ~t[257]);
  assign t[221] = (t[258] & ~t[259]);
  assign t[222] = (t[260] & ~t[261]);
  assign t[223] = (t[262] & ~t[263]);
  assign t[224] = (t[264] & ~t[265]);
  assign t[225] = (t[266] & ~t[267]);
  assign t[226] = (t[268] & ~t[269]);
  assign t[227] = (t[270] & ~t[271]);
  assign t[228] = (t[272] & ~t[273]);
  assign t[229] = (t[274] & ~t[275]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (t[276] & ~t[277]);
  assign t[231] = (t[278] & ~t[279]);
  assign t[232] = (t[280] & ~t[281]);
  assign t[233] = (t[282] & ~t[283]);
  assign t[234] = (t[284] & ~t[285]);
  assign t[235] = (t[286] & ~t[287]);
  assign t[236] = (t[288] & ~t[289]);
  assign t[237] = (t[290] & ~t[291]);
  assign t[238] = (t[292] & ~t[293]);
  assign t[239] = (t[294] & ~t[295]);
  assign t[23] = x[4] ? t[33] : t[32];
  assign t[240] = (t[296] & ~t[297]);
  assign t[241] = (t[298] & ~t[299]);
  assign t[242] = (t[300] & ~t[301]);
  assign t[243] = (t[302] & ~t[303]);
  assign t[244] = (t[304] & ~t[305]);
  assign t[245] = (t[306] & ~t[307]);
  assign t[246] = (t[308] & ~t[309]);
  assign t[247] = (t[310] & ~t[311]);
  assign t[248] = t[312] ^ x[2];
  assign t[249] = t[313] ^ x[1];
  assign t[24] = x[4] ? t[35] : t[34];
  assign t[250] = t[314] ^ x[10];
  assign t[251] = t[315] ^ x[9];
  assign t[252] = t[316] ^ x[13];
  assign t[253] = t[317] ^ x[12];
  assign t[254] = t[318] ^ x[16];
  assign t[255] = t[319] ^ x[15];
  assign t[256] = t[320] ^ x[19];
  assign t[257] = t[321] ^ x[18];
  assign t[258] = t[322] ^ x[22];
  assign t[259] = t[323] ^ x[21];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[324] ^ x[25];
  assign t[261] = t[325] ^ x[24];
  assign t[262] = t[326] ^ x[28];
  assign t[263] = t[327] ^ x[27];
  assign t[264] = t[328] ^ x[31];
  assign t[265] = t[329] ^ x[30];
  assign t[266] = t[330] ^ x[34];
  assign t[267] = t[331] ^ x[33];
  assign t[268] = t[332] ^ x[37];
  assign t[269] = t[333] ^ x[36];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[334] ^ x[40];
  assign t[271] = t[335] ^ x[39];
  assign t[272] = t[336] ^ x[43];
  assign t[273] = t[337] ^ x[42];
  assign t[274] = t[338] ^ x[46];
  assign t[275] = t[339] ^ x[45];
  assign t[276] = t[340] ^ x[51];
  assign t[277] = t[341] ^ x[50];
  assign t[278] = t[342] ^ x[54];
  assign t[279] = t[343] ^ x[53];
  assign t[27] = ~(t[40]);
  assign t[280] = t[344] ^ x[57];
  assign t[281] = t[345] ^ x[56];
  assign t[282] = t[346] ^ x[60];
  assign t[283] = t[347] ^ x[59];
  assign t[284] = t[348] ^ x[65];
  assign t[285] = t[349] ^ x[64];
  assign t[286] = t[350] ^ x[68];
  assign t[287] = t[351] ^ x[67];
  assign t[288] = t[352] ^ x[71];
  assign t[289] = t[353] ^ x[70];
  assign t[28] = ~(t[41] & t[42]);
  assign t[290] = t[354] ^ x[76];
  assign t[291] = t[355] ^ x[75];
  assign t[292] = t[356] ^ x[79];
  assign t[293] = t[357] ^ x[78];
  assign t[294] = t[358] ^ x[82];
  assign t[295] = t[359] ^ x[81];
  assign t[296] = t[360] ^ x[85];
  assign t[297] = t[361] ^ x[84];
  assign t[298] = t[362] ^ x[88];
  assign t[299] = t[363] ^ x[87];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[364] ^ x[91];
  assign t[301] = t[365] ^ x[90];
  assign t[302] = t[366] ^ x[94];
  assign t[303] = t[367] ^ x[93];
  assign t[304] = t[368] ^ x[97];
  assign t[305] = t[369] ^ x[96];
  assign t[306] = t[370] ^ x[100];
  assign t[307] = t[371] ^ x[99];
  assign t[308] = t[372] ^ x[103];
  assign t[309] = t[373] ^ x[102];
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = t[374] ^ x[106];
  assign t[311] = t[375] ^ x[105];
  assign t[312] = (x[0]);
  assign t[313] = (x[0]);
  assign t[314] = (x[8]);
  assign t[315] = (x[8]);
  assign t[316] = (x[11]);
  assign t[317] = (x[11]);
  assign t[318] = (x[14]);
  assign t[319] = (x[14]);
  assign t[31] = ~(t[157] | t[47]);
  assign t[320] = (x[17]);
  assign t[321] = (x[17]);
  assign t[322] = (x[20]);
  assign t[323] = (x[20]);
  assign t[324] = (x[23]);
  assign t[325] = (x[23]);
  assign t[326] = (x[26]);
  assign t[327] = (x[26]);
  assign t[328] = (x[29]);
  assign t[329] = (x[29]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[32]);
  assign t[331] = (x[32]);
  assign t[332] = (x[35]);
  assign t[333] = (x[35]);
  assign t[334] = (x[38]);
  assign t[335] = (x[38]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[44]);
  assign t[339] = (x[44]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[58]);
  assign t[347] = (x[58]);
  assign t[348] = (x[63]);
  assign t[349] = (x[63]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = (x[66]);
  assign t[351] = (x[66]);
  assign t[352] = (x[69]);
  assign t[353] = (x[69]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[37] = ~(t[158] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[155]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = ~(t[67]);
  assign t[44] = t[153] ? t[69] : t[68];
  assign t[45] = ~(t[159]);
  assign t[46] = ~(t[160]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[161] | t[74]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[162] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[163]);
  assign t[57] = ~(t[164]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[165] | t[90]);
  assign t[61] = t[27] ? x[48] : x[47];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[67] | t[93]);
  assign t[64] = ~(t[67] | t[94]);
  assign t[65] = ~(t[154] | t[95]);
  assign t[66] = t[43] & t[153];
  assign t[67] = ~(t[155]);
  assign t[68] = ~(x[4] & t[96]);
  assign t[69] = ~(t[156] & t[97]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[166]);
  assign t[71] = ~(t[159] | t[160]);
  assign t[72] = ~(t[167]);
  assign t[73] = ~(t[168]);
  assign t[74] = ~(t[98] | t[99]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[169] | t[102]);
  assign t[77] = t[103] ? x[62] : x[61];
  assign t[78] = ~(t[104] & t[105]);
  assign t[79] = ~(t[170]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[171]);
  assign t[81] = ~(t[106] | t[107]);
  assign t[82] = ~(t[108] | t[109]);
  assign t[83] = ~(t[172] | t[110]);
  assign t[84] = t[103] ? x[73] : x[72];
  assign t[85] = ~(t[111] & t[42]);
  assign t[86] = ~(t[152]);
  assign t[87] = ~(t[163] | t[164]);
  assign t[88] = ~(t[173]);
  assign t[89] = ~(t[174]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112] | t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = ~(t[115] | t[29]);
  assign t[93] = t[153] ? t[117] : t[116];
  assign t[94] = t[153] ? t[118] : t[68];
  assign t[95] = ~(t[156]);
  assign t[96] = ~(t[154] | t[156]);
  assign t[97] = ~(x[4] | t[119]);
  assign t[98] = ~(t[175]);
  assign t[99] = ~(t[167] | t[168]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [88:0] x;
 output y;

 wire [254:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = t[126] ^ x[10];
  assign t[101] = t[127] ^ x[13];
  assign t[102] = t[128] ^ x[16];
  assign t[103] = t[129] ^ x[19];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[25];
  assign t[106] = t[132] ^ x[28];
  assign t[107] = t[133] ^ x[31];
  assign t[108] = t[134] ^ x[36];
  assign t[109] = t[135] ^ x[39];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[42];
  assign t[111] = t[137] ^ x[47];
  assign t[112] = t[138] ^ x[50];
  assign t[113] = t[139] ^ x[55];
  assign t[114] = t[140] ^ x[58];
  assign t[115] = t[141] ^ x[61];
  assign t[116] = t[142] ^ x[64];
  assign t[117] = t[143] ^ x[67];
  assign t[118] = t[144] ^ x[70];
  assign t[119] = t[145] ^ x[73];
  assign t[11] = ~(x[3]);
  assign t[120] = t[146] ^ x[76];
  assign t[121] = t[147] ^ x[79];
  assign t[122] = t[148] ^ x[82];
  assign t[123] = t[149] ^ x[85];
  assign t[124] = t[150] ^ x[88];
  assign t[125] = (t[151] & ~t[152]);
  assign t[126] = (t[153] & ~t[154]);
  assign t[127] = (t[155] & ~t[156]);
  assign t[128] = (t[157] & ~t[158]);
  assign t[129] = (t[159] & ~t[160]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[161] & ~t[162]);
  assign t[131] = (t[163] & ~t[164]);
  assign t[132] = (t[165] & ~t[166]);
  assign t[133] = (t[167] & ~t[168]);
  assign t[134] = (t[169] & ~t[170]);
  assign t[135] = (t[171] & ~t[172]);
  assign t[136] = (t[173] & ~t[174]);
  assign t[137] = (t[175] & ~t[176]);
  assign t[138] = (t[177] & ~t[178]);
  assign t[139] = (t[179] & ~t[180]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (t[181] & ~t[182]);
  assign t[141] = (t[183] & ~t[184]);
  assign t[142] = (t[185] & ~t[186]);
  assign t[143] = (t[187] & ~t[188]);
  assign t[144] = (t[189] & ~t[190]);
  assign t[145] = (t[191] & ~t[192]);
  assign t[146] = (t[193] & ~t[194]);
  assign t[147] = (t[195] & ~t[196]);
  assign t[148] = (t[197] & ~t[198]);
  assign t[149] = (t[199] & ~t[200]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[201] & ~t[202]);
  assign t[151] = t[203] ^ x[2];
  assign t[152] = t[204] ^ x[1];
  assign t[153] = t[205] ^ x[10];
  assign t[154] = t[206] ^ x[9];
  assign t[155] = t[207] ^ x[13];
  assign t[156] = t[208] ^ x[12];
  assign t[157] = t[209] ^ x[16];
  assign t[158] = t[210] ^ x[15];
  assign t[159] = t[211] ^ x[19];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[212] ^ x[18];
  assign t[161] = t[213] ^ x[22];
  assign t[162] = t[214] ^ x[21];
  assign t[163] = t[215] ^ x[25];
  assign t[164] = t[216] ^ x[24];
  assign t[165] = t[217] ^ x[28];
  assign t[166] = t[218] ^ x[27];
  assign t[167] = t[219] ^ x[31];
  assign t[168] = t[220] ^ x[30];
  assign t[169] = t[221] ^ x[36];
  assign t[16] = ~(t[74] & t[75]);
  assign t[170] = t[222] ^ x[35];
  assign t[171] = t[223] ^ x[39];
  assign t[172] = t[224] ^ x[38];
  assign t[173] = t[225] ^ x[42];
  assign t[174] = t[226] ^ x[41];
  assign t[175] = t[227] ^ x[47];
  assign t[176] = t[228] ^ x[46];
  assign t[177] = t[229] ^ x[50];
  assign t[178] = t[230] ^ x[49];
  assign t[179] = t[231] ^ x[55];
  assign t[17] = ~(t[76] & t[77]);
  assign t[180] = t[232] ^ x[54];
  assign t[181] = t[233] ^ x[58];
  assign t[182] = t[234] ^ x[57];
  assign t[183] = t[235] ^ x[61];
  assign t[184] = t[236] ^ x[60];
  assign t[185] = t[237] ^ x[64];
  assign t[186] = t[238] ^ x[63];
  assign t[187] = t[239] ^ x[67];
  assign t[188] = t[240] ^ x[66];
  assign t[189] = t[241] ^ x[70];
  assign t[18] = ~(t[24]);
  assign t[190] = t[242] ^ x[69];
  assign t[191] = t[243] ^ x[73];
  assign t[192] = t[244] ^ x[72];
  assign t[193] = t[245] ^ x[76];
  assign t[194] = t[246] ^ x[75];
  assign t[195] = t[247] ^ x[79];
  assign t[196] = t[248] ^ x[78];
  assign t[197] = t[249] ^ x[82];
  assign t[198] = t[250] ^ x[81];
  assign t[199] = t[251] ^ x[85];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[252] ^ x[84];
  assign t[201] = t[253] ^ x[88];
  assign t[202] = t[254] ^ x[87];
  assign t[203] = (x[0]);
  assign t[204] = (x[0]);
  assign t[205] = (x[8]);
  assign t[206] = (x[8]);
  assign t[207] = (x[11]);
  assign t[208] = (x[11]);
  assign t[209] = (x[14]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[14]);
  assign t[211] = (x[17]);
  assign t[212] = (x[17]);
  assign t[213] = (x[20]);
  assign t[214] = (x[20]);
  assign t[215] = (x[23]);
  assign t[216] = (x[23]);
  assign t[217] = (x[26]);
  assign t[218] = (x[26]);
  assign t[219] = (x[29]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[29]);
  assign t[221] = (x[34]);
  assign t[222] = (x[34]);
  assign t[223] = (x[37]);
  assign t[224] = (x[37]);
  assign t[225] = (x[40]);
  assign t[226] = (x[40]);
  assign t[227] = (x[45]);
  assign t[228] = (x[45]);
  assign t[229] = (x[48]);
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = (x[48]);
  assign t[231] = (x[53]);
  assign t[232] = (x[53]);
  assign t[233] = (x[56]);
  assign t[234] = (x[56]);
  assign t[235] = (x[59]);
  assign t[236] = (x[59]);
  assign t[237] = (x[62]);
  assign t[238] = (x[62]);
  assign t[239] = (x[65]);
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[65]);
  assign t[241] = (x[68]);
  assign t[242] = (x[68]);
  assign t[243] = (x[71]);
  assign t[244] = (x[71]);
  assign t[245] = (x[74]);
  assign t[246] = (x[74]);
  assign t[247] = (x[77]);
  assign t[248] = (x[77]);
  assign t[249] = (x[80]);
  assign t[24] = ~(t[76]);
  assign t[250] = (x[80]);
  assign t[251] = (x[83]);
  assign t[252] = (x[83]);
  assign t[253] = (x[86]);
  assign t[254] = (x[86]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[78] & t[37]);
  assign t[28] = ~(t[79] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[80] & t[47]);
  assign t[34] = ~(t[81] & t[48]);
  assign t[35] = t[18] ? x[33] : x[32];
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[82]);
  assign t[38] = ~(t[82] & t[51]);
  assign t[39] = ~(t[83] & t[52]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[84] & t[53]);
  assign t[41] = t[54] ? x[44] : x[43];
  assign t[42] = ~(t[55] & t[56]);
  assign t[43] = ~(t[85] & t[57]);
  assign t[44] = ~(t[86] & t[58]);
  assign t[45] = t[54] ? x[52] : x[51];
  assign t[46] = ~(t[59] & t[60]);
  assign t[47] = ~(t[87]);
  assign t[48] = ~(t[87] & t[61]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[78]);
  assign t[52] = ~(t[90]);
  assign t[53] = ~(t[90] & t[64]);
  assign t[54] = ~(t[24]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[80]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[96] & t[70]);
  assign t[64] = ~(t[83]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[97] & t[71]);
  assign t[67] = ~(t[85]);
  assign t[68] = ~(t[98]);
  assign t[69] = ~(t[98] & t[72]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[88]);
  assign t[71] = ~(t[91]);
  assign t[72] = ~(t[94]);
  assign t[73] = (t[99]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = t[125] ^ x[2];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind231(x, y);
 input [88:0] x;
 output y;

 wire [254:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = t[126] ^ x[10];
  assign t[101] = t[127] ^ x[13];
  assign t[102] = t[128] ^ x[16];
  assign t[103] = t[129] ^ x[19];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[25];
  assign t[106] = t[132] ^ x[28];
  assign t[107] = t[133] ^ x[31];
  assign t[108] = t[134] ^ x[36];
  assign t[109] = t[135] ^ x[39];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[42];
  assign t[111] = t[137] ^ x[47];
  assign t[112] = t[138] ^ x[50];
  assign t[113] = t[139] ^ x[55];
  assign t[114] = t[140] ^ x[58];
  assign t[115] = t[141] ^ x[61];
  assign t[116] = t[142] ^ x[64];
  assign t[117] = t[143] ^ x[67];
  assign t[118] = t[144] ^ x[70];
  assign t[119] = t[145] ^ x[73];
  assign t[11] = ~(x[3]);
  assign t[120] = t[146] ^ x[76];
  assign t[121] = t[147] ^ x[79];
  assign t[122] = t[148] ^ x[82];
  assign t[123] = t[149] ^ x[85];
  assign t[124] = t[150] ^ x[88];
  assign t[125] = (t[151] & ~t[152]);
  assign t[126] = (t[153] & ~t[154]);
  assign t[127] = (t[155] & ~t[156]);
  assign t[128] = (t[157] & ~t[158]);
  assign t[129] = (t[159] & ~t[160]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[161] & ~t[162]);
  assign t[131] = (t[163] & ~t[164]);
  assign t[132] = (t[165] & ~t[166]);
  assign t[133] = (t[167] & ~t[168]);
  assign t[134] = (t[169] & ~t[170]);
  assign t[135] = (t[171] & ~t[172]);
  assign t[136] = (t[173] & ~t[174]);
  assign t[137] = (t[175] & ~t[176]);
  assign t[138] = (t[177] & ~t[178]);
  assign t[139] = (t[179] & ~t[180]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (t[181] & ~t[182]);
  assign t[141] = (t[183] & ~t[184]);
  assign t[142] = (t[185] & ~t[186]);
  assign t[143] = (t[187] & ~t[188]);
  assign t[144] = (t[189] & ~t[190]);
  assign t[145] = (t[191] & ~t[192]);
  assign t[146] = (t[193] & ~t[194]);
  assign t[147] = (t[195] & ~t[196]);
  assign t[148] = (t[197] & ~t[198]);
  assign t[149] = (t[199] & ~t[200]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[201] & ~t[202]);
  assign t[151] = t[203] ^ x[2];
  assign t[152] = t[204] ^ x[1];
  assign t[153] = t[205] ^ x[10];
  assign t[154] = t[206] ^ x[9];
  assign t[155] = t[207] ^ x[13];
  assign t[156] = t[208] ^ x[12];
  assign t[157] = t[209] ^ x[16];
  assign t[158] = t[210] ^ x[15];
  assign t[159] = t[211] ^ x[19];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[212] ^ x[18];
  assign t[161] = t[213] ^ x[22];
  assign t[162] = t[214] ^ x[21];
  assign t[163] = t[215] ^ x[25];
  assign t[164] = t[216] ^ x[24];
  assign t[165] = t[217] ^ x[28];
  assign t[166] = t[218] ^ x[27];
  assign t[167] = t[219] ^ x[31];
  assign t[168] = t[220] ^ x[30];
  assign t[169] = t[221] ^ x[36];
  assign t[16] = ~(t[74] & t[75]);
  assign t[170] = t[222] ^ x[35];
  assign t[171] = t[223] ^ x[39];
  assign t[172] = t[224] ^ x[38];
  assign t[173] = t[225] ^ x[42];
  assign t[174] = t[226] ^ x[41];
  assign t[175] = t[227] ^ x[47];
  assign t[176] = t[228] ^ x[46];
  assign t[177] = t[229] ^ x[50];
  assign t[178] = t[230] ^ x[49];
  assign t[179] = t[231] ^ x[55];
  assign t[17] = ~(t[76] & t[77]);
  assign t[180] = t[232] ^ x[54];
  assign t[181] = t[233] ^ x[58];
  assign t[182] = t[234] ^ x[57];
  assign t[183] = t[235] ^ x[61];
  assign t[184] = t[236] ^ x[60];
  assign t[185] = t[237] ^ x[64];
  assign t[186] = t[238] ^ x[63];
  assign t[187] = t[239] ^ x[67];
  assign t[188] = t[240] ^ x[66];
  assign t[189] = t[241] ^ x[70];
  assign t[18] = ~(t[24]);
  assign t[190] = t[242] ^ x[69];
  assign t[191] = t[243] ^ x[73];
  assign t[192] = t[244] ^ x[72];
  assign t[193] = t[245] ^ x[76];
  assign t[194] = t[246] ^ x[75];
  assign t[195] = t[247] ^ x[79];
  assign t[196] = t[248] ^ x[78];
  assign t[197] = t[249] ^ x[82];
  assign t[198] = t[250] ^ x[81];
  assign t[199] = t[251] ^ x[85];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[252] ^ x[84];
  assign t[201] = t[253] ^ x[88];
  assign t[202] = t[254] ^ x[87];
  assign t[203] = (x[0]);
  assign t[204] = (x[0]);
  assign t[205] = (x[8]);
  assign t[206] = (x[8]);
  assign t[207] = (x[11]);
  assign t[208] = (x[11]);
  assign t[209] = (x[14]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[14]);
  assign t[211] = (x[17]);
  assign t[212] = (x[17]);
  assign t[213] = (x[20]);
  assign t[214] = (x[20]);
  assign t[215] = (x[23]);
  assign t[216] = (x[23]);
  assign t[217] = (x[26]);
  assign t[218] = (x[26]);
  assign t[219] = (x[29]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[29]);
  assign t[221] = (x[34]);
  assign t[222] = (x[34]);
  assign t[223] = (x[37]);
  assign t[224] = (x[37]);
  assign t[225] = (x[40]);
  assign t[226] = (x[40]);
  assign t[227] = (x[45]);
  assign t[228] = (x[45]);
  assign t[229] = (x[48]);
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = (x[48]);
  assign t[231] = (x[53]);
  assign t[232] = (x[53]);
  assign t[233] = (x[56]);
  assign t[234] = (x[56]);
  assign t[235] = (x[59]);
  assign t[236] = (x[59]);
  assign t[237] = (x[62]);
  assign t[238] = (x[62]);
  assign t[239] = (x[65]);
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[65]);
  assign t[241] = (x[68]);
  assign t[242] = (x[68]);
  assign t[243] = (x[71]);
  assign t[244] = (x[71]);
  assign t[245] = (x[74]);
  assign t[246] = (x[74]);
  assign t[247] = (x[77]);
  assign t[248] = (x[77]);
  assign t[249] = (x[80]);
  assign t[24] = ~(t[76]);
  assign t[250] = (x[80]);
  assign t[251] = (x[83]);
  assign t[252] = (x[83]);
  assign t[253] = (x[86]);
  assign t[254] = (x[86]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[78] & t[37]);
  assign t[28] = ~(t[79] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[80] & t[47]);
  assign t[34] = ~(t[81] & t[48]);
  assign t[35] = t[18] ? x[33] : x[32];
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[82]);
  assign t[38] = ~(t[82] & t[51]);
  assign t[39] = ~(t[83] & t[52]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[84] & t[53]);
  assign t[41] = t[54] ? x[44] : x[43];
  assign t[42] = ~(t[55] & t[56]);
  assign t[43] = ~(t[85] & t[57]);
  assign t[44] = ~(t[86] & t[58]);
  assign t[45] = t[54] ? x[52] : x[51];
  assign t[46] = ~(t[59] & t[60]);
  assign t[47] = ~(t[87]);
  assign t[48] = ~(t[87] & t[61]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[78]);
  assign t[52] = ~(t[90]);
  assign t[53] = ~(t[90] & t[64]);
  assign t[54] = ~(t[24]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[80]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[96] & t[70]);
  assign t[64] = ~(t[83]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[97] & t[71]);
  assign t[67] = ~(t[85]);
  assign t[68] = ~(t[98]);
  assign t[69] = ~(t[98] & t[72]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[88]);
  assign t[71] = ~(t[91]);
  assign t[72] = ~(t[94]);
  assign t[73] = (t[99]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = t[125] ^ x[2];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [106:0] x;
 output y;

 wire [310:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[2];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[10];
  assign t[121] = t[153] ^ x[13];
  assign t[122] = t[154] ^ x[16];
  assign t[123] = t[155] ^ x[19];
  assign t[124] = t[156] ^ x[22];
  assign t[125] = t[157] ^ x[25];
  assign t[126] = t[158] ^ x[30];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[36];
  assign t[129] = t[161] ^ x[41];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[46];
  assign t[131] = t[163] ^ x[49];
  assign t[132] = t[164] ^ x[52];
  assign t[133] = t[165] ^ x[55];
  assign t[134] = t[166] ^ x[58];
  assign t[135] = t[167] ^ x[61];
  assign t[136] = t[168] ^ x[64];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[70];
  assign t[139] = t[171] ^ x[73];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[76];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[82];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = t[176] ^ x[88];
  assign t[145] = t[177] ^ x[91];
  assign t[146] = t[178] ^ x[94];
  assign t[147] = t[179] ^ x[97];
  assign t[148] = t[180] ^ x[100];
  assign t[149] = t[181] ^ x[103];
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = t[182] ^ x[106];
  assign t[151] = (t[183] & ~t[184]);
  assign t[152] = (t[185] & ~t[186]);
  assign t[153] = (t[187] & ~t[188]);
  assign t[154] = (t[189] & ~t[190]);
  assign t[155] = (t[191] & ~t[192]);
  assign t[156] = (t[193] & ~t[194]);
  assign t[157] = (t[195] & ~t[196]);
  assign t[158] = (t[197] & ~t[198]);
  assign t[159] = (t[199] & ~t[200]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[201] & ~t[202]);
  assign t[161] = (t[203] & ~t[204]);
  assign t[162] = (t[205] & ~t[206]);
  assign t[163] = (t[207] & ~t[208]);
  assign t[164] = (t[209] & ~t[210]);
  assign t[165] = (t[211] & ~t[212]);
  assign t[166] = (t[213] & ~t[214]);
  assign t[167] = (t[215] & ~t[216]);
  assign t[168] = (t[217] & ~t[218]);
  assign t[169] = (t[219] & ~t[220]);
  assign t[16] = ~(t[88] & t[89]);
  assign t[170] = (t[221] & ~t[222]);
  assign t[171] = (t[223] & ~t[224]);
  assign t[172] = (t[225] & ~t[226]);
  assign t[173] = (t[227] & ~t[228]);
  assign t[174] = (t[229] & ~t[230]);
  assign t[175] = (t[231] & ~t[232]);
  assign t[176] = (t[233] & ~t[234]);
  assign t[177] = (t[235] & ~t[236]);
  assign t[178] = (t[237] & ~t[238]);
  assign t[179] = (t[239] & ~t[240]);
  assign t[17] = ~(t[90] & t[91]);
  assign t[180] = (t[241] & ~t[242]);
  assign t[181] = (t[243] & ~t[244]);
  assign t[182] = (t[245] & ~t[246]);
  assign t[183] = t[247] ^ x[2];
  assign t[184] = t[248] ^ x[1];
  assign t[185] = t[249] ^ x[10];
  assign t[186] = t[250] ^ x[9];
  assign t[187] = t[251] ^ x[13];
  assign t[188] = t[252] ^ x[12];
  assign t[189] = t[253] ^ x[16];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[15];
  assign t[191] = t[255] ^ x[19];
  assign t[192] = t[256] ^ x[18];
  assign t[193] = t[257] ^ x[22];
  assign t[194] = t[258] ^ x[21];
  assign t[195] = t[259] ^ x[25];
  assign t[196] = t[260] ^ x[24];
  assign t[197] = t[261] ^ x[30];
  assign t[198] = t[262] ^ x[29];
  assign t[199] = t[263] ^ x[33];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[32];
  assign t[201] = t[265] ^ x[36];
  assign t[202] = t[266] ^ x[35];
  assign t[203] = t[267] ^ x[41];
  assign t[204] = t[268] ^ x[40];
  assign t[205] = t[269] ^ x[46];
  assign t[206] = t[270] ^ x[45];
  assign t[207] = t[271] ^ x[49];
  assign t[208] = t[272] ^ x[48];
  assign t[209] = t[273] ^ x[52];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[51];
  assign t[211] = t[275] ^ x[55];
  assign t[212] = t[276] ^ x[54];
  assign t[213] = t[277] ^ x[58];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[61];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[64];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[67];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[70];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[73];
  assign t[224] = t[288] ^ x[72];
  assign t[225] = t[289] ^ x[76];
  assign t[226] = t[290] ^ x[75];
  assign t[227] = t[291] ^ x[79];
  assign t[228] = t[292] ^ x[78];
  assign t[229] = t[293] ^ x[82];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[81];
  assign t[231] = t[295] ^ x[85];
  assign t[232] = t[296] ^ x[84];
  assign t[233] = t[297] ^ x[88];
  assign t[234] = t[298] ^ x[87];
  assign t[235] = t[299] ^ x[91];
  assign t[236] = t[300] ^ x[90];
  assign t[237] = t[301] ^ x[94];
  assign t[238] = t[302] ^ x[93];
  assign t[239] = t[303] ^ x[97];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = t[304] ^ x[96];
  assign t[241] = t[305] ^ x[100];
  assign t[242] = t[306] ^ x[99];
  assign t[243] = t[307] ^ x[103];
  assign t[244] = t[308] ^ x[102];
  assign t[245] = t[309] ^ x[106];
  assign t[246] = t[310] ^ x[105];
  assign t[247] = (x[0]);
  assign t[248] = (x[0]);
  assign t[249] = (x[8]);
  assign t[24] = ~(t[90]);
  assign t[250] = (x[8]);
  assign t[251] = (x[11]);
  assign t[252] = (x[11]);
  assign t[253] = (x[14]);
  assign t[254] = (x[14]);
  assign t[255] = (x[17]);
  assign t[256] = (x[17]);
  assign t[257] = (x[20]);
  assign t[258] = (x[20]);
  assign t[259] = (x[23]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[23]);
  assign t[261] = (x[28]);
  assign t[262] = (x[28]);
  assign t[263] = (x[31]);
  assign t[264] = (x[31]);
  assign t[265] = (x[34]);
  assign t[266] = (x[34]);
  assign t[267] = (x[39]);
  assign t[268] = (x[39]);
  assign t[269] = (x[44]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[44]);
  assign t[271] = (x[47]);
  assign t[272] = (x[47]);
  assign t[273] = (x[50]);
  assign t[274] = (x[50]);
  assign t[275] = (x[53]);
  assign t[276] = (x[53]);
  assign t[277] = (x[56]);
  assign t[278] = (x[56]);
  assign t[279] = (x[59]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[59]);
  assign t[281] = (x[62]);
  assign t[282] = (x[62]);
  assign t[283] = (x[65]);
  assign t[284] = (x[65]);
  assign t[285] = (x[68]);
  assign t[286] = (x[68]);
  assign t[287] = (x[71]);
  assign t[288] = (x[71]);
  assign t[289] = (x[74]);
  assign t[28] = ~(t[39] & t[92]);
  assign t[290] = (x[74]);
  assign t[291] = (x[77]);
  assign t[292] = (x[77]);
  assign t[293] = (x[80]);
  assign t[294] = (x[80]);
  assign t[295] = (x[83]);
  assign t[296] = (x[83]);
  assign t[297] = (x[86]);
  assign t[298] = (x[86]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[89]);
  assign t[301] = (x[92]);
  assign t[302] = (x[92]);
  assign t[303] = (x[95]);
  assign t[304] = (x[95]);
  assign t[305] = (x[98]);
  assign t[306] = (x[98]);
  assign t[307] = (x[101]);
  assign t[308] = (x[101]);
  assign t[309] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[310] = (x[104]);
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[93]);
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[94]);
  assign t[38] = ~(t[95]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[96]);
  assign t[42] = t[58] ? x[38] : x[37];
  assign t[43] = ~(t[59] & t[60]);
  assign t[44] = ~(t[61] & t[62]);
  assign t[45] = ~(t[63] & t[97]);
  assign t[46] = t[58] ? x[43] : x[42];
  assign t[47] = ~(t[64] & t[65]);
  assign t[48] = ~(t[98]);
  assign t[49] = ~(t[99]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[66] & t[67]);
  assign t[51] = ~(t[68] & t[69]);
  assign t[52] = ~(t[70] & t[100]);
  assign t[53] = ~(t[95] & t[94]);
  assign t[54] = ~(t[101]);
  assign t[55] = ~(t[102]);
  assign t[56] = ~(t[103]);
  assign t[57] = ~(t[71] & t[72]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[73] & t[74]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[75] & t[104]);
  assign t[61] = ~(t[105]);
  assign t[62] = ~(t[106]);
  assign t[63] = ~(t[76] & t[77]);
  assign t[64] = ~(t[78] & t[79]);
  assign t[65] = ~(t[80] & t[107]);
  assign t[66] = ~(t[99] & t[98]);
  assign t[67] = ~(t[87]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [106:0] x;
 output y;

 wire [310:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[2];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[10];
  assign t[121] = t[153] ^ x[13];
  assign t[122] = t[154] ^ x[16];
  assign t[123] = t[155] ^ x[19];
  assign t[124] = t[156] ^ x[22];
  assign t[125] = t[157] ^ x[25];
  assign t[126] = t[158] ^ x[30];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[36];
  assign t[129] = t[161] ^ x[41];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[46];
  assign t[131] = t[163] ^ x[49];
  assign t[132] = t[164] ^ x[52];
  assign t[133] = t[165] ^ x[55];
  assign t[134] = t[166] ^ x[58];
  assign t[135] = t[167] ^ x[61];
  assign t[136] = t[168] ^ x[64];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[70];
  assign t[139] = t[171] ^ x[73];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[76];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[82];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = t[176] ^ x[88];
  assign t[145] = t[177] ^ x[91];
  assign t[146] = t[178] ^ x[94];
  assign t[147] = t[179] ^ x[97];
  assign t[148] = t[180] ^ x[100];
  assign t[149] = t[181] ^ x[103];
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = t[182] ^ x[106];
  assign t[151] = (t[183] & ~t[184]);
  assign t[152] = (t[185] & ~t[186]);
  assign t[153] = (t[187] & ~t[188]);
  assign t[154] = (t[189] & ~t[190]);
  assign t[155] = (t[191] & ~t[192]);
  assign t[156] = (t[193] & ~t[194]);
  assign t[157] = (t[195] & ~t[196]);
  assign t[158] = (t[197] & ~t[198]);
  assign t[159] = (t[199] & ~t[200]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[201] & ~t[202]);
  assign t[161] = (t[203] & ~t[204]);
  assign t[162] = (t[205] & ~t[206]);
  assign t[163] = (t[207] & ~t[208]);
  assign t[164] = (t[209] & ~t[210]);
  assign t[165] = (t[211] & ~t[212]);
  assign t[166] = (t[213] & ~t[214]);
  assign t[167] = (t[215] & ~t[216]);
  assign t[168] = (t[217] & ~t[218]);
  assign t[169] = (t[219] & ~t[220]);
  assign t[16] = ~(t[88] & t[89]);
  assign t[170] = (t[221] & ~t[222]);
  assign t[171] = (t[223] & ~t[224]);
  assign t[172] = (t[225] & ~t[226]);
  assign t[173] = (t[227] & ~t[228]);
  assign t[174] = (t[229] & ~t[230]);
  assign t[175] = (t[231] & ~t[232]);
  assign t[176] = (t[233] & ~t[234]);
  assign t[177] = (t[235] & ~t[236]);
  assign t[178] = (t[237] & ~t[238]);
  assign t[179] = (t[239] & ~t[240]);
  assign t[17] = ~(t[90] & t[91]);
  assign t[180] = (t[241] & ~t[242]);
  assign t[181] = (t[243] & ~t[244]);
  assign t[182] = (t[245] & ~t[246]);
  assign t[183] = t[247] ^ x[2];
  assign t[184] = t[248] ^ x[1];
  assign t[185] = t[249] ^ x[10];
  assign t[186] = t[250] ^ x[9];
  assign t[187] = t[251] ^ x[13];
  assign t[188] = t[252] ^ x[12];
  assign t[189] = t[253] ^ x[16];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[15];
  assign t[191] = t[255] ^ x[19];
  assign t[192] = t[256] ^ x[18];
  assign t[193] = t[257] ^ x[22];
  assign t[194] = t[258] ^ x[21];
  assign t[195] = t[259] ^ x[25];
  assign t[196] = t[260] ^ x[24];
  assign t[197] = t[261] ^ x[30];
  assign t[198] = t[262] ^ x[29];
  assign t[199] = t[263] ^ x[33];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[32];
  assign t[201] = t[265] ^ x[36];
  assign t[202] = t[266] ^ x[35];
  assign t[203] = t[267] ^ x[41];
  assign t[204] = t[268] ^ x[40];
  assign t[205] = t[269] ^ x[46];
  assign t[206] = t[270] ^ x[45];
  assign t[207] = t[271] ^ x[49];
  assign t[208] = t[272] ^ x[48];
  assign t[209] = t[273] ^ x[52];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[51];
  assign t[211] = t[275] ^ x[55];
  assign t[212] = t[276] ^ x[54];
  assign t[213] = t[277] ^ x[58];
  assign t[214] = t[278] ^ x[57];
  assign t[215] = t[279] ^ x[61];
  assign t[216] = t[280] ^ x[60];
  assign t[217] = t[281] ^ x[64];
  assign t[218] = t[282] ^ x[63];
  assign t[219] = t[283] ^ x[67];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[66];
  assign t[221] = t[285] ^ x[70];
  assign t[222] = t[286] ^ x[69];
  assign t[223] = t[287] ^ x[73];
  assign t[224] = t[288] ^ x[72];
  assign t[225] = t[289] ^ x[76];
  assign t[226] = t[290] ^ x[75];
  assign t[227] = t[291] ^ x[79];
  assign t[228] = t[292] ^ x[78];
  assign t[229] = t[293] ^ x[82];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[81];
  assign t[231] = t[295] ^ x[85];
  assign t[232] = t[296] ^ x[84];
  assign t[233] = t[297] ^ x[88];
  assign t[234] = t[298] ^ x[87];
  assign t[235] = t[299] ^ x[91];
  assign t[236] = t[300] ^ x[90];
  assign t[237] = t[301] ^ x[94];
  assign t[238] = t[302] ^ x[93];
  assign t[239] = t[303] ^ x[97];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = t[304] ^ x[96];
  assign t[241] = t[305] ^ x[100];
  assign t[242] = t[306] ^ x[99];
  assign t[243] = t[307] ^ x[103];
  assign t[244] = t[308] ^ x[102];
  assign t[245] = t[309] ^ x[106];
  assign t[246] = t[310] ^ x[105];
  assign t[247] = (x[0]);
  assign t[248] = (x[0]);
  assign t[249] = (x[8]);
  assign t[24] = ~(t[90]);
  assign t[250] = (x[8]);
  assign t[251] = (x[11]);
  assign t[252] = (x[11]);
  assign t[253] = (x[14]);
  assign t[254] = (x[14]);
  assign t[255] = (x[17]);
  assign t[256] = (x[17]);
  assign t[257] = (x[20]);
  assign t[258] = (x[20]);
  assign t[259] = (x[23]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[23]);
  assign t[261] = (x[28]);
  assign t[262] = (x[28]);
  assign t[263] = (x[31]);
  assign t[264] = (x[31]);
  assign t[265] = (x[34]);
  assign t[266] = (x[34]);
  assign t[267] = (x[39]);
  assign t[268] = (x[39]);
  assign t[269] = (x[44]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[44]);
  assign t[271] = (x[47]);
  assign t[272] = (x[47]);
  assign t[273] = (x[50]);
  assign t[274] = (x[50]);
  assign t[275] = (x[53]);
  assign t[276] = (x[53]);
  assign t[277] = (x[56]);
  assign t[278] = (x[56]);
  assign t[279] = (x[59]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[59]);
  assign t[281] = (x[62]);
  assign t[282] = (x[62]);
  assign t[283] = (x[65]);
  assign t[284] = (x[65]);
  assign t[285] = (x[68]);
  assign t[286] = (x[68]);
  assign t[287] = (x[71]);
  assign t[288] = (x[71]);
  assign t[289] = (x[74]);
  assign t[28] = ~(t[39] & t[92]);
  assign t[290] = (x[74]);
  assign t[291] = (x[77]);
  assign t[292] = (x[77]);
  assign t[293] = (x[80]);
  assign t[294] = (x[80]);
  assign t[295] = (x[83]);
  assign t[296] = (x[83]);
  assign t[297] = (x[86]);
  assign t[298] = (x[86]);
  assign t[299] = (x[89]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[89]);
  assign t[301] = (x[92]);
  assign t[302] = (x[92]);
  assign t[303] = (x[95]);
  assign t[304] = (x[95]);
  assign t[305] = (x[98]);
  assign t[306] = (x[98]);
  assign t[307] = (x[101]);
  assign t[308] = (x[101]);
  assign t[309] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[310] = (x[104]);
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[93]);
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[94]);
  assign t[38] = ~(t[95]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[96]);
  assign t[42] = t[58] ? x[38] : x[37];
  assign t[43] = ~(t[59] & t[60]);
  assign t[44] = ~(t[61] & t[62]);
  assign t[45] = ~(t[63] & t[97]);
  assign t[46] = t[58] ? x[43] : x[42];
  assign t[47] = ~(t[64] & t[65]);
  assign t[48] = ~(t[98]);
  assign t[49] = ~(t[99]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[66] & t[67]);
  assign t[51] = ~(t[68] & t[69]);
  assign t[52] = ~(t[70] & t[100]);
  assign t[53] = ~(t[95] & t[94]);
  assign t[54] = ~(t[101]);
  assign t[55] = ~(t[102]);
  assign t[56] = ~(t[103]);
  assign t[57] = ~(t[71] & t[72]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[73] & t[74]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[75] & t[104]);
  assign t[61] = ~(t[105]);
  assign t[62] = ~(t[106]);
  assign t[63] = ~(t[76] & t[77]);
  assign t[64] = ~(t[78] & t[79]);
  assign t[65] = ~(t[80] & t[107]);
  assign t[66] = ~(t[99] & t[98]);
  assign t[67] = ~(t[87]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [106:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[2];
  assign t[113] = t[145] ^ x[10];
  assign t[114] = t[146] ^ x[13];
  assign t[115] = t[147] ^ x[16];
  assign t[116] = t[148] ^ x[19];
  assign t[117] = t[149] ^ x[22];
  assign t[118] = t[150] ^ x[25];
  assign t[119] = t[151] ^ x[30];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[36];
  assign t[122] = t[154] ^ x[41];
  assign t[123] = t[155] ^ x[46];
  assign t[124] = t[156] ^ x[49];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[55];
  assign t[127] = t[159] ^ x[58];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[70];
  assign t[132] = t[164] ^ x[73];
  assign t[133] = t[165] ^ x[76];
  assign t[134] = t[166] ^ x[79];
  assign t[135] = t[167] ^ x[82];
  assign t[136] = t[168] ^ x[85];
  assign t[137] = t[169] ^ x[88];
  assign t[138] = t[170] ^ x[91];
  assign t[139] = t[171] ^ x[94];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[97];
  assign t[141] = t[173] ^ x[100];
  assign t[142] = t[174] ^ x[103];
  assign t[143] = t[175] ^ x[106];
  assign t[144] = (t[176] & ~t[177]);
  assign t[145] = (t[178] & ~t[179]);
  assign t[146] = (t[180] & ~t[181]);
  assign t[147] = (t[182] & ~t[183]);
  assign t[148] = (t[184] & ~t[185]);
  assign t[149] = (t[186] & ~t[187]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[188] & ~t[189]);
  assign t[151] = (t[190] & ~t[191]);
  assign t[152] = (t[192] & ~t[193]);
  assign t[153] = (t[194] & ~t[195]);
  assign t[154] = (t[196] & ~t[197]);
  assign t[155] = (t[198] & ~t[199]);
  assign t[156] = (t[200] & ~t[201]);
  assign t[157] = (t[202] & ~t[203]);
  assign t[158] = (t[204] & ~t[205]);
  assign t[159] = (t[206] & ~t[207]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[208] & ~t[209]);
  assign t[161] = (t[210] & ~t[211]);
  assign t[162] = (t[212] & ~t[213]);
  assign t[163] = (t[214] & ~t[215]);
  assign t[164] = (t[216] & ~t[217]);
  assign t[165] = (t[218] & ~t[219]);
  assign t[166] = (t[220] & ~t[221]);
  assign t[167] = (t[222] & ~t[223]);
  assign t[168] = (t[224] & ~t[225]);
  assign t[169] = (t[226] & ~t[227]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (t[228] & ~t[229]);
  assign t[171] = (t[230] & ~t[231]);
  assign t[172] = (t[232] & ~t[233]);
  assign t[173] = (t[234] & ~t[235]);
  assign t[174] = (t[236] & ~t[237]);
  assign t[175] = (t[238] & ~t[239]);
  assign t[176] = t[240] ^ x[2];
  assign t[177] = t[241] ^ x[1];
  assign t[178] = t[242] ^ x[10];
  assign t[179] = t[243] ^ x[9];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[244] ^ x[13];
  assign t[181] = t[245] ^ x[12];
  assign t[182] = t[246] ^ x[16];
  assign t[183] = t[247] ^ x[15];
  assign t[184] = t[248] ^ x[19];
  assign t[185] = t[249] ^ x[18];
  assign t[186] = t[250] ^ x[22];
  assign t[187] = t[251] ^ x[21];
  assign t[188] = t[252] ^ x[25];
  assign t[189] = t[253] ^ x[24];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[30];
  assign t[191] = t[255] ^ x[29];
  assign t[192] = t[256] ^ x[33];
  assign t[193] = t[257] ^ x[32];
  assign t[194] = t[258] ^ x[36];
  assign t[195] = t[259] ^ x[35];
  assign t[196] = t[260] ^ x[41];
  assign t[197] = t[261] ^ x[40];
  assign t[198] = t[262] ^ x[46];
  assign t[199] = t[263] ^ x[45];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[49];
  assign t[201] = t[265] ^ x[48];
  assign t[202] = t[266] ^ x[52];
  assign t[203] = t[267] ^ x[51];
  assign t[204] = t[268] ^ x[55];
  assign t[205] = t[269] ^ x[54];
  assign t[206] = t[270] ^ x[58];
  assign t[207] = t[271] ^ x[57];
  assign t[208] = t[272] ^ x[61];
  assign t[209] = t[273] ^ x[60];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[64];
  assign t[211] = t[275] ^ x[63];
  assign t[212] = t[276] ^ x[67];
  assign t[213] = t[277] ^ x[66];
  assign t[214] = t[278] ^ x[70];
  assign t[215] = t[279] ^ x[69];
  assign t[216] = t[280] ^ x[73];
  assign t[217] = t[281] ^ x[72];
  assign t[218] = t[282] ^ x[76];
  assign t[219] = t[283] ^ x[75];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[79];
  assign t[221] = t[285] ^ x[78];
  assign t[222] = t[286] ^ x[82];
  assign t[223] = t[287] ^ x[81];
  assign t[224] = t[288] ^ x[85];
  assign t[225] = t[289] ^ x[84];
  assign t[226] = t[290] ^ x[88];
  assign t[227] = t[291] ^ x[87];
  assign t[228] = t[292] ^ x[91];
  assign t[229] = t[293] ^ x[90];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[94];
  assign t[231] = t[295] ^ x[93];
  assign t[232] = t[296] ^ x[97];
  assign t[233] = t[297] ^ x[96];
  assign t[234] = t[298] ^ x[100];
  assign t[235] = t[299] ^ x[99];
  assign t[236] = t[300] ^ x[103];
  assign t[237] = t[301] ^ x[102];
  assign t[238] = t[302] ^ x[106];
  assign t[239] = t[303] ^ x[105];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[0]);
  assign t[241] = (x[0]);
  assign t[242] = (x[8]);
  assign t[243] = (x[8]);
  assign t[244] = (x[11]);
  assign t[245] = (x[11]);
  assign t[246] = (x[14]);
  assign t[247] = (x[14]);
  assign t[248] = (x[17]);
  assign t[249] = (x[17]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[20]);
  assign t[251] = (x[20]);
  assign t[252] = (x[23]);
  assign t[253] = (x[23]);
  assign t[254] = (x[28]);
  assign t[255] = (x[28]);
  assign t[256] = (x[31]);
  assign t[257] = (x[31]);
  assign t[258] = (x[34]);
  assign t[259] = (x[34]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[39]);
  assign t[261] = (x[39]);
  assign t[262] = (x[44]);
  assign t[263] = (x[44]);
  assign t[264] = (x[47]);
  assign t[265] = (x[47]);
  assign t[266] = (x[50]);
  assign t[267] = (x[50]);
  assign t[268] = (x[53]);
  assign t[269] = (x[53]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[56]);
  assign t[271] = (x[56]);
  assign t[272] = (x[59]);
  assign t[273] = (x[59]);
  assign t[274] = (x[62]);
  assign t[275] = (x[62]);
  assign t[276] = (x[65]);
  assign t[277] = (x[65]);
  assign t[278] = (x[68]);
  assign t[279] = (x[68]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[71]);
  assign t[281] = (x[71]);
  assign t[282] = (x[74]);
  assign t[283] = (x[74]);
  assign t[284] = (x[77]);
  assign t[285] = (x[77]);
  assign t[286] = (x[80]);
  assign t[287] = (x[80]);
  assign t[288] = (x[83]);
  assign t[289] = (x[83]);
  assign t[28] = t[39] | t[85];
  assign t[290] = (x[86]);
  assign t[291] = (x[86]);
  assign t[292] = (x[89]);
  assign t[293] = (x[89]);
  assign t[294] = (x[92]);
  assign t[295] = (x[92]);
  assign t[296] = (x[95]);
  assign t[297] = (x[95]);
  assign t[298] = (x[98]);
  assign t[299] = (x[98]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[101]);
  assign t[301] = (x[101]);
  assign t[302] = (x[104]);
  assign t[303] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[57] ? x[38] : x[37];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[60] & t[61]);
  assign t[45] = t[62] | t[90];
  assign t[46] = t[57] ? x[43] : x[42];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[70] & t[71]);
  assign t[59] = t[72] | t[96];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[97]);
  assign t[61] = ~(t[98]);
  assign t[62] = ~(t[73] | t[60]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [106:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[2];
  assign t[113] = t[145] ^ x[10];
  assign t[114] = t[146] ^ x[13];
  assign t[115] = t[147] ^ x[16];
  assign t[116] = t[148] ^ x[19];
  assign t[117] = t[149] ^ x[22];
  assign t[118] = t[150] ^ x[25];
  assign t[119] = t[151] ^ x[30];
  assign t[11] = ~(x[3]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[36];
  assign t[122] = t[154] ^ x[41];
  assign t[123] = t[155] ^ x[46];
  assign t[124] = t[156] ^ x[49];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[55];
  assign t[127] = t[159] ^ x[58];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[70];
  assign t[132] = t[164] ^ x[73];
  assign t[133] = t[165] ^ x[76];
  assign t[134] = t[166] ^ x[79];
  assign t[135] = t[167] ^ x[82];
  assign t[136] = t[168] ^ x[85];
  assign t[137] = t[169] ^ x[88];
  assign t[138] = t[170] ^ x[91];
  assign t[139] = t[171] ^ x[94];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[97];
  assign t[141] = t[173] ^ x[100];
  assign t[142] = t[174] ^ x[103];
  assign t[143] = t[175] ^ x[106];
  assign t[144] = (t[176] & ~t[177]);
  assign t[145] = (t[178] & ~t[179]);
  assign t[146] = (t[180] & ~t[181]);
  assign t[147] = (t[182] & ~t[183]);
  assign t[148] = (t[184] & ~t[185]);
  assign t[149] = (t[186] & ~t[187]);
  assign t[14] = x[4] ? t[21] : t[20];
  assign t[150] = (t[188] & ~t[189]);
  assign t[151] = (t[190] & ~t[191]);
  assign t[152] = (t[192] & ~t[193]);
  assign t[153] = (t[194] & ~t[195]);
  assign t[154] = (t[196] & ~t[197]);
  assign t[155] = (t[198] & ~t[199]);
  assign t[156] = (t[200] & ~t[201]);
  assign t[157] = (t[202] & ~t[203]);
  assign t[158] = (t[204] & ~t[205]);
  assign t[159] = (t[206] & ~t[207]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (t[208] & ~t[209]);
  assign t[161] = (t[210] & ~t[211]);
  assign t[162] = (t[212] & ~t[213]);
  assign t[163] = (t[214] & ~t[215]);
  assign t[164] = (t[216] & ~t[217]);
  assign t[165] = (t[218] & ~t[219]);
  assign t[166] = (t[220] & ~t[221]);
  assign t[167] = (t[222] & ~t[223]);
  assign t[168] = (t[224] & ~t[225]);
  assign t[169] = (t[226] & ~t[227]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (t[228] & ~t[229]);
  assign t[171] = (t[230] & ~t[231]);
  assign t[172] = (t[232] & ~t[233]);
  assign t[173] = (t[234] & ~t[235]);
  assign t[174] = (t[236] & ~t[237]);
  assign t[175] = (t[238] & ~t[239]);
  assign t[176] = t[240] ^ x[2];
  assign t[177] = t[241] ^ x[1];
  assign t[178] = t[242] ^ x[10];
  assign t[179] = t[243] ^ x[9];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[244] ^ x[13];
  assign t[181] = t[245] ^ x[12];
  assign t[182] = t[246] ^ x[16];
  assign t[183] = t[247] ^ x[15];
  assign t[184] = t[248] ^ x[19];
  assign t[185] = t[249] ^ x[18];
  assign t[186] = t[250] ^ x[22];
  assign t[187] = t[251] ^ x[21];
  assign t[188] = t[252] ^ x[25];
  assign t[189] = t[253] ^ x[24];
  assign t[18] = ~(t[24]);
  assign t[190] = t[254] ^ x[30];
  assign t[191] = t[255] ^ x[29];
  assign t[192] = t[256] ^ x[33];
  assign t[193] = t[257] ^ x[32];
  assign t[194] = t[258] ^ x[36];
  assign t[195] = t[259] ^ x[35];
  assign t[196] = t[260] ^ x[41];
  assign t[197] = t[261] ^ x[40];
  assign t[198] = t[262] ^ x[46];
  assign t[199] = t[263] ^ x[45];
  assign t[19] = x[4] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[49];
  assign t[201] = t[265] ^ x[48];
  assign t[202] = t[266] ^ x[52];
  assign t[203] = t[267] ^ x[51];
  assign t[204] = t[268] ^ x[55];
  assign t[205] = t[269] ^ x[54];
  assign t[206] = t[270] ^ x[58];
  assign t[207] = t[271] ^ x[57];
  assign t[208] = t[272] ^ x[61];
  assign t[209] = t[273] ^ x[60];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[274] ^ x[64];
  assign t[211] = t[275] ^ x[63];
  assign t[212] = t[276] ^ x[67];
  assign t[213] = t[277] ^ x[66];
  assign t[214] = t[278] ^ x[70];
  assign t[215] = t[279] ^ x[69];
  assign t[216] = t[280] ^ x[73];
  assign t[217] = t[281] ^ x[72];
  assign t[218] = t[282] ^ x[76];
  assign t[219] = t[283] ^ x[75];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[284] ^ x[79];
  assign t[221] = t[285] ^ x[78];
  assign t[222] = t[286] ^ x[82];
  assign t[223] = t[287] ^ x[81];
  assign t[224] = t[288] ^ x[85];
  assign t[225] = t[289] ^ x[84];
  assign t[226] = t[290] ^ x[88];
  assign t[227] = t[291] ^ x[87];
  assign t[228] = t[292] ^ x[91];
  assign t[229] = t[293] ^ x[90];
  assign t[22] = x[4] ? t[30] : t[29];
  assign t[230] = t[294] ^ x[94];
  assign t[231] = t[295] ^ x[93];
  assign t[232] = t[296] ^ x[97];
  assign t[233] = t[297] ^ x[96];
  assign t[234] = t[298] ^ x[100];
  assign t[235] = t[299] ^ x[99];
  assign t[236] = t[300] ^ x[103];
  assign t[237] = t[301] ^ x[102];
  assign t[238] = t[302] ^ x[106];
  assign t[239] = t[303] ^ x[105];
  assign t[23] = x[4] ? t[32] : t[31];
  assign t[240] = (x[0]);
  assign t[241] = (x[0]);
  assign t[242] = (x[8]);
  assign t[243] = (x[8]);
  assign t[244] = (x[11]);
  assign t[245] = (x[11]);
  assign t[246] = (x[14]);
  assign t[247] = (x[14]);
  assign t[248] = (x[17]);
  assign t[249] = (x[17]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[20]);
  assign t[251] = (x[20]);
  assign t[252] = (x[23]);
  assign t[253] = (x[23]);
  assign t[254] = (x[28]);
  assign t[255] = (x[28]);
  assign t[256] = (x[31]);
  assign t[257] = (x[31]);
  assign t[258] = (x[34]);
  assign t[259] = (x[34]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[39]);
  assign t[261] = (x[39]);
  assign t[262] = (x[44]);
  assign t[263] = (x[44]);
  assign t[264] = (x[47]);
  assign t[265] = (x[47]);
  assign t[266] = (x[50]);
  assign t[267] = (x[50]);
  assign t[268] = (x[53]);
  assign t[269] = (x[53]);
  assign t[26] = t[35] ^ t[36];
  assign t[270] = (x[56]);
  assign t[271] = (x[56]);
  assign t[272] = (x[59]);
  assign t[273] = (x[59]);
  assign t[274] = (x[62]);
  assign t[275] = (x[62]);
  assign t[276] = (x[65]);
  assign t[277] = (x[65]);
  assign t[278] = (x[68]);
  assign t[279] = (x[68]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[280] = (x[71]);
  assign t[281] = (x[71]);
  assign t[282] = (x[74]);
  assign t[283] = (x[74]);
  assign t[284] = (x[77]);
  assign t[285] = (x[77]);
  assign t[286] = (x[80]);
  assign t[287] = (x[80]);
  assign t[288] = (x[83]);
  assign t[289] = (x[83]);
  assign t[28] = t[39] | t[85];
  assign t[290] = (x[86]);
  assign t[291] = (x[86]);
  assign t[292] = (x[89]);
  assign t[293] = (x[89]);
  assign t[294] = (x[92]);
  assign t[295] = (x[92]);
  assign t[296] = (x[95]);
  assign t[297] = (x[95]);
  assign t[298] = (x[98]);
  assign t[299] = (x[98]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[101]);
  assign t[301] = (x[101]);
  assign t[302] = (x[104]);
  assign t[303] = (x[104]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[27] : x[26];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[57] ? x[38] : x[37];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[60] & t[61]);
  assign t[45] = t[62] | t[90];
  assign t[46] = t[57] ? x[43] : x[42];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[70] & t[71]);
  assign t[59] = t[72] | t[96];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[97]);
  assign t[61] = ~(t[98]);
  assign t[62] = ~(t[73] | t[60]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind236(x, y);
 input [151:0] x;
 output y;

 wire [525:0] t;
  assign t[0] = t[1] ? t[2] : t[211];
  assign t[100] = ~(t[234]);
  assign t[101] = ~(t[144] | t[145]);
  assign t[102] = ~(t[146] | t[147]);
  assign t[103] = ~(t[235] | t[148]);
  assign t[104] = t[91] ? x[87] : x[86];
  assign t[105] = ~(t[149] & t[150]);
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[223] | t[224]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151] | t[152]);
  assign t[111] = ~(t[49]);
  assign t[112] = ~(t[137] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[239]);
  assign t[115] = ~(t[240]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = t[111] ? x[104] : x[103];
  assign t[118] = ~(t[158] & t[159]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[160] | t[161]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = ~(t[243] | t[164]);
  assign t[124] = t[111] ? x[115] : x[114];
  assign t[125] = ~(t[84] & t[149]);
  assign t[126] = ~(t[214]);
  assign t[127] = ~(t[165] & t[166]);
  assign t[128] = ~(x[4] & t[167]);
  assign t[129] = ~(t[81] | t[168]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[142] & t[169]);
  assign t[131] = ~(t[126] | t[170]);
  assign t[132] = ~(t[126] | t[171]);
  assign t[133] = ~(t[172] & t[215]);
  assign t[134] = ~(t[173] & t[166]);
  assign t[135] = ~(t[244]);
  assign t[136] = ~(t[229] | t[230]);
  assign t[137] = ~(t[81] | t[174]);
  assign t[138] = t[175] | t[176];
  assign t[139] = ~(t[177] & t[178]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[245]);
  assign t[141] = ~(t[231] | t[232]);
  assign t[142] = ~(t[179] | t[180]);
  assign t[143] = ~(t[181] | t[182]);
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[233] | t[234]);
  assign t[146] = ~(t[247]);
  assign t[147] = ~(t[248]);
  assign t[148] = ~(t[183] | t[184]);
  assign t[149] = ~(t[130] | t[185]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[129] | t[153]);
  assign t[151] = ~(t[249]);
  assign t[152] = ~(t[237] | t[238]);
  assign t[153] = ~(t[81] | t[186]);
  assign t[154] = t[215] & t[187];
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[250]);
  assign t[157] = ~(t[239] | t[240]);
  assign t[158] = ~(t[179] | t[132]);
  assign t[159] = ~(t[188] | t[176]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[241] | t[242]);
  assign t[162] = ~(t[252]);
  assign t[163] = ~(t[253]);
  assign t[164] = ~(t[189] | t[190]);
  assign t[165] = ~(x[4] | t[191]);
  assign t[166] = ~(t[215]);
  assign t[167] = ~(t[213] | t[166]);
  assign t[168] = t[212] ? t[133] : t[134];
  assign t[169] = ~(t[126] & t[192]);
  assign t[16] = ~(t[212] & t[213]);
  assign t[170] = t[212] ? t[193] : t[134];
  assign t[171] = t[212] ? t[127] : t[194];
  assign t[172] = x[4] & t[213];
  assign t[173] = ~(x[4] | t[213]);
  assign t[174] = t[212] ? t[194] : t[195];
  assign t[175] = ~(t[84] & t[196]);
  assign t[176] = ~(t[81] | t[197]);
  assign t[177] = ~(t[198] | t[50]);
  assign t[178] = t[126] | t[199];
  assign t[179] = ~(t[126] | t[200]);
  assign t[17] = ~(t[214] & t[215]);
  assign t[180] = ~(t[81] | t[201]);
  assign t[181] = ~(t[81] | t[202]);
  assign t[182] = ~(t[150] & t[178]);
  assign t[183] = ~(t[254]);
  assign t[184] = ~(t[247] | t[248]);
  assign t[185] = ~(t[203] & t[178]);
  assign t[186] = t[212] ? t[193] : t[204];
  assign t[187] = ~(t[126] | t[212]);
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[255]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[252] | t[253]);
  assign t[191] = ~(t[213]);
  assign t[192] = ~(t[194] & t[195]);
  assign t[193] = ~(t[172] & t[166]);
  assign t[194] = ~(x[4] & t[206]);
  assign t[195] = ~(t[215] & t[165]);
  assign t[196] = ~(t[167] & t[207]);
  assign t[197] = t[212] ? t[195] : t[194];
  assign t[198] = ~(t[208]);
  assign t[199] = t[212] ? t[194] : t[127];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[212] ? t[134] : t[193];
  assign t[201] = t[212] ? t[127] : t[128];
  assign t[202] = t[212] ? t[204] : t[193];
  assign t[203] = ~(t[154] & t[209]);
  assign t[204] = ~(t[173] & t[215]);
  assign t[205] = ~(t[50] | t[153]);
  assign t[206] = ~(t[213] | t[215]);
  assign t[207] = t[81] & t[212];
  assign t[208] = ~(t[187] & t[210]);
  assign t[209] = t[173] | t[172];
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = ~(t[195] & t[128]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = t[301] ^ x[2];
  assign t[257] = t[302] ^ x[10];
  assign t[258] = t[303] ^ x[13];
  assign t[259] = t[304] ^ x[16];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[19];
  assign t[261] = t[306] ^ x[22];
  assign t[262] = t[307] ^ x[25];
  assign t[263] = t[308] ^ x[28];
  assign t[264] = t[309] ^ x[31];
  assign t[265] = t[310] ^ x[34];
  assign t[266] = t[311] ^ x[39];
  assign t[267] = t[312] ^ x[42];
  assign t[268] = t[313] ^ x[45];
  assign t[269] = t[314] ^ x[48];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[51];
  assign t[271] = t[316] ^ x[56];
  assign t[272] = t[317] ^ x[59];
  assign t[273] = t[318] ^ x[62];
  assign t[274] = t[319] ^ x[65];
  assign t[275] = t[320] ^ x[68];
  assign t[276] = t[321] ^ x[71];
  assign t[277] = t[322] ^ x[74];
  assign t[278] = t[323] ^ x[79];
  assign t[279] = t[324] ^ x[82];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[85];
  assign t[281] = t[326] ^ x[90];
  assign t[282] = t[327] ^ x[93];
  assign t[283] = t[328] ^ x[96];
  assign t[284] = t[329] ^ x[99];
  assign t[285] = t[330] ^ x[102];
  assign t[286] = t[331] ^ x[107];
  assign t[287] = t[332] ^ x[110];
  assign t[288] = t[333] ^ x[113];
  assign t[289] = t[334] ^ x[118];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[121];
  assign t[291] = t[336] ^ x[124];
  assign t[292] = t[337] ^ x[127];
  assign t[293] = t[338] ^ x[130];
  assign t[294] = t[339] ^ x[133];
  assign t[295] = t[340] ^ x[136];
  assign t[296] = t[341] ^ x[139];
  assign t[297] = t[342] ^ x[142];
  assign t[298] = t[343] ^ x[145];
  assign t[299] = t[344] ^ x[148];
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[151];
  assign t[301] = (t[346] & ~t[347]);
  assign t[302] = (t[348] & ~t[349]);
  assign t[303] = (t[350] & ~t[351]);
  assign t[304] = (t[352] & ~t[353]);
  assign t[305] = (t[354] & ~t[355]);
  assign t[306] = (t[356] & ~t[357]);
  assign t[307] = (t[358] & ~t[359]);
  assign t[308] = (t[360] & ~t[361]);
  assign t[309] = (t[362] & ~t[363]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[364] & ~t[365]);
  assign t[311] = (t[366] & ~t[367]);
  assign t[312] = (t[368] & ~t[369]);
  assign t[313] = (t[370] & ~t[371]);
  assign t[314] = (t[372] & ~t[373]);
  assign t[315] = (t[374] & ~t[375]);
  assign t[316] = (t[376] & ~t[377]);
  assign t[317] = (t[378] & ~t[379]);
  assign t[318] = (t[380] & ~t[381]);
  assign t[319] = (t[382] & ~t[383]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[384] & ~t[385]);
  assign t[321] = (t[386] & ~t[387]);
  assign t[322] = (t[388] & ~t[389]);
  assign t[323] = (t[390] & ~t[391]);
  assign t[324] = (t[392] & ~t[393]);
  assign t[325] = (t[394] & ~t[395]);
  assign t[326] = (t[396] & ~t[397]);
  assign t[327] = (t[398] & ~t[399]);
  assign t[328] = (t[400] & ~t[401]);
  assign t[329] = (t[402] & ~t[403]);
  assign t[32] = ~(t[52]);
  assign t[330] = (t[404] & ~t[405]);
  assign t[331] = (t[406] & ~t[407]);
  assign t[332] = (t[408] & ~t[409]);
  assign t[333] = (t[410] & ~t[411]);
  assign t[334] = (t[412] & ~t[413]);
  assign t[335] = (t[414] & ~t[415]);
  assign t[336] = (t[416] & ~t[417]);
  assign t[337] = (t[418] & ~t[419]);
  assign t[338] = (t[420] & ~t[421]);
  assign t[339] = (t[422] & ~t[423]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = (t[424] & ~t[425]);
  assign t[341] = (t[426] & ~t[427]);
  assign t[342] = (t[428] & ~t[429]);
  assign t[343] = (t[430] & ~t[431]);
  assign t[344] = (t[432] & ~t[433]);
  assign t[345] = (t[434] & ~t[435]);
  assign t[346] = t[436] ^ x[2];
  assign t[347] = t[437] ^ x[1];
  assign t[348] = t[438] ^ x[10];
  assign t[349] = t[439] ^ x[9];
  assign t[34] = ~(t[216] | t[55]);
  assign t[350] = t[440] ^ x[13];
  assign t[351] = t[441] ^ x[12];
  assign t[352] = t[442] ^ x[16];
  assign t[353] = t[443] ^ x[15];
  assign t[354] = t[444] ^ x[19];
  assign t[355] = t[445] ^ x[18];
  assign t[356] = t[446] ^ x[22];
  assign t[357] = t[447] ^ x[21];
  assign t[358] = t[448] ^ x[25];
  assign t[359] = t[449] ^ x[24];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[450] ^ x[28];
  assign t[361] = t[451] ^ x[27];
  assign t[362] = t[452] ^ x[31];
  assign t[363] = t[453] ^ x[30];
  assign t[364] = t[454] ^ x[34];
  assign t[365] = t[455] ^ x[33];
  assign t[366] = t[456] ^ x[39];
  assign t[367] = t[457] ^ x[38];
  assign t[368] = t[458] ^ x[42];
  assign t[369] = t[459] ^ x[41];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[460] ^ x[45];
  assign t[371] = t[461] ^ x[44];
  assign t[372] = t[462] ^ x[48];
  assign t[373] = t[463] ^ x[47];
  assign t[374] = t[464] ^ x[51];
  assign t[375] = t[465] ^ x[50];
  assign t[376] = t[466] ^ x[56];
  assign t[377] = t[467] ^ x[55];
  assign t[378] = t[468] ^ x[59];
  assign t[379] = t[469] ^ x[58];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[470] ^ x[62];
  assign t[381] = t[471] ^ x[61];
  assign t[382] = t[472] ^ x[65];
  assign t[383] = t[473] ^ x[64];
  assign t[384] = t[474] ^ x[68];
  assign t[385] = t[475] ^ x[67];
  assign t[386] = t[476] ^ x[71];
  assign t[387] = t[477] ^ x[70];
  assign t[388] = t[478] ^ x[74];
  assign t[389] = t[479] ^ x[73];
  assign t[38] = ~(t[47] ^ t[62]);
  assign t[390] = t[480] ^ x[79];
  assign t[391] = t[481] ^ x[78];
  assign t[392] = t[482] ^ x[82];
  assign t[393] = t[483] ^ x[81];
  assign t[394] = t[484] ^ x[85];
  assign t[395] = t[485] ^ x[84];
  assign t[396] = t[486] ^ x[90];
  assign t[397] = t[487] ^ x[89];
  assign t[398] = t[488] ^ x[93];
  assign t[399] = t[489] ^ x[92];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[96];
  assign t[401] = t[491] ^ x[95];
  assign t[402] = t[492] ^ x[99];
  assign t[403] = t[493] ^ x[98];
  assign t[404] = t[494] ^ x[102];
  assign t[405] = t[495] ^ x[101];
  assign t[406] = t[496] ^ x[107];
  assign t[407] = t[497] ^ x[106];
  assign t[408] = t[498] ^ x[110];
  assign t[409] = t[499] ^ x[109];
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[410] = t[500] ^ x[113];
  assign t[411] = t[501] ^ x[112];
  assign t[412] = t[502] ^ x[118];
  assign t[413] = t[503] ^ x[117];
  assign t[414] = t[504] ^ x[121];
  assign t[415] = t[505] ^ x[120];
  assign t[416] = t[506] ^ x[124];
  assign t[417] = t[507] ^ x[123];
  assign t[418] = t[508] ^ x[127];
  assign t[419] = t[509] ^ x[126];
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = t[510] ^ x[130];
  assign t[421] = t[511] ^ x[129];
  assign t[422] = t[512] ^ x[133];
  assign t[423] = t[513] ^ x[132];
  assign t[424] = t[514] ^ x[136];
  assign t[425] = t[515] ^ x[135];
  assign t[426] = t[516] ^ x[139];
  assign t[427] = t[517] ^ x[138];
  assign t[428] = t[518] ^ x[142];
  assign t[429] = t[519] ^ x[141];
  assign t[42] = ~(t[217] | t[69]);
  assign t[430] = t[520] ^ x[145];
  assign t[431] = t[521] ^ x[144];
  assign t[432] = t[522] ^ x[148];
  assign t[433] = t[523] ^ x[147];
  assign t[434] = t[524] ^ x[151];
  assign t[435] = t[525] ^ x[150];
  assign t[436] = (x[0]);
  assign t[437] = (x[0]);
  assign t[438] = (x[8]);
  assign t[439] = (x[8]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[11]);
  assign t[441] = (x[11]);
  assign t[442] = (x[14]);
  assign t[443] = (x[14]);
  assign t[444] = (x[17]);
  assign t[445] = (x[17]);
  assign t[446] = (x[20]);
  assign t[447] = (x[20]);
  assign t[448] = (x[23]);
  assign t[449] = (x[23]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[26]);
  assign t[451] = (x[26]);
  assign t[452] = (x[29]);
  assign t[453] = (x[29]);
  assign t[454] = (x[32]);
  assign t[455] = (x[32]);
  assign t[456] = (x[37]);
  assign t[457] = (x[37]);
  assign t[458] = (x[40]);
  assign t[459] = (x[40]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[43]);
  assign t[461] = (x[43]);
  assign t[462] = (x[46]);
  assign t[463] = (x[46]);
  assign t[464] = (x[49]);
  assign t[465] = (x[49]);
  assign t[466] = (x[54]);
  assign t[467] = (x[54]);
  assign t[468] = (x[57]);
  assign t[469] = (x[57]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = (x[60]);
  assign t[471] = (x[60]);
  assign t[472] = (x[63]);
  assign t[473] = (x[63]);
  assign t[474] = (x[66]);
  assign t[475] = (x[66]);
  assign t[476] = (x[69]);
  assign t[477] = (x[69]);
  assign t[478] = (x[72]);
  assign t[479] = (x[72]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[77]);
  assign t[481] = (x[77]);
  assign t[482] = (x[80]);
  assign t[483] = (x[80]);
  assign t[484] = (x[83]);
  assign t[485] = (x[83]);
  assign t[486] = (x[88]);
  assign t[487] = (x[88]);
  assign t[488] = (x[91]);
  assign t[489] = (x[91]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = (x[94]);
  assign t[491] = (x[94]);
  assign t[492] = (x[97]);
  assign t[493] = (x[97]);
  assign t[494] = (x[100]);
  assign t[495] = (x[100]);
  assign t[496] = (x[105]);
  assign t[497] = (x[105]);
  assign t[498] = (x[108]);
  assign t[499] = (x[108]);
  assign t[49] = ~(t[214]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[111]);
  assign t[501] = (x[111]);
  assign t[502] = (x[116]);
  assign t[503] = (x[116]);
  assign t[504] = (x[119]);
  assign t[505] = (x[119]);
  assign t[506] = (x[122]);
  assign t[507] = (x[122]);
  assign t[508] = (x[125]);
  assign t[509] = (x[125]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (x[128]);
  assign t[511] = (x[128]);
  assign t[512] = (x[131]);
  assign t[513] = (x[131]);
  assign t[514] = (x[134]);
  assign t[515] = (x[134]);
  assign t[516] = (x[137]);
  assign t[517] = (x[137]);
  assign t[518] = (x[140]);
  assign t[519] = (x[140]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[520] = (x[143]);
  assign t[521] = (x[143]);
  assign t[522] = (x[146]);
  assign t[523] = (x[146]);
  assign t[524] = (x[149]);
  assign t[525] = (x[149]);
  assign t[52] = ~(t[81] | t[85]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[220] | t[90]);
  assign t[58] = t[91] ? x[36] : x[35];
  assign t[59] = ~(t[92] & t[93]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[221] | t[96]);
  assign t[62] = ~(t[97] ^ t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[222] | t[101]);
  assign t[65] = ~(t[102] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[223]);
  assign t[68] = ~(t[224]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[225] | t[110]);
  assign t[72] = t[111] ? x[53] : x[52];
  assign t[73] = ~(t[112] & t[113]);
  assign t[74] = ~(t[114] | t[115]);
  assign t[75] = ~(t[226] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[227] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[212] ? t[128] : t[127];
  assign t[83] = ~(t[129] | t[130]);
  assign t[84] = ~(t[131] | t[132]);
  assign t[85] = t[212] ? t[134] : t[133];
  assign t[86] = ~(t[228]);
  assign t[87] = ~(t[218] | t[219]);
  assign t[88] = ~(t[229]);
  assign t[89] = ~(t[230]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[135] | t[136]);
  assign t[91] = ~(t[49]);
  assign t[92] = ~(t[129] | t[137]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[231]);
  assign t[95] = ~(t[232]);
  assign t[96] = ~(t[140] | t[141]);
  assign t[97] = t[91] ? x[76] : x[75];
  assign t[98] = ~(t[142] & t[143]);
  assign t[99] = ~(t[233]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [151:0] x;
 output y;

 wire [525:0] t;
  assign t[0] = t[1] ? t[2] : t[211];
  assign t[100] = ~(t[234]);
  assign t[101] = ~(t[144] | t[145]);
  assign t[102] = ~(t[146] | t[147]);
  assign t[103] = ~(t[235] | t[148]);
  assign t[104] = t[91] ? x[87] : x[86];
  assign t[105] = ~(t[149] & t[150]);
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[223] | t[224]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151] | t[152]);
  assign t[111] = ~(t[49]);
  assign t[112] = ~(t[137] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[239]);
  assign t[115] = ~(t[240]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = t[111] ? x[104] : x[103];
  assign t[118] = ~(t[158] & t[159]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[160] | t[161]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = ~(t[243] | t[164]);
  assign t[124] = t[111] ? x[115] : x[114];
  assign t[125] = ~(t[84] & t[149]);
  assign t[126] = ~(t[214]);
  assign t[127] = ~(t[165] & t[166]);
  assign t[128] = ~(x[4] & t[167]);
  assign t[129] = ~(t[81] | t[168]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[142] & t[169]);
  assign t[131] = ~(t[126] | t[170]);
  assign t[132] = ~(t[126] | t[171]);
  assign t[133] = ~(t[172] & t[215]);
  assign t[134] = ~(t[173] & t[166]);
  assign t[135] = ~(t[244]);
  assign t[136] = ~(t[229] | t[230]);
  assign t[137] = ~(t[81] | t[174]);
  assign t[138] = t[175] | t[176];
  assign t[139] = ~(t[177] & t[178]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[245]);
  assign t[141] = ~(t[231] | t[232]);
  assign t[142] = ~(t[179] | t[180]);
  assign t[143] = ~(t[181] | t[182]);
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[233] | t[234]);
  assign t[146] = ~(t[247]);
  assign t[147] = ~(t[248]);
  assign t[148] = ~(t[183] | t[184]);
  assign t[149] = ~(t[130] | t[185]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[129] | t[153]);
  assign t[151] = ~(t[249]);
  assign t[152] = ~(t[237] | t[238]);
  assign t[153] = ~(t[81] | t[186]);
  assign t[154] = t[215] & t[187];
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[250]);
  assign t[157] = ~(t[239] | t[240]);
  assign t[158] = ~(t[179] | t[132]);
  assign t[159] = ~(t[188] | t[176]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[241] | t[242]);
  assign t[162] = ~(t[252]);
  assign t[163] = ~(t[253]);
  assign t[164] = ~(t[189] | t[190]);
  assign t[165] = ~(x[4] | t[191]);
  assign t[166] = ~(t[215]);
  assign t[167] = ~(t[213] | t[166]);
  assign t[168] = t[212] ? t[133] : t[134];
  assign t[169] = ~(t[126] & t[192]);
  assign t[16] = ~(t[212] & t[213]);
  assign t[170] = t[212] ? t[193] : t[134];
  assign t[171] = t[212] ? t[127] : t[194];
  assign t[172] = x[4] & t[213];
  assign t[173] = ~(x[4] | t[213]);
  assign t[174] = t[212] ? t[194] : t[195];
  assign t[175] = ~(t[84] & t[196]);
  assign t[176] = ~(t[81] | t[197]);
  assign t[177] = ~(t[198] | t[50]);
  assign t[178] = t[126] | t[199];
  assign t[179] = ~(t[126] | t[200]);
  assign t[17] = ~(t[214] & t[215]);
  assign t[180] = ~(t[81] | t[201]);
  assign t[181] = ~(t[81] | t[202]);
  assign t[182] = ~(t[150] & t[178]);
  assign t[183] = ~(t[254]);
  assign t[184] = ~(t[247] | t[248]);
  assign t[185] = ~(t[203] & t[178]);
  assign t[186] = t[212] ? t[193] : t[204];
  assign t[187] = ~(t[126] | t[212]);
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[255]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[252] | t[253]);
  assign t[191] = ~(t[213]);
  assign t[192] = ~(t[194] & t[195]);
  assign t[193] = ~(t[172] & t[166]);
  assign t[194] = ~(x[4] & t[206]);
  assign t[195] = ~(t[215] & t[165]);
  assign t[196] = ~(t[167] & t[207]);
  assign t[197] = t[212] ? t[195] : t[194];
  assign t[198] = ~(t[208]);
  assign t[199] = t[212] ? t[194] : t[127];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[212] ? t[134] : t[193];
  assign t[201] = t[212] ? t[127] : t[128];
  assign t[202] = t[212] ? t[204] : t[193];
  assign t[203] = ~(t[154] & t[209]);
  assign t[204] = ~(t[173] & t[215]);
  assign t[205] = ~(t[50] | t[153]);
  assign t[206] = ~(t[213] | t[215]);
  assign t[207] = t[81] & t[212];
  assign t[208] = ~(t[187] & t[210]);
  assign t[209] = t[173] | t[172];
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = ~(t[195] & t[128]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = t[301] ^ x[2];
  assign t[257] = t[302] ^ x[10];
  assign t[258] = t[303] ^ x[13];
  assign t[259] = t[304] ^ x[16];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[19];
  assign t[261] = t[306] ^ x[22];
  assign t[262] = t[307] ^ x[25];
  assign t[263] = t[308] ^ x[28];
  assign t[264] = t[309] ^ x[31];
  assign t[265] = t[310] ^ x[34];
  assign t[266] = t[311] ^ x[39];
  assign t[267] = t[312] ^ x[42];
  assign t[268] = t[313] ^ x[45];
  assign t[269] = t[314] ^ x[48];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[51];
  assign t[271] = t[316] ^ x[56];
  assign t[272] = t[317] ^ x[59];
  assign t[273] = t[318] ^ x[62];
  assign t[274] = t[319] ^ x[65];
  assign t[275] = t[320] ^ x[68];
  assign t[276] = t[321] ^ x[71];
  assign t[277] = t[322] ^ x[74];
  assign t[278] = t[323] ^ x[79];
  assign t[279] = t[324] ^ x[82];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[85];
  assign t[281] = t[326] ^ x[90];
  assign t[282] = t[327] ^ x[93];
  assign t[283] = t[328] ^ x[96];
  assign t[284] = t[329] ^ x[99];
  assign t[285] = t[330] ^ x[102];
  assign t[286] = t[331] ^ x[107];
  assign t[287] = t[332] ^ x[110];
  assign t[288] = t[333] ^ x[113];
  assign t[289] = t[334] ^ x[118];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[121];
  assign t[291] = t[336] ^ x[124];
  assign t[292] = t[337] ^ x[127];
  assign t[293] = t[338] ^ x[130];
  assign t[294] = t[339] ^ x[133];
  assign t[295] = t[340] ^ x[136];
  assign t[296] = t[341] ^ x[139];
  assign t[297] = t[342] ^ x[142];
  assign t[298] = t[343] ^ x[145];
  assign t[299] = t[344] ^ x[148];
  assign t[29] = x[4] ? t[48] : t[47];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[151];
  assign t[301] = (t[346] & ~t[347]);
  assign t[302] = (t[348] & ~t[349]);
  assign t[303] = (t[350] & ~t[351]);
  assign t[304] = (t[352] & ~t[353]);
  assign t[305] = (t[354] & ~t[355]);
  assign t[306] = (t[356] & ~t[357]);
  assign t[307] = (t[358] & ~t[359]);
  assign t[308] = (t[360] & ~t[361]);
  assign t[309] = (t[362] & ~t[363]);
  assign t[30] = ~(t[49]);
  assign t[310] = (t[364] & ~t[365]);
  assign t[311] = (t[366] & ~t[367]);
  assign t[312] = (t[368] & ~t[369]);
  assign t[313] = (t[370] & ~t[371]);
  assign t[314] = (t[372] & ~t[373]);
  assign t[315] = (t[374] & ~t[375]);
  assign t[316] = (t[376] & ~t[377]);
  assign t[317] = (t[378] & ~t[379]);
  assign t[318] = (t[380] & ~t[381]);
  assign t[319] = (t[382] & ~t[383]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (t[384] & ~t[385]);
  assign t[321] = (t[386] & ~t[387]);
  assign t[322] = (t[388] & ~t[389]);
  assign t[323] = (t[390] & ~t[391]);
  assign t[324] = (t[392] & ~t[393]);
  assign t[325] = (t[394] & ~t[395]);
  assign t[326] = (t[396] & ~t[397]);
  assign t[327] = (t[398] & ~t[399]);
  assign t[328] = (t[400] & ~t[401]);
  assign t[329] = (t[402] & ~t[403]);
  assign t[32] = ~(t[52]);
  assign t[330] = (t[404] & ~t[405]);
  assign t[331] = (t[406] & ~t[407]);
  assign t[332] = (t[408] & ~t[409]);
  assign t[333] = (t[410] & ~t[411]);
  assign t[334] = (t[412] & ~t[413]);
  assign t[335] = (t[414] & ~t[415]);
  assign t[336] = (t[416] & ~t[417]);
  assign t[337] = (t[418] & ~t[419]);
  assign t[338] = (t[420] & ~t[421]);
  assign t[339] = (t[422] & ~t[423]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = (t[424] & ~t[425]);
  assign t[341] = (t[426] & ~t[427]);
  assign t[342] = (t[428] & ~t[429]);
  assign t[343] = (t[430] & ~t[431]);
  assign t[344] = (t[432] & ~t[433]);
  assign t[345] = (t[434] & ~t[435]);
  assign t[346] = t[436] ^ x[2];
  assign t[347] = t[437] ^ x[1];
  assign t[348] = t[438] ^ x[10];
  assign t[349] = t[439] ^ x[9];
  assign t[34] = ~(t[216] | t[55]);
  assign t[350] = t[440] ^ x[13];
  assign t[351] = t[441] ^ x[12];
  assign t[352] = t[442] ^ x[16];
  assign t[353] = t[443] ^ x[15];
  assign t[354] = t[444] ^ x[19];
  assign t[355] = t[445] ^ x[18];
  assign t[356] = t[446] ^ x[22];
  assign t[357] = t[447] ^ x[21];
  assign t[358] = t[448] ^ x[25];
  assign t[359] = t[449] ^ x[24];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[450] ^ x[28];
  assign t[361] = t[451] ^ x[27];
  assign t[362] = t[452] ^ x[31];
  assign t[363] = t[453] ^ x[30];
  assign t[364] = t[454] ^ x[34];
  assign t[365] = t[455] ^ x[33];
  assign t[366] = t[456] ^ x[39];
  assign t[367] = t[457] ^ x[38];
  assign t[368] = t[458] ^ x[42];
  assign t[369] = t[459] ^ x[41];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[460] ^ x[45];
  assign t[371] = t[461] ^ x[44];
  assign t[372] = t[462] ^ x[48];
  assign t[373] = t[463] ^ x[47];
  assign t[374] = t[464] ^ x[51];
  assign t[375] = t[465] ^ x[50];
  assign t[376] = t[466] ^ x[56];
  assign t[377] = t[467] ^ x[55];
  assign t[378] = t[468] ^ x[59];
  assign t[379] = t[469] ^ x[58];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[470] ^ x[62];
  assign t[381] = t[471] ^ x[61];
  assign t[382] = t[472] ^ x[65];
  assign t[383] = t[473] ^ x[64];
  assign t[384] = t[474] ^ x[68];
  assign t[385] = t[475] ^ x[67];
  assign t[386] = t[476] ^ x[71];
  assign t[387] = t[477] ^ x[70];
  assign t[388] = t[478] ^ x[74];
  assign t[389] = t[479] ^ x[73];
  assign t[38] = ~(t[47] ^ t[62]);
  assign t[390] = t[480] ^ x[79];
  assign t[391] = t[481] ^ x[78];
  assign t[392] = t[482] ^ x[82];
  assign t[393] = t[483] ^ x[81];
  assign t[394] = t[484] ^ x[85];
  assign t[395] = t[485] ^ x[84];
  assign t[396] = t[486] ^ x[90];
  assign t[397] = t[487] ^ x[89];
  assign t[398] = t[488] ^ x[93];
  assign t[399] = t[489] ^ x[92];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[490] ^ x[96];
  assign t[401] = t[491] ^ x[95];
  assign t[402] = t[492] ^ x[99];
  assign t[403] = t[493] ^ x[98];
  assign t[404] = t[494] ^ x[102];
  assign t[405] = t[495] ^ x[101];
  assign t[406] = t[496] ^ x[107];
  assign t[407] = t[497] ^ x[106];
  assign t[408] = t[498] ^ x[110];
  assign t[409] = t[499] ^ x[109];
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[410] = t[500] ^ x[113];
  assign t[411] = t[501] ^ x[112];
  assign t[412] = t[502] ^ x[118];
  assign t[413] = t[503] ^ x[117];
  assign t[414] = t[504] ^ x[121];
  assign t[415] = t[505] ^ x[120];
  assign t[416] = t[506] ^ x[124];
  assign t[417] = t[507] ^ x[123];
  assign t[418] = t[508] ^ x[127];
  assign t[419] = t[509] ^ x[126];
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = t[510] ^ x[130];
  assign t[421] = t[511] ^ x[129];
  assign t[422] = t[512] ^ x[133];
  assign t[423] = t[513] ^ x[132];
  assign t[424] = t[514] ^ x[136];
  assign t[425] = t[515] ^ x[135];
  assign t[426] = t[516] ^ x[139];
  assign t[427] = t[517] ^ x[138];
  assign t[428] = t[518] ^ x[142];
  assign t[429] = t[519] ^ x[141];
  assign t[42] = ~(t[217] | t[69]);
  assign t[430] = t[520] ^ x[145];
  assign t[431] = t[521] ^ x[144];
  assign t[432] = t[522] ^ x[148];
  assign t[433] = t[523] ^ x[147];
  assign t[434] = t[524] ^ x[151];
  assign t[435] = t[525] ^ x[150];
  assign t[436] = (x[0]);
  assign t[437] = (x[0]);
  assign t[438] = (x[8]);
  assign t[439] = (x[8]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[11]);
  assign t[441] = (x[11]);
  assign t[442] = (x[14]);
  assign t[443] = (x[14]);
  assign t[444] = (x[17]);
  assign t[445] = (x[17]);
  assign t[446] = (x[20]);
  assign t[447] = (x[20]);
  assign t[448] = (x[23]);
  assign t[449] = (x[23]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[26]);
  assign t[451] = (x[26]);
  assign t[452] = (x[29]);
  assign t[453] = (x[29]);
  assign t[454] = (x[32]);
  assign t[455] = (x[32]);
  assign t[456] = (x[37]);
  assign t[457] = (x[37]);
  assign t[458] = (x[40]);
  assign t[459] = (x[40]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[43]);
  assign t[461] = (x[43]);
  assign t[462] = (x[46]);
  assign t[463] = (x[46]);
  assign t[464] = (x[49]);
  assign t[465] = (x[49]);
  assign t[466] = (x[54]);
  assign t[467] = (x[54]);
  assign t[468] = (x[57]);
  assign t[469] = (x[57]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = (x[60]);
  assign t[471] = (x[60]);
  assign t[472] = (x[63]);
  assign t[473] = (x[63]);
  assign t[474] = (x[66]);
  assign t[475] = (x[66]);
  assign t[476] = (x[69]);
  assign t[477] = (x[69]);
  assign t[478] = (x[72]);
  assign t[479] = (x[72]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (x[77]);
  assign t[481] = (x[77]);
  assign t[482] = (x[80]);
  assign t[483] = (x[80]);
  assign t[484] = (x[83]);
  assign t[485] = (x[83]);
  assign t[486] = (x[88]);
  assign t[487] = (x[88]);
  assign t[488] = (x[91]);
  assign t[489] = (x[91]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = (x[94]);
  assign t[491] = (x[94]);
  assign t[492] = (x[97]);
  assign t[493] = (x[97]);
  assign t[494] = (x[100]);
  assign t[495] = (x[100]);
  assign t[496] = (x[105]);
  assign t[497] = (x[105]);
  assign t[498] = (x[108]);
  assign t[499] = (x[108]);
  assign t[49] = ~(t[214]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[500] = (x[111]);
  assign t[501] = (x[111]);
  assign t[502] = (x[116]);
  assign t[503] = (x[116]);
  assign t[504] = (x[119]);
  assign t[505] = (x[119]);
  assign t[506] = (x[122]);
  assign t[507] = (x[122]);
  assign t[508] = (x[125]);
  assign t[509] = (x[125]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (x[128]);
  assign t[511] = (x[128]);
  assign t[512] = (x[131]);
  assign t[513] = (x[131]);
  assign t[514] = (x[134]);
  assign t[515] = (x[134]);
  assign t[516] = (x[137]);
  assign t[517] = (x[137]);
  assign t[518] = (x[140]);
  assign t[519] = (x[140]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[520] = (x[143]);
  assign t[521] = (x[143]);
  assign t[522] = (x[146]);
  assign t[523] = (x[146]);
  assign t[524] = (x[149]);
  assign t[525] = (x[149]);
  assign t[52] = ~(t[81] | t[85]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[220] | t[90]);
  assign t[58] = t[91] ? x[36] : x[35];
  assign t[59] = ~(t[92] & t[93]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[221] | t[96]);
  assign t[62] = ~(t[97] ^ t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[222] | t[101]);
  assign t[65] = ~(t[102] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[223]);
  assign t[68] = ~(t[224]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[225] | t[110]);
  assign t[72] = t[111] ? x[53] : x[52];
  assign t[73] = ~(t[112] & t[113]);
  assign t[74] = ~(t[114] | t[115]);
  assign t[75] = ~(t[226] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[227] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[212] ? t[128] : t[127];
  assign t[83] = ~(t[129] | t[130]);
  assign t[84] = ~(t[131] | t[132]);
  assign t[85] = t[212] ? t[134] : t[133];
  assign t[86] = ~(t[228]);
  assign t[87] = ~(t[218] | t[219]);
  assign t[88] = ~(t[229]);
  assign t[89] = ~(t[230]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[135] | t[136]);
  assign t[91] = ~(t[49]);
  assign t[92] = ~(t[129] | t[137]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[231]);
  assign t[95] = ~(t[232]);
  assign t[96] = ~(t[140] | t[141]);
  assign t[97] = t[91] ? x[76] : x[75];
  assign t[98] = ~(t[142] & t[143]);
  assign t[99] = ~(t[233]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[42];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ? x[35] : x[34];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[44];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[60] ? x[52] : x[51];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[48] ? x[60] : x[59];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[25]);
  assign t[61] = ~(t[117] & t[80]);
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[60] ? x[77] : x[76];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[121] & t[86]);
  assign t[68] = ~(t[122] & t[87]);
  assign t[69] = t[60] ? x[85] : x[84];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131] & t[96]);
  assign t[86] = ~(t[132]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[134]);
  assign t[96] = ~(t[134] & t[99]);
  assign t[97] = ~(t[121]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[130]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [121:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[2];
  assign t[136] = t[171] ^ x[10];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[16];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[22];
  assign t[141] = t[176] ^ x[25];
  assign t[142] = t[177] ^ x[30];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[38];
  assign t[145] = t[180] ^ x[41];
  assign t[146] = t[181] ^ x[44];
  assign t[147] = t[182] ^ x[47];
  assign t[148] = t[183] ^ x[50];
  assign t[149] = t[184] ^ x[55];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[58];
  assign t[151] = t[186] ^ x[63];
  assign t[152] = t[187] ^ x[66];
  assign t[153] = t[188] ^ x[69];
  assign t[154] = t[189] ^ x[72];
  assign t[155] = t[190] ^ x[75];
  assign t[156] = t[191] ^ x[80];
  assign t[157] = t[192] ^ x[83];
  assign t[158] = t[193] ^ x[88];
  assign t[159] = t[194] ^ x[91];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[94];
  assign t[161] = t[196] ^ x[97];
  assign t[162] = t[197] ^ x[100];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[106];
  assign t[165] = t[200] ^ x[109];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[115];
  assign t[168] = t[203] ^ x[118];
  assign t[169] = t[204] ^ x[121];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (t[205] & ~t[206]);
  assign t[171] = (t[207] & ~t[208]);
  assign t[172] = (t[209] & ~t[210]);
  assign t[173] = (t[211] & ~t[212]);
  assign t[174] = (t[213] & ~t[214]);
  assign t[175] = (t[215] & ~t[216]);
  assign t[176] = (t[217] & ~t[218]);
  assign t[177] = (t[219] & ~t[220]);
  assign t[178] = (t[221] & ~t[222]);
  assign t[179] = (t[223] & ~t[224]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (t[225] & ~t[226]);
  assign t[181] = (t[227] & ~t[228]);
  assign t[182] = (t[229] & ~t[230]);
  assign t[183] = (t[231] & ~t[232]);
  assign t[184] = (t[233] & ~t[234]);
  assign t[185] = (t[235] & ~t[236]);
  assign t[186] = (t[237] & ~t[238]);
  assign t[187] = (t[239] & ~t[240]);
  assign t[188] = (t[241] & ~t[242]);
  assign t[189] = (t[243] & ~t[244]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[245] & ~t[246]);
  assign t[191] = (t[247] & ~t[248]);
  assign t[192] = (t[249] & ~t[250]);
  assign t[193] = (t[251] & ~t[252]);
  assign t[194] = (t[253] & ~t[254]);
  assign t[195] = (t[255] & ~t[256]);
  assign t[196] = (t[257] & ~t[258]);
  assign t[197] = (t[259] & ~t[260]);
  assign t[198] = (t[261] & ~t[262]);
  assign t[199] = (t[263] & ~t[264]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[265] & ~t[266]);
  assign t[201] = (t[267] & ~t[268]);
  assign t[202] = (t[269] & ~t[270]);
  assign t[203] = (t[271] & ~t[272]);
  assign t[204] = (t[273] & ~t[274]);
  assign t[205] = t[275] ^ x[2];
  assign t[206] = t[276] ^ x[1];
  assign t[207] = t[277] ^ x[10];
  assign t[208] = t[278] ^ x[9];
  assign t[209] = t[279] ^ x[13];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[280] ^ x[12];
  assign t[211] = t[281] ^ x[16];
  assign t[212] = t[282] ^ x[15];
  assign t[213] = t[283] ^ x[19];
  assign t[214] = t[284] ^ x[18];
  assign t[215] = t[285] ^ x[22];
  assign t[216] = t[286] ^ x[21];
  assign t[217] = t[287] ^ x[25];
  assign t[218] = t[288] ^ x[24];
  assign t[219] = t[289] ^ x[30];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[290] ^ x[29];
  assign t[221] = t[291] ^ x[33];
  assign t[222] = t[292] ^ x[32];
  assign t[223] = t[293] ^ x[38];
  assign t[224] = t[294] ^ x[37];
  assign t[225] = t[295] ^ x[41];
  assign t[226] = t[296] ^ x[40];
  assign t[227] = t[297] ^ x[44];
  assign t[228] = t[298] ^ x[43];
  assign t[229] = t[299] ^ x[47];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[300] ^ x[46];
  assign t[231] = t[301] ^ x[50];
  assign t[232] = t[302] ^ x[49];
  assign t[233] = t[303] ^ x[55];
  assign t[234] = t[304] ^ x[54];
  assign t[235] = t[305] ^ x[58];
  assign t[236] = t[306] ^ x[57];
  assign t[237] = t[307] ^ x[63];
  assign t[238] = t[308] ^ x[62];
  assign t[239] = t[309] ^ x[66];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[310] ^ x[65];
  assign t[241] = t[311] ^ x[69];
  assign t[242] = t[312] ^ x[68];
  assign t[243] = t[313] ^ x[72];
  assign t[244] = t[314] ^ x[71];
  assign t[245] = t[315] ^ x[75];
  assign t[246] = t[316] ^ x[74];
  assign t[247] = t[317] ^ x[80];
  assign t[248] = t[318] ^ x[79];
  assign t[249] = t[319] ^ x[83];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[320] ^ x[82];
  assign t[251] = t[321] ^ x[88];
  assign t[252] = t[322] ^ x[87];
  assign t[253] = t[323] ^ x[91];
  assign t[254] = t[324] ^ x[90];
  assign t[255] = t[325] ^ x[94];
  assign t[256] = t[326] ^ x[93];
  assign t[257] = t[327] ^ x[97];
  assign t[258] = t[328] ^ x[96];
  assign t[259] = t[329] ^ x[100];
  assign t[25] = ~(t[103]);
  assign t[260] = t[330] ^ x[99];
  assign t[261] = t[331] ^ x[103];
  assign t[262] = t[332] ^ x[102];
  assign t[263] = t[333] ^ x[106];
  assign t[264] = t[334] ^ x[105];
  assign t[265] = t[335] ^ x[109];
  assign t[266] = t[336] ^ x[108];
  assign t[267] = t[337] ^ x[112];
  assign t[268] = t[338] ^ x[111];
  assign t[269] = t[339] ^ x[115];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[340] ^ x[114];
  assign t[271] = t[341] ^ x[118];
  assign t[272] = t[342] ^ x[117];
  assign t[273] = t[343] ^ x[121];
  assign t[274] = t[344] ^ x[120];
  assign t[275] = (x[0]);
  assign t[276] = (x[0]);
  assign t[277] = (x[8]);
  assign t[278] = (x[8]);
  assign t[279] = (x[11]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[11]);
  assign t[281] = (x[14]);
  assign t[282] = (x[14]);
  assign t[283] = (x[17]);
  assign t[284] = (x[17]);
  assign t[285] = (x[20]);
  assign t[286] = (x[20]);
  assign t[287] = (x[23]);
  assign t[288] = (x[23]);
  assign t[289] = (x[28]);
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = (x[28]);
  assign t[291] = (x[31]);
  assign t[292] = (x[31]);
  assign t[293] = (x[36]);
  assign t[294] = (x[36]);
  assign t[295] = (x[39]);
  assign t[296] = (x[39]);
  assign t[297] = (x[42]);
  assign t[298] = (x[42]);
  assign t[299] = (x[45]);
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[45]);
  assign t[301] = (x[48]);
  assign t[302] = (x[48]);
  assign t[303] = (x[53]);
  assign t[304] = (x[53]);
  assign t[305] = (x[56]);
  assign t[306] = (x[56]);
  assign t[307] = (x[61]);
  assign t[308] = (x[61]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[310] = (x[64]);
  assign t[311] = (x[67]);
  assign t[312] = (x[67]);
  assign t[313] = (x[70]);
  assign t[314] = (x[70]);
  assign t[315] = (x[73]);
  assign t[316] = (x[73]);
  assign t[317] = (x[78]);
  assign t[318] = (x[78]);
  assign t[319] = (x[81]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[320] = (x[81]);
  assign t[321] = (x[86]);
  assign t[322] = (x[86]);
  assign t[323] = (x[89]);
  assign t[324] = (x[89]);
  assign t[325] = (x[92]);
  assign t[326] = (x[92]);
  assign t[327] = (x[95]);
  assign t[328] = (x[95]);
  assign t[329] = (x[98]);
  assign t[32] = t[48] ? x[27] : x[26];
  assign t[330] = (x[98]);
  assign t[331] = (x[101]);
  assign t[332] = (x[101]);
  assign t[333] = (x[104]);
  assign t[334] = (x[104]);
  assign t[335] = (x[107]);
  assign t[336] = (x[107]);
  assign t[337] = (x[110]);
  assign t[338] = (x[110]);
  assign t[339] = (x[113]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[113]);
  assign t[341] = (x[116]);
  assign t[342] = (x[116]);
  assign t[343] = (x[119]);
  assign t[344] = (x[119]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[42];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ? x[35] : x[34];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[44];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[60] ? x[52] : x[51];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[48] ? x[60] : x[59];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[25]);
  assign t[61] = ~(t[117] & t[80]);
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[60] ? x[77] : x[76];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[121] & t[86]);
  assign t[68] = ~(t[122] & t[87]);
  assign t[69] = t[60] ? x[85] : x[84];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131] & t[96]);
  assign t[86] = ~(t[132]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[134]);
  assign t[96] = ~(t[134] & t[99]);
  assign t[97] = ~(t[121]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[130]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [151:0] x;
 output y;

 wire [434:0] t;
  assign t[0] = t[1] ? t[2] : t[120];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[156]);
  assign t[104] = ~(t[116] & t[117]);
  assign t[105] = ~(t[144] & t[143]);
  assign t[106] = ~(t[157]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[151] & t[150]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[162]);
  assign t[115] = ~(t[118] & t[119]);
  assign t[116] = ~(t[156] & t[155]);
  assign t[117] = ~(t[163]);
  assign t[118] = ~(t[162] & t[161]);
  assign t[119] = ~(t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = (t[209]);
  assign t[165] = t[210] ^ x[2];
  assign t[166] = t[211] ^ x[10];
  assign t[167] = t[212] ^ x[13];
  assign t[168] = t[213] ^ x[16];
  assign t[169] = t[214] ^ x[19];
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = t[215] ^ x[22];
  assign t[171] = t[216] ^ x[27];
  assign t[172] = t[217] ^ x[32];
  assign t[173] = t[218] ^ x[35];
  assign t[174] = t[219] ^ x[38];
  assign t[175] = t[220] ^ x[41];
  assign t[176] = t[221] ^ x[46];
  assign t[177] = t[222] ^ x[51];
  assign t[178] = t[223] ^ x[54];
  assign t[179] = t[224] ^ x[57];
  assign t[17] = ~(t[123] & t[124]);
  assign t[180] = t[225] ^ x[60];
  assign t[181] = t[226] ^ x[65];
  assign t[182] = t[227] ^ x[70];
  assign t[183] = t[228] ^ x[73];
  assign t[184] = t[229] ^ x[76];
  assign t[185] = t[230] ^ x[79];
  assign t[186] = t[231] ^ x[82];
  assign t[187] = t[232] ^ x[85];
  assign t[188] = t[233] ^ x[88];
  assign t[189] = t[234] ^ x[91];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[94];
  assign t[191] = t[236] ^ x[97];
  assign t[192] = t[237] ^ x[100];
  assign t[193] = t[238] ^ x[103];
  assign t[194] = t[239] ^ x[106];
  assign t[195] = t[240] ^ x[109];
  assign t[196] = t[241] ^ x[112];
  assign t[197] = t[242] ^ x[115];
  assign t[198] = t[243] ^ x[118];
  assign t[199] = t[244] ^ x[121];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[124];
  assign t[201] = t[246] ^ x[127];
  assign t[202] = t[247] ^ x[130];
  assign t[203] = t[248] ^ x[133];
  assign t[204] = t[249] ^ x[136];
  assign t[205] = t[250] ^ x[139];
  assign t[206] = t[251] ^ x[142];
  assign t[207] = t[252] ^ x[145];
  assign t[208] = t[253] ^ x[148];
  assign t[209] = t[254] ^ x[151];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[255] & ~t[256]);
  assign t[211] = (t[257] & ~t[258]);
  assign t[212] = (t[259] & ~t[260]);
  assign t[213] = (t[261] & ~t[262]);
  assign t[214] = (t[263] & ~t[264]);
  assign t[215] = (t[265] & ~t[266]);
  assign t[216] = (t[267] & ~t[268]);
  assign t[217] = (t[269] & ~t[270]);
  assign t[218] = (t[271] & ~t[272]);
  assign t[219] = (t[273] & ~t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[275] & ~t[276]);
  assign t[221] = (t[277] & ~t[278]);
  assign t[222] = (t[279] & ~t[280]);
  assign t[223] = (t[281] & ~t[282]);
  assign t[224] = (t[283] & ~t[284]);
  assign t[225] = (t[285] & ~t[286]);
  assign t[226] = (t[287] & ~t[288]);
  assign t[227] = (t[289] & ~t[290]);
  assign t[228] = (t[291] & ~t[292]);
  assign t[229] = (t[293] & ~t[294]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[295] & ~t[296]);
  assign t[231] = (t[297] & ~t[298]);
  assign t[232] = (t[299] & ~t[300]);
  assign t[233] = (t[301] & ~t[302]);
  assign t[234] = (t[303] & ~t[304]);
  assign t[235] = (t[305] & ~t[306]);
  assign t[236] = (t[307] & ~t[308]);
  assign t[237] = (t[309] & ~t[310]);
  assign t[238] = (t[311] & ~t[312]);
  assign t[239] = (t[313] & ~t[314]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[315] & ~t[316]);
  assign t[241] = (t[317] & ~t[318]);
  assign t[242] = (t[319] & ~t[320]);
  assign t[243] = (t[321] & ~t[322]);
  assign t[244] = (t[323] & ~t[324]);
  assign t[245] = (t[325] & ~t[326]);
  assign t[246] = (t[327] & ~t[328]);
  assign t[247] = (t[329] & ~t[330]);
  assign t[248] = (t[331] & ~t[332]);
  assign t[249] = (t[333] & ~t[334]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[335] & ~t[336]);
  assign t[251] = (t[337] & ~t[338]);
  assign t[252] = (t[339] & ~t[340]);
  assign t[253] = (t[341] & ~t[342]);
  assign t[254] = (t[343] & ~t[344]);
  assign t[255] = t[345] ^ x[2];
  assign t[256] = t[346] ^ x[1];
  assign t[257] = t[347] ^ x[10];
  assign t[258] = t[348] ^ x[9];
  assign t[259] = t[349] ^ x[13];
  assign t[25] = ~(t[123]);
  assign t[260] = t[350] ^ x[12];
  assign t[261] = t[351] ^ x[16];
  assign t[262] = t[352] ^ x[15];
  assign t[263] = t[353] ^ x[19];
  assign t[264] = t[354] ^ x[18];
  assign t[265] = t[355] ^ x[22];
  assign t[266] = t[356] ^ x[21];
  assign t[267] = t[357] ^ x[27];
  assign t[268] = t[358] ^ x[26];
  assign t[269] = t[359] ^ x[32];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[31];
  assign t[271] = t[361] ^ x[35];
  assign t[272] = t[362] ^ x[34];
  assign t[273] = t[363] ^ x[38];
  assign t[274] = t[364] ^ x[37];
  assign t[275] = t[365] ^ x[41];
  assign t[276] = t[366] ^ x[40];
  assign t[277] = t[367] ^ x[46];
  assign t[278] = t[368] ^ x[45];
  assign t[279] = t[369] ^ x[51];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[50];
  assign t[281] = t[371] ^ x[54];
  assign t[282] = t[372] ^ x[53];
  assign t[283] = t[373] ^ x[57];
  assign t[284] = t[374] ^ x[56];
  assign t[285] = t[375] ^ x[60];
  assign t[286] = t[376] ^ x[59];
  assign t[287] = t[377] ^ x[65];
  assign t[288] = t[378] ^ x[64];
  assign t[289] = t[379] ^ x[70];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[69];
  assign t[291] = t[381] ^ x[73];
  assign t[292] = t[382] ^ x[72];
  assign t[293] = t[383] ^ x[76];
  assign t[294] = t[384] ^ x[75];
  assign t[295] = t[385] ^ x[79];
  assign t[296] = t[386] ^ x[78];
  assign t[297] = t[387] ^ x[82];
  assign t[298] = t[388] ^ x[81];
  assign t[299] = t[389] ^ x[85];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[84];
  assign t[301] = t[391] ^ x[88];
  assign t[302] = t[392] ^ x[87];
  assign t[303] = t[393] ^ x[91];
  assign t[304] = t[394] ^ x[90];
  assign t[305] = t[395] ^ x[94];
  assign t[306] = t[396] ^ x[93];
  assign t[307] = t[397] ^ x[97];
  assign t[308] = t[398] ^ x[96];
  assign t[309] = t[399] ^ x[100];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[99];
  assign t[311] = t[401] ^ x[103];
  assign t[312] = t[402] ^ x[102];
  assign t[313] = t[403] ^ x[106];
  assign t[314] = t[404] ^ x[105];
  assign t[315] = t[405] ^ x[109];
  assign t[316] = t[406] ^ x[108];
  assign t[317] = t[407] ^ x[112];
  assign t[318] = t[408] ^ x[111];
  assign t[319] = t[409] ^ x[115];
  assign t[31] = ~(t[48] & t[125]);
  assign t[320] = t[410] ^ x[114];
  assign t[321] = t[411] ^ x[118];
  assign t[322] = t[412] ^ x[117];
  assign t[323] = t[413] ^ x[121];
  assign t[324] = t[414] ^ x[120];
  assign t[325] = t[415] ^ x[124];
  assign t[326] = t[416] ^ x[123];
  assign t[327] = t[417] ^ x[127];
  assign t[328] = t[418] ^ x[126];
  assign t[329] = t[419] ^ x[130];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[129];
  assign t[331] = t[421] ^ x[133];
  assign t[332] = t[422] ^ x[132];
  assign t[333] = t[423] ^ x[136];
  assign t[334] = t[424] ^ x[135];
  assign t[335] = t[425] ^ x[139];
  assign t[336] = t[426] ^ x[138];
  assign t[337] = t[427] ^ x[142];
  assign t[338] = t[428] ^ x[141];
  assign t[339] = t[429] ^ x[145];
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = t[430] ^ x[144];
  assign t[341] = t[431] ^ x[148];
  assign t[342] = t[432] ^ x[147];
  assign t[343] = t[433] ^ x[151];
  assign t[344] = t[434] ^ x[150];
  assign t[345] = (x[0]);
  assign t[346] = (x[0]);
  assign t[347] = (x[8]);
  assign t[348] = (x[8]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[11]);
  assign t[351] = (x[14]);
  assign t[352] = (x[14]);
  assign t[353] = (x[17]);
  assign t[354] = (x[17]);
  assign t[355] = (x[20]);
  assign t[356] = (x[20]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[30]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[30]);
  assign t[361] = (x[33]);
  assign t[362] = (x[33]);
  assign t[363] = (x[36]);
  assign t[364] = (x[36]);
  assign t[365] = (x[39]);
  assign t[366] = (x[39]);
  assign t[367] = (x[44]);
  assign t[368] = (x[44]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[49]);
  assign t[371] = (x[52]);
  assign t[372] = (x[52]);
  assign t[373] = (x[55]);
  assign t[374] = (x[55]);
  assign t[375] = (x[58]);
  assign t[376] = (x[58]);
  assign t[377] = (x[63]);
  assign t[378] = (x[63]);
  assign t[379] = (x[68]);
  assign t[37] = t[58] ^ t[44];
  assign t[380] = (x[68]);
  assign t[381] = (x[71]);
  assign t[382] = (x[71]);
  assign t[383] = (x[74]);
  assign t[384] = (x[74]);
  assign t[385] = (x[77]);
  assign t[386] = (x[77]);
  assign t[387] = (x[80]);
  assign t[388] = (x[80]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[83]);
  assign t[391] = (x[86]);
  assign t[392] = (x[86]);
  assign t[393] = (x[89]);
  assign t[394] = (x[89]);
  assign t[395] = (x[92]);
  assign t[396] = (x[92]);
  assign t[397] = (x[95]);
  assign t[398] = (x[95]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[61] & t[126]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[98]);
  assign t[401] = (x[101]);
  assign t[402] = (x[101]);
  assign t[403] = (x[104]);
  assign t[404] = (x[104]);
  assign t[405] = (x[107]);
  assign t[406] = (x[107]);
  assign t[407] = (x[110]);
  assign t[408] = (x[110]);
  assign t[409] = (x[113]);
  assign t[40] = t[62] ? x[29] : x[28];
  assign t[410] = (x[113]);
  assign t[411] = (x[116]);
  assign t[412] = (x[116]);
  assign t[413] = (x[119]);
  assign t[414] = (x[119]);
  assign t[415] = (x[122]);
  assign t[416] = (x[122]);
  assign t[417] = (x[125]);
  assign t[418] = (x[125]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[420] = (x[128]);
  assign t[421] = (x[131]);
  assign t[422] = (x[131]);
  assign t[423] = (x[134]);
  assign t[424] = (x[134]);
  assign t[425] = (x[137]);
  assign t[426] = (x[137]);
  assign t[427] = (x[140]);
  assign t[428] = (x[140]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[430] = (x[143]);
  assign t[431] = (x[146]);
  assign t[432] = (x[146]);
  assign t[433] = (x[149]);
  assign t[434] = (x[149]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[127]);
  assign t[47] = ~(t[128]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[129]);
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[130]);
  assign t[54] = t[49] ? x[43] : x[42];
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = ~(t[82] & t[83]);
  assign t[57] = ~(t[84] & t[131]);
  assign t[58] = t[18] ? x[48] : x[47];
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[133]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[134]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[135]);
  assign t[67] = t[62] ? x[62] : x[61];
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = ~(t[95] & t[136]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[67] : x[66];
  assign t[71] = ~(t[96] & t[97]);
  assign t[72] = ~(t[128] & t[127]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[98] & t[99]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[102] & t[103]);
  assign t[81] = ~(t[104] & t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[105] & t[106]);
  assign t[85] = ~(t[133] & t[132]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[147]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[109] & t[110]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[151]);
  assign t[95] = ~(t[111] & t[112]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[115] & t[152]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[153]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind241(x, y);
 input [151:0] x;
 output y;

 wire [434:0] t;
  assign t[0] = t[1] ? t[2] : t[120];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[156]);
  assign t[104] = ~(t[116] & t[117]);
  assign t[105] = ~(t[144] & t[143]);
  assign t[106] = ~(t[157]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[151] & t[150]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[162]);
  assign t[115] = ~(t[118] & t[119]);
  assign t[116] = ~(t[156] & t[155]);
  assign t[117] = ~(t[163]);
  assign t[118] = ~(t[162] & t[161]);
  assign t[119] = ~(t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = (t[209]);
  assign t[165] = t[210] ^ x[2];
  assign t[166] = t[211] ^ x[10];
  assign t[167] = t[212] ^ x[13];
  assign t[168] = t[213] ^ x[16];
  assign t[169] = t[214] ^ x[19];
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = t[215] ^ x[22];
  assign t[171] = t[216] ^ x[27];
  assign t[172] = t[217] ^ x[32];
  assign t[173] = t[218] ^ x[35];
  assign t[174] = t[219] ^ x[38];
  assign t[175] = t[220] ^ x[41];
  assign t[176] = t[221] ^ x[46];
  assign t[177] = t[222] ^ x[51];
  assign t[178] = t[223] ^ x[54];
  assign t[179] = t[224] ^ x[57];
  assign t[17] = ~(t[123] & t[124]);
  assign t[180] = t[225] ^ x[60];
  assign t[181] = t[226] ^ x[65];
  assign t[182] = t[227] ^ x[70];
  assign t[183] = t[228] ^ x[73];
  assign t[184] = t[229] ^ x[76];
  assign t[185] = t[230] ^ x[79];
  assign t[186] = t[231] ^ x[82];
  assign t[187] = t[232] ^ x[85];
  assign t[188] = t[233] ^ x[88];
  assign t[189] = t[234] ^ x[91];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[94];
  assign t[191] = t[236] ^ x[97];
  assign t[192] = t[237] ^ x[100];
  assign t[193] = t[238] ^ x[103];
  assign t[194] = t[239] ^ x[106];
  assign t[195] = t[240] ^ x[109];
  assign t[196] = t[241] ^ x[112];
  assign t[197] = t[242] ^ x[115];
  assign t[198] = t[243] ^ x[118];
  assign t[199] = t[244] ^ x[121];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[124];
  assign t[201] = t[246] ^ x[127];
  assign t[202] = t[247] ^ x[130];
  assign t[203] = t[248] ^ x[133];
  assign t[204] = t[249] ^ x[136];
  assign t[205] = t[250] ^ x[139];
  assign t[206] = t[251] ^ x[142];
  assign t[207] = t[252] ^ x[145];
  assign t[208] = t[253] ^ x[148];
  assign t[209] = t[254] ^ x[151];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[255] & ~t[256]);
  assign t[211] = (t[257] & ~t[258]);
  assign t[212] = (t[259] & ~t[260]);
  assign t[213] = (t[261] & ~t[262]);
  assign t[214] = (t[263] & ~t[264]);
  assign t[215] = (t[265] & ~t[266]);
  assign t[216] = (t[267] & ~t[268]);
  assign t[217] = (t[269] & ~t[270]);
  assign t[218] = (t[271] & ~t[272]);
  assign t[219] = (t[273] & ~t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[275] & ~t[276]);
  assign t[221] = (t[277] & ~t[278]);
  assign t[222] = (t[279] & ~t[280]);
  assign t[223] = (t[281] & ~t[282]);
  assign t[224] = (t[283] & ~t[284]);
  assign t[225] = (t[285] & ~t[286]);
  assign t[226] = (t[287] & ~t[288]);
  assign t[227] = (t[289] & ~t[290]);
  assign t[228] = (t[291] & ~t[292]);
  assign t[229] = (t[293] & ~t[294]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[295] & ~t[296]);
  assign t[231] = (t[297] & ~t[298]);
  assign t[232] = (t[299] & ~t[300]);
  assign t[233] = (t[301] & ~t[302]);
  assign t[234] = (t[303] & ~t[304]);
  assign t[235] = (t[305] & ~t[306]);
  assign t[236] = (t[307] & ~t[308]);
  assign t[237] = (t[309] & ~t[310]);
  assign t[238] = (t[311] & ~t[312]);
  assign t[239] = (t[313] & ~t[314]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[315] & ~t[316]);
  assign t[241] = (t[317] & ~t[318]);
  assign t[242] = (t[319] & ~t[320]);
  assign t[243] = (t[321] & ~t[322]);
  assign t[244] = (t[323] & ~t[324]);
  assign t[245] = (t[325] & ~t[326]);
  assign t[246] = (t[327] & ~t[328]);
  assign t[247] = (t[329] & ~t[330]);
  assign t[248] = (t[331] & ~t[332]);
  assign t[249] = (t[333] & ~t[334]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (t[335] & ~t[336]);
  assign t[251] = (t[337] & ~t[338]);
  assign t[252] = (t[339] & ~t[340]);
  assign t[253] = (t[341] & ~t[342]);
  assign t[254] = (t[343] & ~t[344]);
  assign t[255] = t[345] ^ x[2];
  assign t[256] = t[346] ^ x[1];
  assign t[257] = t[347] ^ x[10];
  assign t[258] = t[348] ^ x[9];
  assign t[259] = t[349] ^ x[13];
  assign t[25] = ~(t[123]);
  assign t[260] = t[350] ^ x[12];
  assign t[261] = t[351] ^ x[16];
  assign t[262] = t[352] ^ x[15];
  assign t[263] = t[353] ^ x[19];
  assign t[264] = t[354] ^ x[18];
  assign t[265] = t[355] ^ x[22];
  assign t[266] = t[356] ^ x[21];
  assign t[267] = t[357] ^ x[27];
  assign t[268] = t[358] ^ x[26];
  assign t[269] = t[359] ^ x[32];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[31];
  assign t[271] = t[361] ^ x[35];
  assign t[272] = t[362] ^ x[34];
  assign t[273] = t[363] ^ x[38];
  assign t[274] = t[364] ^ x[37];
  assign t[275] = t[365] ^ x[41];
  assign t[276] = t[366] ^ x[40];
  assign t[277] = t[367] ^ x[46];
  assign t[278] = t[368] ^ x[45];
  assign t[279] = t[369] ^ x[51];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[50];
  assign t[281] = t[371] ^ x[54];
  assign t[282] = t[372] ^ x[53];
  assign t[283] = t[373] ^ x[57];
  assign t[284] = t[374] ^ x[56];
  assign t[285] = t[375] ^ x[60];
  assign t[286] = t[376] ^ x[59];
  assign t[287] = t[377] ^ x[65];
  assign t[288] = t[378] ^ x[64];
  assign t[289] = t[379] ^ x[70];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[69];
  assign t[291] = t[381] ^ x[73];
  assign t[292] = t[382] ^ x[72];
  assign t[293] = t[383] ^ x[76];
  assign t[294] = t[384] ^ x[75];
  assign t[295] = t[385] ^ x[79];
  assign t[296] = t[386] ^ x[78];
  assign t[297] = t[387] ^ x[82];
  assign t[298] = t[388] ^ x[81];
  assign t[299] = t[389] ^ x[85];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[84];
  assign t[301] = t[391] ^ x[88];
  assign t[302] = t[392] ^ x[87];
  assign t[303] = t[393] ^ x[91];
  assign t[304] = t[394] ^ x[90];
  assign t[305] = t[395] ^ x[94];
  assign t[306] = t[396] ^ x[93];
  assign t[307] = t[397] ^ x[97];
  assign t[308] = t[398] ^ x[96];
  assign t[309] = t[399] ^ x[100];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[99];
  assign t[311] = t[401] ^ x[103];
  assign t[312] = t[402] ^ x[102];
  assign t[313] = t[403] ^ x[106];
  assign t[314] = t[404] ^ x[105];
  assign t[315] = t[405] ^ x[109];
  assign t[316] = t[406] ^ x[108];
  assign t[317] = t[407] ^ x[112];
  assign t[318] = t[408] ^ x[111];
  assign t[319] = t[409] ^ x[115];
  assign t[31] = ~(t[48] & t[125]);
  assign t[320] = t[410] ^ x[114];
  assign t[321] = t[411] ^ x[118];
  assign t[322] = t[412] ^ x[117];
  assign t[323] = t[413] ^ x[121];
  assign t[324] = t[414] ^ x[120];
  assign t[325] = t[415] ^ x[124];
  assign t[326] = t[416] ^ x[123];
  assign t[327] = t[417] ^ x[127];
  assign t[328] = t[418] ^ x[126];
  assign t[329] = t[419] ^ x[130];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[129];
  assign t[331] = t[421] ^ x[133];
  assign t[332] = t[422] ^ x[132];
  assign t[333] = t[423] ^ x[136];
  assign t[334] = t[424] ^ x[135];
  assign t[335] = t[425] ^ x[139];
  assign t[336] = t[426] ^ x[138];
  assign t[337] = t[427] ^ x[142];
  assign t[338] = t[428] ^ x[141];
  assign t[339] = t[429] ^ x[145];
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = t[430] ^ x[144];
  assign t[341] = t[431] ^ x[148];
  assign t[342] = t[432] ^ x[147];
  assign t[343] = t[433] ^ x[151];
  assign t[344] = t[434] ^ x[150];
  assign t[345] = (x[0]);
  assign t[346] = (x[0]);
  assign t[347] = (x[8]);
  assign t[348] = (x[8]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[11]);
  assign t[351] = (x[14]);
  assign t[352] = (x[14]);
  assign t[353] = (x[17]);
  assign t[354] = (x[17]);
  assign t[355] = (x[20]);
  assign t[356] = (x[20]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[30]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[30]);
  assign t[361] = (x[33]);
  assign t[362] = (x[33]);
  assign t[363] = (x[36]);
  assign t[364] = (x[36]);
  assign t[365] = (x[39]);
  assign t[366] = (x[39]);
  assign t[367] = (x[44]);
  assign t[368] = (x[44]);
  assign t[369] = (x[49]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[49]);
  assign t[371] = (x[52]);
  assign t[372] = (x[52]);
  assign t[373] = (x[55]);
  assign t[374] = (x[55]);
  assign t[375] = (x[58]);
  assign t[376] = (x[58]);
  assign t[377] = (x[63]);
  assign t[378] = (x[63]);
  assign t[379] = (x[68]);
  assign t[37] = t[58] ^ t[44];
  assign t[380] = (x[68]);
  assign t[381] = (x[71]);
  assign t[382] = (x[71]);
  assign t[383] = (x[74]);
  assign t[384] = (x[74]);
  assign t[385] = (x[77]);
  assign t[386] = (x[77]);
  assign t[387] = (x[80]);
  assign t[388] = (x[80]);
  assign t[389] = (x[83]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[83]);
  assign t[391] = (x[86]);
  assign t[392] = (x[86]);
  assign t[393] = (x[89]);
  assign t[394] = (x[89]);
  assign t[395] = (x[92]);
  assign t[396] = (x[92]);
  assign t[397] = (x[95]);
  assign t[398] = (x[95]);
  assign t[399] = (x[98]);
  assign t[39] = ~(t[61] & t[126]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[98]);
  assign t[401] = (x[101]);
  assign t[402] = (x[101]);
  assign t[403] = (x[104]);
  assign t[404] = (x[104]);
  assign t[405] = (x[107]);
  assign t[406] = (x[107]);
  assign t[407] = (x[110]);
  assign t[408] = (x[110]);
  assign t[409] = (x[113]);
  assign t[40] = t[62] ? x[29] : x[28];
  assign t[410] = (x[113]);
  assign t[411] = (x[116]);
  assign t[412] = (x[116]);
  assign t[413] = (x[119]);
  assign t[414] = (x[119]);
  assign t[415] = (x[122]);
  assign t[416] = (x[122]);
  assign t[417] = (x[125]);
  assign t[418] = (x[125]);
  assign t[419] = (x[128]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[420] = (x[128]);
  assign t[421] = (x[131]);
  assign t[422] = (x[131]);
  assign t[423] = (x[134]);
  assign t[424] = (x[134]);
  assign t[425] = (x[137]);
  assign t[426] = (x[137]);
  assign t[427] = (x[140]);
  assign t[428] = (x[140]);
  assign t[429] = (x[143]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[430] = (x[143]);
  assign t[431] = (x[146]);
  assign t[432] = (x[146]);
  assign t[433] = (x[149]);
  assign t[434] = (x[149]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[127]);
  assign t[47] = ~(t[128]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[129]);
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[130]);
  assign t[54] = t[49] ? x[43] : x[42];
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = ~(t[82] & t[83]);
  assign t[57] = ~(t[84] & t[131]);
  assign t[58] = t[18] ? x[48] : x[47];
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[133]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[134]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[135]);
  assign t[67] = t[62] ? x[62] : x[61];
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = ~(t[95] & t[136]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[67] : x[66];
  assign t[71] = ~(t[96] & t[97]);
  assign t[72] = ~(t[128] & t[127]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[98] & t[99]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[102] & t[103]);
  assign t[81] = ~(t[104] & t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[105] & t[106]);
  assign t[85] = ~(t[133] & t[132]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[147]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[109] & t[110]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[151]);
  assign t[95] = ~(t[111] & t[112]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[115] & t[152]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[153]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[58] ^ t[44];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[62] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[72] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = t[75] | t[119];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[120];
  assign t[54] = t[49] ? x[43] : x[42];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = t[83] | t[121];
  assign t[58] = t[62] ? x[48] : x[47];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[84] | t[59]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[124];
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = t[90] | t[125];
  assign t[67] = t[62] ? x[62] : x[61];
  assign t[68] = ~(t[91] & t[92]);
  assign t[69] = t[93] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[67] : x[66];
  assign t[71] = ~(t[94] & t[95]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[96] | t[73]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[97] | t[76]);
  assign t[79] = ~(t[98] & t[99]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[100] | t[132];
  assign t[81] = ~(t[133]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[101] | t[81]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [151:0] x;
 output y;

 wire [424:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[2];
  assign t[156] = t[201] ^ x[10];
  assign t[157] = t[202] ^ x[13];
  assign t[158] = t[203] ^ x[16];
  assign t[159] = t[204] ^ x[19];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[22];
  assign t[161] = t[206] ^ x[27];
  assign t[162] = t[207] ^ x[32];
  assign t[163] = t[208] ^ x[35];
  assign t[164] = t[209] ^ x[38];
  assign t[165] = t[210] ^ x[41];
  assign t[166] = t[211] ^ x[46];
  assign t[167] = t[212] ^ x[51];
  assign t[168] = t[213] ^ x[54];
  assign t[169] = t[214] ^ x[57];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[60];
  assign t[171] = t[216] ^ x[65];
  assign t[172] = t[217] ^ x[70];
  assign t[173] = t[218] ^ x[73];
  assign t[174] = t[219] ^ x[76];
  assign t[175] = t[220] ^ x[79];
  assign t[176] = t[221] ^ x[82];
  assign t[177] = t[222] ^ x[85];
  assign t[178] = t[223] ^ x[88];
  assign t[179] = t[224] ^ x[91];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[94];
  assign t[181] = t[226] ^ x[97];
  assign t[182] = t[227] ^ x[100];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[106];
  assign t[185] = t[230] ^ x[109];
  assign t[186] = t[231] ^ x[112];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[118];
  assign t[189] = t[234] ^ x[121];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[124];
  assign t[191] = t[236] ^ x[127];
  assign t[192] = t[237] ^ x[130];
  assign t[193] = t[238] ^ x[133];
  assign t[194] = t[239] ^ x[136];
  assign t[195] = t[240] ^ x[139];
  assign t[196] = t[241] ^ x[142];
  assign t[197] = t[242] ^ x[145];
  assign t[198] = t[243] ^ x[148];
  assign t[199] = t[244] ^ x[151];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[245] & ~t[246]);
  assign t[201] = (t[247] & ~t[248]);
  assign t[202] = (t[249] & ~t[250]);
  assign t[203] = (t[251] & ~t[252]);
  assign t[204] = (t[253] & ~t[254]);
  assign t[205] = (t[255] & ~t[256]);
  assign t[206] = (t[257] & ~t[258]);
  assign t[207] = (t[259] & ~t[260]);
  assign t[208] = (t[261] & ~t[262]);
  assign t[209] = (t[263] & ~t[264]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[265] & ~t[266]);
  assign t[211] = (t[267] & ~t[268]);
  assign t[212] = (t[269] & ~t[270]);
  assign t[213] = (t[271] & ~t[272]);
  assign t[214] = (t[273] & ~t[274]);
  assign t[215] = (t[275] & ~t[276]);
  assign t[216] = (t[277] & ~t[278]);
  assign t[217] = (t[279] & ~t[280]);
  assign t[218] = (t[281] & ~t[282]);
  assign t[219] = (t[283] & ~t[284]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[285] & ~t[286]);
  assign t[221] = (t[287] & ~t[288]);
  assign t[222] = (t[289] & ~t[290]);
  assign t[223] = (t[291] & ~t[292]);
  assign t[224] = (t[293] & ~t[294]);
  assign t[225] = (t[295] & ~t[296]);
  assign t[226] = (t[297] & ~t[298]);
  assign t[227] = (t[299] & ~t[300]);
  assign t[228] = (t[301] & ~t[302]);
  assign t[229] = (t[303] & ~t[304]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[305] & ~t[306]);
  assign t[231] = (t[307] & ~t[308]);
  assign t[232] = (t[309] & ~t[310]);
  assign t[233] = (t[311] & ~t[312]);
  assign t[234] = (t[313] & ~t[314]);
  assign t[235] = (t[315] & ~t[316]);
  assign t[236] = (t[317] & ~t[318]);
  assign t[237] = (t[319] & ~t[320]);
  assign t[238] = (t[321] & ~t[322]);
  assign t[239] = (t[323] & ~t[324]);
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = (t[325] & ~t[326]);
  assign t[241] = (t[327] & ~t[328]);
  assign t[242] = (t[329] & ~t[330]);
  assign t[243] = (t[331] & ~t[332]);
  assign t[244] = (t[333] & ~t[334]);
  assign t[245] = t[335] ^ x[2];
  assign t[246] = t[336] ^ x[1];
  assign t[247] = t[337] ^ x[10];
  assign t[248] = t[338] ^ x[9];
  assign t[249] = t[339] ^ x[13];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[340] ^ x[12];
  assign t[251] = t[341] ^ x[16];
  assign t[252] = t[342] ^ x[15];
  assign t[253] = t[343] ^ x[19];
  assign t[254] = t[344] ^ x[18];
  assign t[255] = t[345] ^ x[22];
  assign t[256] = t[346] ^ x[21];
  assign t[257] = t[347] ^ x[27];
  assign t[258] = t[348] ^ x[26];
  assign t[259] = t[349] ^ x[32];
  assign t[25] = ~(t[113]);
  assign t[260] = t[350] ^ x[31];
  assign t[261] = t[351] ^ x[35];
  assign t[262] = t[352] ^ x[34];
  assign t[263] = t[353] ^ x[38];
  assign t[264] = t[354] ^ x[37];
  assign t[265] = t[355] ^ x[41];
  assign t[266] = t[356] ^ x[40];
  assign t[267] = t[357] ^ x[46];
  assign t[268] = t[358] ^ x[45];
  assign t[269] = t[359] ^ x[51];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[360] ^ x[50];
  assign t[271] = t[361] ^ x[54];
  assign t[272] = t[362] ^ x[53];
  assign t[273] = t[363] ^ x[57];
  assign t[274] = t[364] ^ x[56];
  assign t[275] = t[365] ^ x[60];
  assign t[276] = t[366] ^ x[59];
  assign t[277] = t[367] ^ x[65];
  assign t[278] = t[368] ^ x[64];
  assign t[279] = t[369] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[370] ^ x[69];
  assign t[281] = t[371] ^ x[73];
  assign t[282] = t[372] ^ x[72];
  assign t[283] = t[373] ^ x[76];
  assign t[284] = t[374] ^ x[75];
  assign t[285] = t[375] ^ x[79];
  assign t[286] = t[376] ^ x[78];
  assign t[287] = t[377] ^ x[82];
  assign t[288] = t[378] ^ x[81];
  assign t[289] = t[379] ^ x[85];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[290] = t[380] ^ x[84];
  assign t[291] = t[381] ^ x[88];
  assign t[292] = t[382] ^ x[87];
  assign t[293] = t[383] ^ x[91];
  assign t[294] = t[384] ^ x[90];
  assign t[295] = t[385] ^ x[94];
  assign t[296] = t[386] ^ x[93];
  assign t[297] = t[387] ^ x[97];
  assign t[298] = t[388] ^ x[96];
  assign t[299] = t[389] ^ x[100];
  assign t[29] = x[4] ? t[45] : t[44];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[390] ^ x[99];
  assign t[301] = t[391] ^ x[103];
  assign t[302] = t[392] ^ x[102];
  assign t[303] = t[393] ^ x[106];
  assign t[304] = t[394] ^ x[105];
  assign t[305] = t[395] ^ x[109];
  assign t[306] = t[396] ^ x[108];
  assign t[307] = t[397] ^ x[112];
  assign t[308] = t[398] ^ x[111];
  assign t[309] = t[399] ^ x[115];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[400] ^ x[114];
  assign t[311] = t[401] ^ x[118];
  assign t[312] = t[402] ^ x[117];
  assign t[313] = t[403] ^ x[121];
  assign t[314] = t[404] ^ x[120];
  assign t[315] = t[405] ^ x[124];
  assign t[316] = t[406] ^ x[123];
  assign t[317] = t[407] ^ x[127];
  assign t[318] = t[408] ^ x[126];
  assign t[319] = t[409] ^ x[130];
  assign t[31] = t[48] | t[115];
  assign t[320] = t[410] ^ x[129];
  assign t[321] = t[411] ^ x[133];
  assign t[322] = t[412] ^ x[132];
  assign t[323] = t[413] ^ x[136];
  assign t[324] = t[414] ^ x[135];
  assign t[325] = t[415] ^ x[139];
  assign t[326] = t[416] ^ x[138];
  assign t[327] = t[417] ^ x[142];
  assign t[328] = t[418] ^ x[141];
  assign t[329] = t[419] ^ x[145];
  assign t[32] = t[49] ? x[24] : x[23];
  assign t[330] = t[420] ^ x[144];
  assign t[331] = t[421] ^ x[148];
  assign t[332] = t[422] ^ x[147];
  assign t[333] = t[423] ^ x[151];
  assign t[334] = t[424] ^ x[150];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[8]);
  assign t[338] = (x[8]);
  assign t[339] = (x[11]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[11]);
  assign t[341] = (x[14]);
  assign t[342] = (x[14]);
  assign t[343] = (x[17]);
  assign t[344] = (x[17]);
  assign t[345] = (x[20]);
  assign t[346] = (x[20]);
  assign t[347] = (x[25]);
  assign t[348] = (x[25]);
  assign t[349] = (x[30]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[30]);
  assign t[351] = (x[33]);
  assign t[352] = (x[33]);
  assign t[353] = (x[36]);
  assign t[354] = (x[36]);
  assign t[355] = (x[39]);
  assign t[356] = (x[39]);
  assign t[357] = (x[44]);
  assign t[358] = (x[44]);
  assign t[359] = (x[49]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[49]);
  assign t[361] = (x[52]);
  assign t[362] = (x[52]);
  assign t[363] = (x[55]);
  assign t[364] = (x[55]);
  assign t[365] = (x[58]);
  assign t[366] = (x[58]);
  assign t[367] = (x[63]);
  assign t[368] = (x[63]);
  assign t[369] = (x[68]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[68]);
  assign t[371] = (x[71]);
  assign t[372] = (x[71]);
  assign t[373] = (x[74]);
  assign t[374] = (x[74]);
  assign t[375] = (x[77]);
  assign t[376] = (x[77]);
  assign t[377] = (x[80]);
  assign t[378] = (x[80]);
  assign t[379] = (x[83]);
  assign t[37] = t[58] ^ t[44];
  assign t[380] = (x[83]);
  assign t[381] = (x[86]);
  assign t[382] = (x[86]);
  assign t[383] = (x[89]);
  assign t[384] = (x[89]);
  assign t[385] = (x[92]);
  assign t[386] = (x[92]);
  assign t[387] = (x[95]);
  assign t[388] = (x[95]);
  assign t[389] = (x[98]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[390] = (x[98]);
  assign t[391] = (x[101]);
  assign t[392] = (x[101]);
  assign t[393] = (x[104]);
  assign t[394] = (x[104]);
  assign t[395] = (x[107]);
  assign t[396] = (x[107]);
  assign t[397] = (x[110]);
  assign t[398] = (x[110]);
  assign t[399] = (x[113]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[113]);
  assign t[401] = (x[116]);
  assign t[402] = (x[116]);
  assign t[403] = (x[119]);
  assign t[404] = (x[119]);
  assign t[405] = (x[122]);
  assign t[406] = (x[122]);
  assign t[407] = (x[125]);
  assign t[408] = (x[125]);
  assign t[409] = (x[128]);
  assign t[40] = t[62] ? x[29] : x[28];
  assign t[410] = (x[128]);
  assign t[411] = (x[131]);
  assign t[412] = (x[131]);
  assign t[413] = (x[134]);
  assign t[414] = (x[134]);
  assign t[415] = (x[137]);
  assign t[416] = (x[137]);
  assign t[417] = (x[140]);
  assign t[418] = (x[140]);
  assign t[419] = (x[143]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[420] = (x[143]);
  assign t[421] = (x[146]);
  assign t[422] = (x[146]);
  assign t[423] = (x[149]);
  assign t[424] = (x[149]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[72] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = t[75] | t[119];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[120];
  assign t[54] = t[49] ? x[43] : x[42];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = t[83] | t[121];
  assign t[58] = t[62] ? x[48] : x[47];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[84] | t[59]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[124];
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = t[90] | t[125];
  assign t[67] = t[62] ? x[62] : x[61];
  assign t[68] = ~(t[91] & t[92]);
  assign t[69] = t[93] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[67] : x[66];
  assign t[71] = ~(t[94] & t[95]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[96] | t[73]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[97] | t[76]);
  assign t[79] = ~(t[98] & t[99]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[100] | t[132];
  assign t[81] = ~(t[133]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[101] | t[81]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[48]);
  assign t[106] = ~(t[129] | t[142]);
  assign t[107] = ~(t[127]);
  assign t[108] = ~(t[226]);
  assign t[109] = ~(t[227]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[143] | t[144]);
  assign t[111] = t[30] ? x[95] : x[94];
  assign t[112] = ~(t[145] & t[146]);
  assign t[113] = ~(t[228]);
  assign t[114] = ~(t[229]);
  assign t[115] = ~(t[147] | t[148]);
  assign t[116] = ~(t[149] | t[150]);
  assign t[117] = ~(t[230] | t[151]);
  assign t[118] = t[30] ? x[106] : x[105];
  assign t[119] = ~(t[83] & t[152]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[204]);
  assign t[121] = ~(t[205] & t[153]);
  assign t[122] = ~(x[4] & t[154]);
  assign t[123] = ~(t[155] & t[205]);
  assign t[124] = ~(t[156] & t[157]);
  assign t[125] = ~(t[120] | t[158]);
  assign t[126] = ~(t[120] | t[159]);
  assign t[127] = ~(t[79] | t[160]);
  assign t[128] = ~(t[161] & t[162]);
  assign t[129] = ~(t[79] | t[163]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[231]);
  assign t[131] = ~(t[218] | t[219]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[233]);
  assign t[134] = ~(t[164] | t[165]);
  assign t[135] = ~(t[138] | t[166]);
  assign t[136] = ~(t[234]);
  assign t[137] = ~(t[221] | t[222]);
  assign t[138] = ~(t[167] & t[168]);
  assign t[139] = ~(t[169] & t[31]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[235]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[170] & t[83]);
  assign t[143] = ~(t[236]);
  assign t[144] = ~(t[226] | t[227]);
  assign t[145] = ~(t[171] | t[126]);
  assign t[146] = ~(t[172] | t[173]);
  assign t[147] = ~(t[237]);
  assign t[148] = ~(t[228] | t[229]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[239]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[176] | t[177]);
  assign t[153] = ~(x[4] | t[178]);
  assign t[154] = ~(t[203] | t[205]);
  assign t[155] = ~(x[4] | t[203]);
  assign t[156] = x[4] & t[203];
  assign t[157] = ~(t[205]);
  assign t[158] = t[202] ? t[124] : t[179];
  assign t[159] = t[202] ? t[180] : t[122];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[202] ? t[179] : t[181];
  assign t[161] = ~(t[182] | t[49]);
  assign t[162] = ~(t[51] & t[183]);
  assign t[163] = t[202] ? t[184] : t[180];
  assign t[164] = ~(t[240]);
  assign t[165] = ~(t[232] | t[233]);
  assign t[166] = ~(t[185] & t[186]);
  assign t[167] = ~(t[82] & t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[127] | t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[182] | t[176]);
  assign t[171] = ~(t[120] | t[191]);
  assign t[172] = ~(t[87]);
  assign t[173] = ~(t[79] | t[192]);
  assign t[174] = ~(t[241]);
  assign t[175] = ~(t[238] | t[239]);
  assign t[176] = ~(t[193] & t[194]);
  assign t[177] = ~(t[162] & t[186]);
  assign t[178] = ~(t[203]);
  assign t[179] = ~(t[155] & t[157]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[153] & t[157]);
  assign t[181] = ~(t[156] & t[205]);
  assign t[182] = ~(t[79] | t[195]);
  assign t[183] = t[155] | t[156];
  assign t[184] = ~(x[4] & t[188]);
  assign t[185] = ~(t[126]);
  assign t[186] = t[120] | t[196];
  assign t[187] = ~(t[121] & t[184]);
  assign t[188] = ~(t[203] | t[157]);
  assign t[189] = t[79] & t[202];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[197]);
  assign t[191] = t[202] ? t[179] : t[124];
  assign t[192] = t[202] ? t[121] : t[122];
  assign t[193] = ~(t[171] | t[198]);
  assign t[194] = ~(t[120] & t[199]);
  assign t[195] = t[202] ? t[181] : t[179];
  assign t[196] = t[202] ? t[122] : t[180];
  assign t[197] = t[202] ? t[123] : t[124];
  assign t[198] = ~(t[79] | t[200]);
  assign t[199] = ~(t[122] & t[121]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[180] : t[184];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[10];
  assign t[244] = t[285] ^ x[13];
  assign t[245] = t[286] ^ x[16];
  assign t[246] = t[287] ^ x[19];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[36];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[68];
  assign t[262] = t[303] ^ x[73];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[81];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[98];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[10];
  assign t[327] = t[409] ^ x[9];
  assign t[328] = t[410] ^ x[13];
  assign t[329] = t[411] ^ x[12];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[16];
  assign t[331] = t[413] ^ x[15];
  assign t[332] = t[414] ^ x[19];
  assign t[333] = t[415] ^ x[18];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[36];
  assign t[343] = t[425] ^ x[35];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[68];
  assign t[363] = t[445] ^ x[67];
  assign t[364] = t[446] ^ x[73];
  assign t[365] = t[447] ^ x[72];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[81];
  assign t[369] = t[451] ^ x[80];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[98];
  assign t[379] = t[461] ^ x[97];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[38] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[8]);
  assign t[409] = (x[8]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[11]);
  assign t[411] = (x[11]);
  assign t[412] = (x[14]);
  assign t[413] = (x[14]);
  assign t[414] = (x[17]);
  assign t[415] = (x[17]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[207] | t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[34]);
  assign t[425] = (x[34]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[66]);
  assign t[445] = (x[66]);
  assign t[446] = (x[71]);
  assign t[447] = (x[71]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[79]);
  assign t[451] = (x[79]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[44] ^ t[74]);
  assign t[460] = (x[96]);
  assign t[461] = (x[96]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[204]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = t[205] & t[82];
  assign t[52] = ~(t[83]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[204] ? x[33] : x[32];
  assign t[57] = ~(t[86] & t[87]);
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[210] | t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91] | t[92]);
  assign t[61] = ~(t[93] ^ t[94]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[63] = ~(t[211] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[214] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[105] ? x[50] : x[49];
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[108] | t[109]);
  assign t[73] = ~(t[215] | t[110]);
  assign t[74] = ~(t[111] ^ t[112]);
  assign t[75] = ~(t[113] | t[114]);
  assign t[76] = ~(t[216] | t[115]);
  assign t[77] = ~(t[116] | t[117]);
  assign t[78] = ~(t[118] ^ t[119]);
  assign t[79] = ~(t[120]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[202] ? t[122] : t[121];
  assign t[81] = t[202] ? t[124] : t[123];
  assign t[82] = ~(t[120] | t[202]);
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = ~(t[217]);
  assign t[85] = ~(t[208] | t[209]);
  assign t[86] = ~(t[127] | t[128]);
  assign t[87] = ~(t[129] | t[50]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[220] | t[134]);
  assign t[93] = t[105] ? x[70] : x[69];
  assign t[94] = ~(t[135] & t[107]);
  assign t[95] = ~(t[221]);
  assign t[96] = ~(t[222]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[204] ? x[78] : x[77];
  assign t[99] = t[138] | t[139];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [139:0] x;
 output y;

 wire [487:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[48]);
  assign t[106] = ~(t[129] | t[142]);
  assign t[107] = ~(t[127]);
  assign t[108] = ~(t[226]);
  assign t[109] = ~(t[227]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[143] | t[144]);
  assign t[111] = t[30] ? x[95] : x[94];
  assign t[112] = ~(t[145] & t[146]);
  assign t[113] = ~(t[228]);
  assign t[114] = ~(t[229]);
  assign t[115] = ~(t[147] | t[148]);
  assign t[116] = ~(t[149] | t[150]);
  assign t[117] = ~(t[230] | t[151]);
  assign t[118] = t[30] ? x[106] : x[105];
  assign t[119] = ~(t[83] & t[152]);
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[204]);
  assign t[121] = ~(t[205] & t[153]);
  assign t[122] = ~(x[4] & t[154]);
  assign t[123] = ~(t[155] & t[205]);
  assign t[124] = ~(t[156] & t[157]);
  assign t[125] = ~(t[120] | t[158]);
  assign t[126] = ~(t[120] | t[159]);
  assign t[127] = ~(t[79] | t[160]);
  assign t[128] = ~(t[161] & t[162]);
  assign t[129] = ~(t[79] | t[163]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[231]);
  assign t[131] = ~(t[218] | t[219]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[233]);
  assign t[134] = ~(t[164] | t[165]);
  assign t[135] = ~(t[138] | t[166]);
  assign t[136] = ~(t[234]);
  assign t[137] = ~(t[221] | t[222]);
  assign t[138] = ~(t[167] & t[168]);
  assign t[139] = ~(t[169] & t[31]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[235]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[170] & t[83]);
  assign t[143] = ~(t[236]);
  assign t[144] = ~(t[226] | t[227]);
  assign t[145] = ~(t[171] | t[126]);
  assign t[146] = ~(t[172] | t[173]);
  assign t[147] = ~(t[237]);
  assign t[148] = ~(t[228] | t[229]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[239]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[176] | t[177]);
  assign t[153] = ~(x[4] | t[178]);
  assign t[154] = ~(t[203] | t[205]);
  assign t[155] = ~(x[4] | t[203]);
  assign t[156] = x[4] & t[203];
  assign t[157] = ~(t[205]);
  assign t[158] = t[202] ? t[124] : t[179];
  assign t[159] = t[202] ? t[180] : t[122];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[202] ? t[179] : t[181];
  assign t[161] = ~(t[182] | t[49]);
  assign t[162] = ~(t[51] & t[183]);
  assign t[163] = t[202] ? t[184] : t[180];
  assign t[164] = ~(t[240]);
  assign t[165] = ~(t[232] | t[233]);
  assign t[166] = ~(t[185] & t[186]);
  assign t[167] = ~(t[82] & t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[127] | t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[182] | t[176]);
  assign t[171] = ~(t[120] | t[191]);
  assign t[172] = ~(t[87]);
  assign t[173] = ~(t[79] | t[192]);
  assign t[174] = ~(t[241]);
  assign t[175] = ~(t[238] | t[239]);
  assign t[176] = ~(t[193] & t[194]);
  assign t[177] = ~(t[162] & t[186]);
  assign t[178] = ~(t[203]);
  assign t[179] = ~(t[155] & t[157]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[153] & t[157]);
  assign t[181] = ~(t[156] & t[205]);
  assign t[182] = ~(t[79] | t[195]);
  assign t[183] = t[155] | t[156];
  assign t[184] = ~(x[4] & t[188]);
  assign t[185] = ~(t[126]);
  assign t[186] = t[120] | t[196];
  assign t[187] = ~(t[121] & t[184]);
  assign t[188] = ~(t[203] | t[157]);
  assign t[189] = t[79] & t[202];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[197]);
  assign t[191] = t[202] ? t[179] : t[124];
  assign t[192] = t[202] ? t[121] : t[122];
  assign t[193] = ~(t[171] | t[198]);
  assign t[194] = ~(t[120] & t[199]);
  assign t[195] = t[202] ? t[181] : t[179];
  assign t[196] = t[202] ? t[122] : t[180];
  assign t[197] = t[202] ? t[123] : t[124];
  assign t[198] = ~(t[79] | t[200]);
  assign t[199] = ~(t[122] & t[121]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[180] : t[184];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[2];
  assign t[243] = t[284] ^ x[10];
  assign t[244] = t[285] ^ x[13];
  assign t[245] = t[286] ^ x[16];
  assign t[246] = t[287] ^ x[19];
  assign t[247] = t[288] ^ x[22];
  assign t[248] = t[289] ^ x[25];
  assign t[249] = t[290] ^ x[28];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[31];
  assign t[251] = t[292] ^ x[36];
  assign t[252] = t[293] ^ x[39];
  assign t[253] = t[294] ^ x[42];
  assign t[254] = t[295] ^ x[45];
  assign t[255] = t[296] ^ x[48];
  assign t[256] = t[297] ^ x[53];
  assign t[257] = t[298] ^ x[56];
  assign t[258] = t[299] ^ x[59];
  assign t[259] = t[300] ^ x[62];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[65];
  assign t[261] = t[302] ^ x[68];
  assign t[262] = t[303] ^ x[73];
  assign t[263] = t[304] ^ x[76];
  assign t[264] = t[305] ^ x[81];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[87];
  assign t[267] = t[308] ^ x[90];
  assign t[268] = t[309] ^ x[93];
  assign t[269] = t[310] ^ x[98];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[104];
  assign t[272] = t[313] ^ x[109];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[115];
  assign t[275] = t[316] ^ x[118];
  assign t[276] = t[317] ^ x[121];
  assign t[277] = t[318] ^ x[124];
  assign t[278] = t[319] ^ x[127];
  assign t[279] = t[320] ^ x[130];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[133];
  assign t[281] = t[322] ^ x[136];
  assign t[282] = t[323] ^ x[139];
  assign t[283] = (t[324] & ~t[325]);
  assign t[284] = (t[326] & ~t[327]);
  assign t[285] = (t[328] & ~t[329]);
  assign t[286] = (t[330] & ~t[331]);
  assign t[287] = (t[332] & ~t[333]);
  assign t[288] = (t[334] & ~t[335]);
  assign t[289] = (t[336] & ~t[337]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[338] & ~t[339]);
  assign t[291] = (t[340] & ~t[341]);
  assign t[292] = (t[342] & ~t[343]);
  assign t[293] = (t[344] & ~t[345]);
  assign t[294] = (t[346] & ~t[347]);
  assign t[295] = (t[348] & ~t[349]);
  assign t[296] = (t[350] & ~t[351]);
  assign t[297] = (t[352] & ~t[353]);
  assign t[298] = (t[354] & ~t[355]);
  assign t[299] = (t[356] & ~t[357]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[358] & ~t[359]);
  assign t[301] = (t[360] & ~t[361]);
  assign t[302] = (t[362] & ~t[363]);
  assign t[303] = (t[364] & ~t[365]);
  assign t[304] = (t[366] & ~t[367]);
  assign t[305] = (t[368] & ~t[369]);
  assign t[306] = (t[370] & ~t[371]);
  assign t[307] = (t[372] & ~t[373]);
  assign t[308] = (t[374] & ~t[375]);
  assign t[309] = (t[376] & ~t[377]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[378] & ~t[379]);
  assign t[311] = (t[380] & ~t[381]);
  assign t[312] = (t[382] & ~t[383]);
  assign t[313] = (t[384] & ~t[385]);
  assign t[314] = (t[386] & ~t[387]);
  assign t[315] = (t[388] & ~t[389]);
  assign t[316] = (t[390] & ~t[391]);
  assign t[317] = (t[392] & ~t[393]);
  assign t[318] = (t[394] & ~t[395]);
  assign t[319] = (t[396] & ~t[397]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[398] & ~t[399]);
  assign t[321] = (t[400] & ~t[401]);
  assign t[322] = (t[402] & ~t[403]);
  assign t[323] = (t[404] & ~t[405]);
  assign t[324] = t[406] ^ x[2];
  assign t[325] = t[407] ^ x[1];
  assign t[326] = t[408] ^ x[10];
  assign t[327] = t[409] ^ x[9];
  assign t[328] = t[410] ^ x[13];
  assign t[329] = t[411] ^ x[12];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[16];
  assign t[331] = t[413] ^ x[15];
  assign t[332] = t[414] ^ x[19];
  assign t[333] = t[415] ^ x[18];
  assign t[334] = t[416] ^ x[22];
  assign t[335] = t[417] ^ x[21];
  assign t[336] = t[418] ^ x[25];
  assign t[337] = t[419] ^ x[24];
  assign t[338] = t[420] ^ x[28];
  assign t[339] = t[421] ^ x[27];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[31];
  assign t[341] = t[423] ^ x[30];
  assign t[342] = t[424] ^ x[36];
  assign t[343] = t[425] ^ x[35];
  assign t[344] = t[426] ^ x[39];
  assign t[345] = t[427] ^ x[38];
  assign t[346] = t[428] ^ x[42];
  assign t[347] = t[429] ^ x[41];
  assign t[348] = t[430] ^ x[45];
  assign t[349] = t[431] ^ x[44];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[432] ^ x[48];
  assign t[351] = t[433] ^ x[47];
  assign t[352] = t[434] ^ x[53];
  assign t[353] = t[435] ^ x[52];
  assign t[354] = t[436] ^ x[56];
  assign t[355] = t[437] ^ x[55];
  assign t[356] = t[438] ^ x[59];
  assign t[357] = t[439] ^ x[58];
  assign t[358] = t[440] ^ x[62];
  assign t[359] = t[441] ^ x[61];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[442] ^ x[65];
  assign t[361] = t[443] ^ x[64];
  assign t[362] = t[444] ^ x[68];
  assign t[363] = t[445] ^ x[67];
  assign t[364] = t[446] ^ x[73];
  assign t[365] = t[447] ^ x[72];
  assign t[366] = t[448] ^ x[76];
  assign t[367] = t[449] ^ x[75];
  assign t[368] = t[450] ^ x[81];
  assign t[369] = t[451] ^ x[80];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[452] ^ x[84];
  assign t[371] = t[453] ^ x[83];
  assign t[372] = t[454] ^ x[87];
  assign t[373] = t[455] ^ x[86];
  assign t[374] = t[456] ^ x[90];
  assign t[375] = t[457] ^ x[89];
  assign t[376] = t[458] ^ x[93];
  assign t[377] = t[459] ^ x[92];
  assign t[378] = t[460] ^ x[98];
  assign t[379] = t[461] ^ x[97];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[462] ^ x[101];
  assign t[381] = t[463] ^ x[100];
  assign t[382] = t[464] ^ x[104];
  assign t[383] = t[465] ^ x[103];
  assign t[384] = t[466] ^ x[109];
  assign t[385] = t[467] ^ x[108];
  assign t[386] = t[468] ^ x[112];
  assign t[387] = t[469] ^ x[111];
  assign t[388] = t[470] ^ x[115];
  assign t[389] = t[471] ^ x[114];
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = t[472] ^ x[118];
  assign t[391] = t[473] ^ x[117];
  assign t[392] = t[474] ^ x[121];
  assign t[393] = t[475] ^ x[120];
  assign t[394] = t[476] ^ x[124];
  assign t[395] = t[477] ^ x[123];
  assign t[396] = t[478] ^ x[127];
  assign t[397] = t[479] ^ x[126];
  assign t[398] = t[480] ^ x[130];
  assign t[399] = t[481] ^ x[129];
  assign t[39] = ~(t[38] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[133];
  assign t[401] = t[483] ^ x[132];
  assign t[402] = t[484] ^ x[136];
  assign t[403] = t[485] ^ x[135];
  assign t[404] = t[486] ^ x[139];
  assign t[405] = t[487] ^ x[138];
  assign t[406] = (x[0]);
  assign t[407] = (x[0]);
  assign t[408] = (x[8]);
  assign t[409] = (x[8]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[11]);
  assign t[411] = (x[11]);
  assign t[412] = (x[14]);
  assign t[413] = (x[14]);
  assign t[414] = (x[17]);
  assign t[415] = (x[17]);
  assign t[416] = (x[20]);
  assign t[417] = (x[20]);
  assign t[418] = (x[23]);
  assign t[419] = (x[23]);
  assign t[41] = ~(t[207] | t[67]);
  assign t[420] = (x[26]);
  assign t[421] = (x[26]);
  assign t[422] = (x[29]);
  assign t[423] = (x[29]);
  assign t[424] = (x[34]);
  assign t[425] = (x[34]);
  assign t[426] = (x[37]);
  assign t[427] = (x[37]);
  assign t[428] = (x[40]);
  assign t[429] = (x[40]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[43]);
  assign t[431] = (x[43]);
  assign t[432] = (x[46]);
  assign t[433] = (x[46]);
  assign t[434] = (x[51]);
  assign t[435] = (x[51]);
  assign t[436] = (x[54]);
  assign t[437] = (x[54]);
  assign t[438] = (x[57]);
  assign t[439] = (x[57]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = (x[60]);
  assign t[441] = (x[60]);
  assign t[442] = (x[63]);
  assign t[443] = (x[63]);
  assign t[444] = (x[66]);
  assign t[445] = (x[66]);
  assign t[446] = (x[71]);
  assign t[447] = (x[71]);
  assign t[448] = (x[74]);
  assign t[449] = (x[74]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = (x[79]);
  assign t[451] = (x[79]);
  assign t[452] = (x[82]);
  assign t[453] = (x[82]);
  assign t[454] = (x[85]);
  assign t[455] = (x[85]);
  assign t[456] = (x[88]);
  assign t[457] = (x[88]);
  assign t[458] = (x[91]);
  assign t[459] = (x[91]);
  assign t[45] = ~(t[44] ^ t[74]);
  assign t[460] = (x[96]);
  assign t[461] = (x[96]);
  assign t[462] = (x[99]);
  assign t[463] = (x[99]);
  assign t[464] = (x[102]);
  assign t[465] = (x[102]);
  assign t[466] = (x[107]);
  assign t[467] = (x[107]);
  assign t[468] = (x[110]);
  assign t[469] = (x[110]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[113]);
  assign t[471] = (x[113]);
  assign t[472] = (x[116]);
  assign t[473] = (x[116]);
  assign t[474] = (x[119]);
  assign t[475] = (x[119]);
  assign t[476] = (x[122]);
  assign t[477] = (x[122]);
  assign t[478] = (x[125]);
  assign t[479] = (x[125]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[128]);
  assign t[481] = (x[128]);
  assign t[482] = (x[131]);
  assign t[483] = (x[131]);
  assign t[484] = (x[134]);
  assign t[485] = (x[134]);
  assign t[486] = (x[137]);
  assign t[487] = (x[137]);
  assign t[48] = ~(t[204]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = t[205] & t[82];
  assign t[52] = ~(t[83]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[204] ? x[33] : x[32];
  assign t[57] = ~(t[86] & t[87]);
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[210] | t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91] | t[92]);
  assign t[61] = ~(t[93] ^ t[94]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[63] = ~(t[211] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[214] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[105] ? x[50] : x[49];
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[108] | t[109]);
  assign t[73] = ~(t[215] | t[110]);
  assign t[74] = ~(t[111] ^ t[112]);
  assign t[75] = ~(t[113] | t[114]);
  assign t[76] = ~(t[216] | t[115]);
  assign t[77] = ~(t[116] | t[117]);
  assign t[78] = ~(t[118] ^ t[119]);
  assign t[79] = ~(t[120]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[202] ? t[122] : t[121];
  assign t[81] = t[202] ? t[124] : t[123];
  assign t[82] = ~(t[120] | t[202]);
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = ~(t[217]);
  assign t[85] = ~(t[208] | t[209]);
  assign t[86] = ~(t[127] | t[128]);
  assign t[87] = ~(t[129] | t[50]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[220] | t[134]);
  assign t[93] = t[105] ? x[70] : x[69];
  assign t[94] = ~(t[135] & t[107]);
  assign t[95] = ~(t[221]);
  assign t[96] = ~(t[222]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[204] ? x[78] : x[77];
  assign t[99] = t[138] | t[139];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind246(x, y);
 input [112:0] x;
 output y;

 wire [316:0] t;
  assign t[0] = t[1] ? t[2] : t[93];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = t[157] ^ x[2];
  assign t[126] = t[158] ^ x[10];
  assign t[127] = t[159] ^ x[13];
  assign t[128] = t[160] ^ x[16];
  assign t[129] = t[161] ^ x[19];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[25];
  assign t[132] = t[164] ^ x[30];
  assign t[133] = t[165] ^ x[33];
  assign t[134] = t[166] ^ x[38];
  assign t[135] = t[167] ^ x[41];
  assign t[136] = t[168] ^ x[44];
  assign t[137] = t[169] ^ x[49];
  assign t[138] = t[170] ^ x[52];
  assign t[139] = t[171] ^ x[57];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[60];
  assign t[141] = t[173] ^ x[63];
  assign t[142] = t[174] ^ x[66];
  assign t[143] = t[175] ^ x[69];
  assign t[144] = t[176] ^ x[74];
  assign t[145] = t[177] ^ x[77];
  assign t[146] = t[178] ^ x[82];
  assign t[147] = t[179] ^ x[85];
  assign t[148] = t[180] ^ x[88];
  assign t[149] = t[181] ^ x[91];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[94];
  assign t[151] = t[183] ^ x[97];
  assign t[152] = t[184] ^ x[100];
  assign t[153] = t[185] ^ x[103];
  assign t[154] = t[186] ^ x[106];
  assign t[155] = t[187] ^ x[109];
  assign t[156] = t[188] ^ x[112];
  assign t[157] = (t[189] & ~t[190]);
  assign t[158] = (t[191] & ~t[192]);
  assign t[159] = (t[193] & ~t[194]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[195] & ~t[196]);
  assign t[161] = (t[197] & ~t[198]);
  assign t[162] = (t[199] & ~t[200]);
  assign t[163] = (t[201] & ~t[202]);
  assign t[164] = (t[203] & ~t[204]);
  assign t[165] = (t[205] & ~t[206]);
  assign t[166] = (t[207] & ~t[208]);
  assign t[167] = (t[209] & ~t[210]);
  assign t[168] = (t[211] & ~t[212]);
  assign t[169] = (t[213] & ~t[214]);
  assign t[16] = ~(t[94] & t[95]);
  assign t[170] = (t[215] & ~t[216]);
  assign t[171] = (t[217] & ~t[218]);
  assign t[172] = (t[219] & ~t[220]);
  assign t[173] = (t[221] & ~t[222]);
  assign t[174] = (t[223] & ~t[224]);
  assign t[175] = (t[225] & ~t[226]);
  assign t[176] = (t[227] & ~t[228]);
  assign t[177] = (t[229] & ~t[230]);
  assign t[178] = (t[231] & ~t[232]);
  assign t[179] = (t[233] & ~t[234]);
  assign t[17] = ~(t[96] & t[97]);
  assign t[180] = (t[235] & ~t[236]);
  assign t[181] = (t[237] & ~t[238]);
  assign t[182] = (t[239] & ~t[240]);
  assign t[183] = (t[241] & ~t[242]);
  assign t[184] = (t[243] & ~t[244]);
  assign t[185] = (t[245] & ~t[246]);
  assign t[186] = (t[247] & ~t[248]);
  assign t[187] = (t[249] & ~t[250]);
  assign t[188] = (t[251] & ~t[252]);
  assign t[189] = t[253] ^ x[2];
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[1];
  assign t[191] = t[255] ^ x[10];
  assign t[192] = t[256] ^ x[9];
  assign t[193] = t[257] ^ x[13];
  assign t[194] = t[258] ^ x[12];
  assign t[195] = t[259] ^ x[16];
  assign t[196] = t[260] ^ x[15];
  assign t[197] = t[261] ^ x[19];
  assign t[198] = t[262] ^ x[18];
  assign t[199] = t[263] ^ x[22];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[21];
  assign t[201] = t[265] ^ x[25];
  assign t[202] = t[266] ^ x[24];
  assign t[203] = t[267] ^ x[30];
  assign t[204] = t[268] ^ x[29];
  assign t[205] = t[269] ^ x[33];
  assign t[206] = t[270] ^ x[32];
  assign t[207] = t[271] ^ x[38];
  assign t[208] = t[272] ^ x[37];
  assign t[209] = t[273] ^ x[41];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[40];
  assign t[211] = t[275] ^ x[44];
  assign t[212] = t[276] ^ x[43];
  assign t[213] = t[277] ^ x[49];
  assign t[214] = t[278] ^ x[48];
  assign t[215] = t[279] ^ x[52];
  assign t[216] = t[280] ^ x[51];
  assign t[217] = t[281] ^ x[57];
  assign t[218] = t[282] ^ x[56];
  assign t[219] = t[283] ^ x[60];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[59];
  assign t[221] = t[285] ^ x[63];
  assign t[222] = t[286] ^ x[62];
  assign t[223] = t[287] ^ x[66];
  assign t[224] = t[288] ^ x[65];
  assign t[225] = t[289] ^ x[69];
  assign t[226] = t[290] ^ x[68];
  assign t[227] = t[291] ^ x[74];
  assign t[228] = t[292] ^ x[73];
  assign t[229] = t[293] ^ x[77];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[294] ^ x[76];
  assign t[231] = t[295] ^ x[82];
  assign t[232] = t[296] ^ x[81];
  assign t[233] = t[297] ^ x[85];
  assign t[234] = t[298] ^ x[84];
  assign t[235] = t[299] ^ x[88];
  assign t[236] = t[300] ^ x[87];
  assign t[237] = t[301] ^ x[91];
  assign t[238] = t[302] ^ x[90];
  assign t[239] = t[303] ^ x[94];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[93];
  assign t[241] = t[305] ^ x[97];
  assign t[242] = t[306] ^ x[96];
  assign t[243] = t[307] ^ x[100];
  assign t[244] = t[308] ^ x[99];
  assign t[245] = t[309] ^ x[103];
  assign t[246] = t[310] ^ x[102];
  assign t[247] = t[311] ^ x[106];
  assign t[248] = t[312] ^ x[105];
  assign t[249] = t[313] ^ x[109];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[108];
  assign t[251] = t[315] ^ x[112];
  assign t[252] = t[316] ^ x[111];
  assign t[253] = (x[0]);
  assign t[254] = (x[0]);
  assign t[255] = (x[8]);
  assign t[256] = (x[8]);
  assign t[257] = (x[11]);
  assign t[258] = (x[11]);
  assign t[259] = (x[14]);
  assign t[25] = ~(t[96]);
  assign t[260] = (x[14]);
  assign t[261] = (x[17]);
  assign t[262] = (x[17]);
  assign t[263] = (x[20]);
  assign t[264] = (x[20]);
  assign t[265] = (x[23]);
  assign t[266] = (x[23]);
  assign t[267] = (x[28]);
  assign t[268] = (x[28]);
  assign t[269] = (x[31]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[36]);
  assign t[272] = (x[36]);
  assign t[273] = (x[39]);
  assign t[274] = (x[39]);
  assign t[275] = (x[42]);
  assign t[276] = (x[42]);
  assign t[277] = (x[47]);
  assign t[278] = (x[47]);
  assign t[279] = (x[50]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[55]);
  assign t[282] = (x[55]);
  assign t[283] = (x[58]);
  assign t[284] = (x[58]);
  assign t[285] = (x[61]);
  assign t[286] = (x[61]);
  assign t[287] = (x[64]);
  assign t[288] = (x[64]);
  assign t[289] = (x[67]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[72]);
  assign t[292] = (x[72]);
  assign t[293] = (x[75]);
  assign t[294] = (x[75]);
  assign t[295] = (x[80]);
  assign t[296] = (x[80]);
  assign t[297] = (x[83]);
  assign t[298] = (x[83]);
  assign t[299] = (x[86]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[89]);
  assign t[302] = (x[89]);
  assign t[303] = (x[92]);
  assign t[304] = (x[92]);
  assign t[305] = (x[95]);
  assign t[306] = (x[95]);
  assign t[307] = (x[98]);
  assign t[308] = (x[98]);
  assign t[309] = (x[101]);
  assign t[30] = ~(t[98] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[104]);
  assign t[312] = (x[104]);
  assign t[313] = (x[107]);
  assign t[314] = (x[107]);
  assign t[315] = (x[110]);
  assign t[316] = (x[110]);
  assign t[31] = ~(t[99] & t[46]);
  assign t[32] = t[96] ? x[27] : x[26];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[33];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = t[52] ^ t[53];
  assign t[37] = ~(t[100] & t[54]);
  assign t[38] = ~(t[101] & t[55]);
  assign t[39] = t[56] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[62];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[43];
  assign t[45] = ~(t[102]);
  assign t[46] = ~(t[102] & t[66]);
  assign t[47] = ~(t[103] & t[67]);
  assign t[48] = ~(t[104] & t[68]);
  assign t[49] = t[96] ? x[46] : x[45];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[96] ? x[54] : x[53];
  assign t[53] = ~(t[71] & t[72]);
  assign t[54] = ~(t[107]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[25]);
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[111] & t[77]);
  assign t[61] = t[18] ? x[71] : x[70];
  assign t[62] = ~(t[78] & t[79]);
  assign t[63] = ~(t[112] & t[80]);
  assign t[64] = ~(t[113] & t[81]);
  assign t[65] = t[18] ? x[79] : x[78];
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[114]);
  assign t[68] = ~(t[114] & t[82]);
  assign t[69] = ~(t[115]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[118]);
  assign t[75] = ~(t[118] & t[86]);
  assign t[76] = ~(t[119]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[123]);
  assign t[85] = ~(t[123] & t[91]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[124]);
  assign t[89] = ~(t[124] & t[92]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[120]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [112:0] x;
 output y;

 wire [316:0] t;
  assign t[0] = t[1] ? t[2] : t[93];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = t[157] ^ x[2];
  assign t[126] = t[158] ^ x[10];
  assign t[127] = t[159] ^ x[13];
  assign t[128] = t[160] ^ x[16];
  assign t[129] = t[161] ^ x[19];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[25];
  assign t[132] = t[164] ^ x[30];
  assign t[133] = t[165] ^ x[33];
  assign t[134] = t[166] ^ x[38];
  assign t[135] = t[167] ^ x[41];
  assign t[136] = t[168] ^ x[44];
  assign t[137] = t[169] ^ x[49];
  assign t[138] = t[170] ^ x[52];
  assign t[139] = t[171] ^ x[57];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[60];
  assign t[141] = t[173] ^ x[63];
  assign t[142] = t[174] ^ x[66];
  assign t[143] = t[175] ^ x[69];
  assign t[144] = t[176] ^ x[74];
  assign t[145] = t[177] ^ x[77];
  assign t[146] = t[178] ^ x[82];
  assign t[147] = t[179] ^ x[85];
  assign t[148] = t[180] ^ x[88];
  assign t[149] = t[181] ^ x[91];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[94];
  assign t[151] = t[183] ^ x[97];
  assign t[152] = t[184] ^ x[100];
  assign t[153] = t[185] ^ x[103];
  assign t[154] = t[186] ^ x[106];
  assign t[155] = t[187] ^ x[109];
  assign t[156] = t[188] ^ x[112];
  assign t[157] = (t[189] & ~t[190]);
  assign t[158] = (t[191] & ~t[192]);
  assign t[159] = (t[193] & ~t[194]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[195] & ~t[196]);
  assign t[161] = (t[197] & ~t[198]);
  assign t[162] = (t[199] & ~t[200]);
  assign t[163] = (t[201] & ~t[202]);
  assign t[164] = (t[203] & ~t[204]);
  assign t[165] = (t[205] & ~t[206]);
  assign t[166] = (t[207] & ~t[208]);
  assign t[167] = (t[209] & ~t[210]);
  assign t[168] = (t[211] & ~t[212]);
  assign t[169] = (t[213] & ~t[214]);
  assign t[16] = ~(t[94] & t[95]);
  assign t[170] = (t[215] & ~t[216]);
  assign t[171] = (t[217] & ~t[218]);
  assign t[172] = (t[219] & ~t[220]);
  assign t[173] = (t[221] & ~t[222]);
  assign t[174] = (t[223] & ~t[224]);
  assign t[175] = (t[225] & ~t[226]);
  assign t[176] = (t[227] & ~t[228]);
  assign t[177] = (t[229] & ~t[230]);
  assign t[178] = (t[231] & ~t[232]);
  assign t[179] = (t[233] & ~t[234]);
  assign t[17] = ~(t[96] & t[97]);
  assign t[180] = (t[235] & ~t[236]);
  assign t[181] = (t[237] & ~t[238]);
  assign t[182] = (t[239] & ~t[240]);
  assign t[183] = (t[241] & ~t[242]);
  assign t[184] = (t[243] & ~t[244]);
  assign t[185] = (t[245] & ~t[246]);
  assign t[186] = (t[247] & ~t[248]);
  assign t[187] = (t[249] & ~t[250]);
  assign t[188] = (t[251] & ~t[252]);
  assign t[189] = t[253] ^ x[2];
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[1];
  assign t[191] = t[255] ^ x[10];
  assign t[192] = t[256] ^ x[9];
  assign t[193] = t[257] ^ x[13];
  assign t[194] = t[258] ^ x[12];
  assign t[195] = t[259] ^ x[16];
  assign t[196] = t[260] ^ x[15];
  assign t[197] = t[261] ^ x[19];
  assign t[198] = t[262] ^ x[18];
  assign t[199] = t[263] ^ x[22];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[21];
  assign t[201] = t[265] ^ x[25];
  assign t[202] = t[266] ^ x[24];
  assign t[203] = t[267] ^ x[30];
  assign t[204] = t[268] ^ x[29];
  assign t[205] = t[269] ^ x[33];
  assign t[206] = t[270] ^ x[32];
  assign t[207] = t[271] ^ x[38];
  assign t[208] = t[272] ^ x[37];
  assign t[209] = t[273] ^ x[41];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[40];
  assign t[211] = t[275] ^ x[44];
  assign t[212] = t[276] ^ x[43];
  assign t[213] = t[277] ^ x[49];
  assign t[214] = t[278] ^ x[48];
  assign t[215] = t[279] ^ x[52];
  assign t[216] = t[280] ^ x[51];
  assign t[217] = t[281] ^ x[57];
  assign t[218] = t[282] ^ x[56];
  assign t[219] = t[283] ^ x[60];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[59];
  assign t[221] = t[285] ^ x[63];
  assign t[222] = t[286] ^ x[62];
  assign t[223] = t[287] ^ x[66];
  assign t[224] = t[288] ^ x[65];
  assign t[225] = t[289] ^ x[69];
  assign t[226] = t[290] ^ x[68];
  assign t[227] = t[291] ^ x[74];
  assign t[228] = t[292] ^ x[73];
  assign t[229] = t[293] ^ x[77];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[294] ^ x[76];
  assign t[231] = t[295] ^ x[82];
  assign t[232] = t[296] ^ x[81];
  assign t[233] = t[297] ^ x[85];
  assign t[234] = t[298] ^ x[84];
  assign t[235] = t[299] ^ x[88];
  assign t[236] = t[300] ^ x[87];
  assign t[237] = t[301] ^ x[91];
  assign t[238] = t[302] ^ x[90];
  assign t[239] = t[303] ^ x[94];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[304] ^ x[93];
  assign t[241] = t[305] ^ x[97];
  assign t[242] = t[306] ^ x[96];
  assign t[243] = t[307] ^ x[100];
  assign t[244] = t[308] ^ x[99];
  assign t[245] = t[309] ^ x[103];
  assign t[246] = t[310] ^ x[102];
  assign t[247] = t[311] ^ x[106];
  assign t[248] = t[312] ^ x[105];
  assign t[249] = t[313] ^ x[109];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[314] ^ x[108];
  assign t[251] = t[315] ^ x[112];
  assign t[252] = t[316] ^ x[111];
  assign t[253] = (x[0]);
  assign t[254] = (x[0]);
  assign t[255] = (x[8]);
  assign t[256] = (x[8]);
  assign t[257] = (x[11]);
  assign t[258] = (x[11]);
  assign t[259] = (x[14]);
  assign t[25] = ~(t[96]);
  assign t[260] = (x[14]);
  assign t[261] = (x[17]);
  assign t[262] = (x[17]);
  assign t[263] = (x[20]);
  assign t[264] = (x[20]);
  assign t[265] = (x[23]);
  assign t[266] = (x[23]);
  assign t[267] = (x[28]);
  assign t[268] = (x[28]);
  assign t[269] = (x[31]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[31]);
  assign t[271] = (x[36]);
  assign t[272] = (x[36]);
  assign t[273] = (x[39]);
  assign t[274] = (x[39]);
  assign t[275] = (x[42]);
  assign t[276] = (x[42]);
  assign t[277] = (x[47]);
  assign t[278] = (x[47]);
  assign t[279] = (x[50]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[50]);
  assign t[281] = (x[55]);
  assign t[282] = (x[55]);
  assign t[283] = (x[58]);
  assign t[284] = (x[58]);
  assign t[285] = (x[61]);
  assign t[286] = (x[61]);
  assign t[287] = (x[64]);
  assign t[288] = (x[64]);
  assign t[289] = (x[67]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[72]);
  assign t[292] = (x[72]);
  assign t[293] = (x[75]);
  assign t[294] = (x[75]);
  assign t[295] = (x[80]);
  assign t[296] = (x[80]);
  assign t[297] = (x[83]);
  assign t[298] = (x[83]);
  assign t[299] = (x[86]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[89]);
  assign t[302] = (x[89]);
  assign t[303] = (x[92]);
  assign t[304] = (x[92]);
  assign t[305] = (x[95]);
  assign t[306] = (x[95]);
  assign t[307] = (x[98]);
  assign t[308] = (x[98]);
  assign t[309] = (x[101]);
  assign t[30] = ~(t[98] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[104]);
  assign t[312] = (x[104]);
  assign t[313] = (x[107]);
  assign t[314] = (x[107]);
  assign t[315] = (x[110]);
  assign t[316] = (x[110]);
  assign t[31] = ~(t[99] & t[46]);
  assign t[32] = t[96] ? x[27] : x[26];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[33];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = t[52] ^ t[53];
  assign t[37] = ~(t[100] & t[54]);
  assign t[38] = ~(t[101] & t[55]);
  assign t[39] = t[56] ? x[35] : x[34];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[62];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[43];
  assign t[45] = ~(t[102]);
  assign t[46] = ~(t[102] & t[66]);
  assign t[47] = ~(t[103] & t[67]);
  assign t[48] = ~(t[104] & t[68]);
  assign t[49] = t[96] ? x[46] : x[45];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[96] ? x[54] : x[53];
  assign t[53] = ~(t[71] & t[72]);
  assign t[54] = ~(t[107]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[25]);
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[111] & t[77]);
  assign t[61] = t[18] ? x[71] : x[70];
  assign t[62] = ~(t[78] & t[79]);
  assign t[63] = ~(t[112] & t[80]);
  assign t[64] = ~(t[113] & t[81]);
  assign t[65] = t[18] ? x[79] : x[78];
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[114]);
  assign t[68] = ~(t[114] & t[82]);
  assign t[69] = ~(t[115]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[118]);
  assign t[75] = ~(t[118] & t[86]);
  assign t[76] = ~(t[119]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[123]);
  assign t[85] = ~(t[123] & t[91]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[124]);
  assign t[89] = ~(t[124] & t[92]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[120]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = t[32] ^ t[26];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = ~(t[114]);
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[114] ? x[24] : x[23];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[35];
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[120]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[114] ? x[40] : x[39];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = ~(t[77] & t[121]);
  assign t[54] = t[114] ? x[45] : x[44];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[124]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = ~(t[85] & t[125]);
  assign t[63] = t[18] ? x[59] : x[58];
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = ~(t[88] & t[126]);
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[89] & t[90]);
  assign t[68] = ~(t[119] & t[118]);
  assign t[69] = ~(t[127]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[93] & t[94]);
  assign t[74] = ~(t[95] & t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[132]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [139:0] x;
 output y;

 wire [397:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[2];
  assign t[153] = t[194] ^ x[10];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[27];
  assign t[159] = t[200] ^ x[32];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[35];
  assign t[161] = t[202] ^ x[38];
  assign t[162] = t[203] ^ x[43];
  assign t[163] = t[204] ^ x[48];
  assign t[164] = t[205] ^ x[51];
  assign t[165] = t[206] ^ x[54];
  assign t[166] = t[207] ^ x[57];
  assign t[167] = t[208] ^ x[62];
  assign t[168] = t[209] ^ x[67];
  assign t[169] = t[210] ^ x[70];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[73];
  assign t[171] = t[212] ^ x[76];
  assign t[172] = t[213] ^ x[79];
  assign t[173] = t[214] ^ x[82];
  assign t[174] = t[215] ^ x[85];
  assign t[175] = t[216] ^ x[88];
  assign t[176] = t[217] ^ x[91];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[97];
  assign t[179] = t[220] ^ x[100];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[106];
  assign t[182] = t[223] ^ x[109];
  assign t[183] = t[224] ^ x[112];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = t[226] ^ x[118];
  assign t[186] = t[227] ^ x[121];
  assign t[187] = t[228] ^ x[124];
  assign t[188] = t[229] ^ x[127];
  assign t[189] = t[230] ^ x[130];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[133];
  assign t[191] = t[232] ^ x[136];
  assign t[192] = t[233] ^ x[139];
  assign t[193] = (t[234] & ~t[235]);
  assign t[194] = (t[236] & ~t[237]);
  assign t[195] = (t[238] & ~t[239]);
  assign t[196] = (t[240] & ~t[241]);
  assign t[197] = (t[242] & ~t[243]);
  assign t[198] = (t[244] & ~t[245]);
  assign t[199] = (t[246] & ~t[247]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[248] & ~t[249]);
  assign t[201] = (t[250] & ~t[251]);
  assign t[202] = (t[252] & ~t[253]);
  assign t[203] = (t[254] & ~t[255]);
  assign t[204] = (t[256] & ~t[257]);
  assign t[205] = (t[258] & ~t[259]);
  assign t[206] = (t[260] & ~t[261]);
  assign t[207] = (t[262] & ~t[263]);
  assign t[208] = (t[264] & ~t[265]);
  assign t[209] = (t[266] & ~t[267]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[268] & ~t[269]);
  assign t[211] = (t[270] & ~t[271]);
  assign t[212] = (t[272] & ~t[273]);
  assign t[213] = (t[274] & ~t[275]);
  assign t[214] = (t[276] & ~t[277]);
  assign t[215] = (t[278] & ~t[279]);
  assign t[216] = (t[280] & ~t[281]);
  assign t[217] = (t[282] & ~t[283]);
  assign t[218] = (t[284] & ~t[285]);
  assign t[219] = (t[286] & ~t[287]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[288] & ~t[289]);
  assign t[221] = (t[290] & ~t[291]);
  assign t[222] = (t[292] & ~t[293]);
  assign t[223] = (t[294] & ~t[295]);
  assign t[224] = (t[296] & ~t[297]);
  assign t[225] = (t[298] & ~t[299]);
  assign t[226] = (t[300] & ~t[301]);
  assign t[227] = (t[302] & ~t[303]);
  assign t[228] = (t[304] & ~t[305]);
  assign t[229] = (t[306] & ~t[307]);
  assign t[22] = t[32] ^ t[26];
  assign t[230] = (t[308] & ~t[309]);
  assign t[231] = (t[310] & ~t[311]);
  assign t[232] = (t[312] & ~t[313]);
  assign t[233] = (t[314] & ~t[315]);
  assign t[234] = t[316] ^ x[2];
  assign t[235] = t[317] ^ x[1];
  assign t[236] = t[318] ^ x[10];
  assign t[237] = t[319] ^ x[9];
  assign t[238] = t[320] ^ x[13];
  assign t[239] = t[321] ^ x[12];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[16];
  assign t[241] = t[323] ^ x[15];
  assign t[242] = t[324] ^ x[19];
  assign t[243] = t[325] ^ x[18];
  assign t[244] = t[326] ^ x[22];
  assign t[245] = t[327] ^ x[21];
  assign t[246] = t[328] ^ x[27];
  assign t[247] = t[329] ^ x[26];
  assign t[248] = t[330] ^ x[32];
  assign t[249] = t[331] ^ x[31];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[35];
  assign t[251] = t[333] ^ x[34];
  assign t[252] = t[334] ^ x[38];
  assign t[253] = t[335] ^ x[37];
  assign t[254] = t[336] ^ x[43];
  assign t[255] = t[337] ^ x[42];
  assign t[256] = t[338] ^ x[48];
  assign t[257] = t[339] ^ x[47];
  assign t[258] = t[340] ^ x[51];
  assign t[259] = t[341] ^ x[50];
  assign t[25] = ~(t[114]);
  assign t[260] = t[342] ^ x[54];
  assign t[261] = t[343] ^ x[53];
  assign t[262] = t[344] ^ x[57];
  assign t[263] = t[345] ^ x[56];
  assign t[264] = t[346] ^ x[62];
  assign t[265] = t[347] ^ x[61];
  assign t[266] = t[348] ^ x[67];
  assign t[267] = t[349] ^ x[66];
  assign t[268] = t[350] ^ x[70];
  assign t[269] = t[351] ^ x[69];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[73];
  assign t[271] = t[353] ^ x[72];
  assign t[272] = t[354] ^ x[76];
  assign t[273] = t[355] ^ x[75];
  assign t[274] = t[356] ^ x[79];
  assign t[275] = t[357] ^ x[78];
  assign t[276] = t[358] ^ x[82];
  assign t[277] = t[359] ^ x[81];
  assign t[278] = t[360] ^ x[85];
  assign t[279] = t[361] ^ x[84];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[88];
  assign t[281] = t[363] ^ x[87];
  assign t[282] = t[364] ^ x[91];
  assign t[283] = t[365] ^ x[90];
  assign t[284] = t[366] ^ x[94];
  assign t[285] = t[367] ^ x[93];
  assign t[286] = t[368] ^ x[97];
  assign t[287] = t[369] ^ x[96];
  assign t[288] = t[370] ^ x[100];
  assign t[289] = t[371] ^ x[99];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[103];
  assign t[291] = t[373] ^ x[102];
  assign t[292] = t[374] ^ x[106];
  assign t[293] = t[375] ^ x[105];
  assign t[294] = t[376] ^ x[109];
  assign t[295] = t[377] ^ x[108];
  assign t[296] = t[378] ^ x[112];
  assign t[297] = t[379] ^ x[111];
  assign t[298] = t[380] ^ x[115];
  assign t[299] = t[381] ^ x[114];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[118];
  assign t[301] = t[383] ^ x[117];
  assign t[302] = t[384] ^ x[121];
  assign t[303] = t[385] ^ x[120];
  assign t[304] = t[386] ^ x[124];
  assign t[305] = t[387] ^ x[123];
  assign t[306] = t[388] ^ x[127];
  assign t[307] = t[389] ^ x[126];
  assign t[308] = t[390] ^ x[130];
  assign t[309] = t[391] ^ x[129];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[133];
  assign t[311] = t[393] ^ x[132];
  assign t[312] = t[394] ^ x[136];
  assign t[313] = t[395] ^ x[135];
  assign t[314] = t[396] ^ x[139];
  assign t[315] = t[397] ^ x[138];
  assign t[316] = (x[0]);
  assign t[317] = (x[0]);
  assign t[318] = (x[8]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[11]);
  assign t[321] = (x[11]);
  assign t[322] = (x[14]);
  assign t[323] = (x[14]);
  assign t[324] = (x[17]);
  assign t[325] = (x[17]);
  assign t[326] = (x[20]);
  assign t[327] = (x[20]);
  assign t[328] = (x[25]);
  assign t[329] = (x[25]);
  assign t[32] = t[114] ? x[24] : x[23];
  assign t[330] = (x[30]);
  assign t[331] = (x[30]);
  assign t[332] = (x[33]);
  assign t[333] = (x[33]);
  assign t[334] = (x[36]);
  assign t[335] = (x[36]);
  assign t[336] = (x[41]);
  assign t[337] = (x[41]);
  assign t[338] = (x[46]);
  assign t[339] = (x[46]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[49]);
  assign t[341] = (x[49]);
  assign t[342] = (x[52]);
  assign t[343] = (x[52]);
  assign t[344] = (x[55]);
  assign t[345] = (x[55]);
  assign t[346] = (x[60]);
  assign t[347] = (x[60]);
  assign t[348] = (x[65]);
  assign t[349] = (x[65]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[68]);
  assign t[351] = (x[68]);
  assign t[352] = (x[71]);
  assign t[353] = (x[71]);
  assign t[354] = (x[74]);
  assign t[355] = (x[74]);
  assign t[356] = (x[77]);
  assign t[357] = (x[77]);
  assign t[358] = (x[80]);
  assign t[359] = (x[80]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[83]);
  assign t[361] = (x[83]);
  assign t[362] = (x[86]);
  assign t[363] = (x[86]);
  assign t[364] = (x[89]);
  assign t[365] = (x[89]);
  assign t[366] = (x[92]);
  assign t[367] = (x[92]);
  assign t[368] = (x[95]);
  assign t[369] = (x[95]);
  assign t[36] = t[54] ^ t[35];
  assign t[370] = (x[98]);
  assign t[371] = (x[98]);
  assign t[372] = (x[101]);
  assign t[373] = (x[101]);
  assign t[374] = (x[104]);
  assign t[375] = (x[104]);
  assign t[376] = (x[107]);
  assign t[377] = (x[107]);
  assign t[378] = (x[110]);
  assign t[379] = (x[110]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[113]);
  assign t[381] = (x[113]);
  assign t[382] = (x[116]);
  assign t[383] = (x[116]);
  assign t[384] = (x[119]);
  assign t[385] = (x[119]);
  assign t[386] = (x[122]);
  assign t[387] = (x[122]);
  assign t[388] = (x[125]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[390] = (x[128]);
  assign t[391] = (x[128]);
  assign t[392] = (x[131]);
  assign t[393] = (x[131]);
  assign t[394] = (x[134]);
  assign t[395] = (x[134]);
  assign t[396] = (x[137]);
  assign t[397] = (x[137]);
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[120]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[114] ? x[40] : x[39];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = ~(t[77] & t[121]);
  assign t[54] = t[114] ? x[45] : x[44];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[124]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = ~(t[85] & t[125]);
  assign t[63] = t[18] ? x[59] : x[58];
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = ~(t[88] & t[126]);
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[89] & t[90]);
  assign t[68] = ~(t[119] & t[118]);
  assign t[69] = ~(t[127]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[93] & t[94]);
  assign t[74] = ~(t[95] & t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[132]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [139:0] x;
 output y;

 wire [388:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[2];
  assign t[144] = t[185] ^ x[10];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[27];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[32];
  assign t[151] = t[192] ^ x[35];
  assign t[152] = t[193] ^ x[38];
  assign t[153] = t[194] ^ x[43];
  assign t[154] = t[195] ^ x[48];
  assign t[155] = t[196] ^ x[51];
  assign t[156] = t[197] ^ x[54];
  assign t[157] = t[198] ^ x[57];
  assign t[158] = t[199] ^ x[62];
  assign t[159] = t[200] ^ x[67];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[70];
  assign t[161] = t[202] ^ x[73];
  assign t[162] = t[203] ^ x[76];
  assign t[163] = t[204] ^ x[79];
  assign t[164] = t[205] ^ x[82];
  assign t[165] = t[206] ^ x[85];
  assign t[166] = t[207] ^ x[88];
  assign t[167] = t[208] ^ x[91];
  assign t[168] = t[209] ^ x[94];
  assign t[169] = t[210] ^ x[97];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[100];
  assign t[171] = t[212] ^ x[103];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[109];
  assign t[174] = t[215] ^ x[112];
  assign t[175] = t[216] ^ x[115];
  assign t[176] = t[217] ^ x[118];
  assign t[177] = t[218] ^ x[121];
  assign t[178] = t[219] ^ x[124];
  assign t[179] = t[220] ^ x[127];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[130];
  assign t[181] = t[222] ^ x[133];
  assign t[182] = t[223] ^ x[136];
  assign t[183] = t[224] ^ x[139];
  assign t[184] = (t[225] & ~t[226]);
  assign t[185] = (t[227] & ~t[228]);
  assign t[186] = (t[229] & ~t[230]);
  assign t[187] = (t[231] & ~t[232]);
  assign t[188] = (t[233] & ~t[234]);
  assign t[189] = (t[235] & ~t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[237] & ~t[238]);
  assign t[191] = (t[239] & ~t[240]);
  assign t[192] = (t[241] & ~t[242]);
  assign t[193] = (t[243] & ~t[244]);
  assign t[194] = (t[245] & ~t[246]);
  assign t[195] = (t[247] & ~t[248]);
  assign t[196] = (t[249] & ~t[250]);
  assign t[197] = (t[251] & ~t[252]);
  assign t[198] = (t[253] & ~t[254]);
  assign t[199] = (t[255] & ~t[256]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[257] & ~t[258]);
  assign t[201] = (t[259] & ~t[260]);
  assign t[202] = (t[261] & ~t[262]);
  assign t[203] = (t[263] & ~t[264]);
  assign t[204] = (t[265] & ~t[266]);
  assign t[205] = (t[267] & ~t[268]);
  assign t[206] = (t[269] & ~t[270]);
  assign t[207] = (t[271] & ~t[272]);
  assign t[208] = (t[273] & ~t[274]);
  assign t[209] = (t[275] & ~t[276]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[277] & ~t[278]);
  assign t[211] = (t[279] & ~t[280]);
  assign t[212] = (t[281] & ~t[282]);
  assign t[213] = (t[283] & ~t[284]);
  assign t[214] = (t[285] & ~t[286]);
  assign t[215] = (t[287] & ~t[288]);
  assign t[216] = (t[289] & ~t[290]);
  assign t[217] = (t[291] & ~t[292]);
  assign t[218] = (t[293] & ~t[294]);
  assign t[219] = (t[295] & ~t[296]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[297] & ~t[298]);
  assign t[221] = (t[299] & ~t[300]);
  assign t[222] = (t[301] & ~t[302]);
  assign t[223] = (t[303] & ~t[304]);
  assign t[224] = (t[305] & ~t[306]);
  assign t[225] = t[307] ^ x[2];
  assign t[226] = t[308] ^ x[1];
  assign t[227] = t[309] ^ x[10];
  assign t[228] = t[310] ^ x[9];
  assign t[229] = t[311] ^ x[13];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[312] ^ x[12];
  assign t[231] = t[313] ^ x[16];
  assign t[232] = t[314] ^ x[15];
  assign t[233] = t[315] ^ x[19];
  assign t[234] = t[316] ^ x[18];
  assign t[235] = t[317] ^ x[22];
  assign t[236] = t[318] ^ x[21];
  assign t[237] = t[319] ^ x[27];
  assign t[238] = t[320] ^ x[26];
  assign t[239] = t[321] ^ x[32];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[31];
  assign t[241] = t[323] ^ x[35];
  assign t[242] = t[324] ^ x[34];
  assign t[243] = t[325] ^ x[38];
  assign t[244] = t[326] ^ x[37];
  assign t[245] = t[327] ^ x[43];
  assign t[246] = t[328] ^ x[42];
  assign t[247] = t[329] ^ x[48];
  assign t[248] = t[330] ^ x[47];
  assign t[249] = t[331] ^ x[51];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[50];
  assign t[251] = t[333] ^ x[54];
  assign t[252] = t[334] ^ x[53];
  assign t[253] = t[335] ^ x[57];
  assign t[254] = t[336] ^ x[56];
  assign t[255] = t[337] ^ x[62];
  assign t[256] = t[338] ^ x[61];
  assign t[257] = t[339] ^ x[67];
  assign t[258] = t[340] ^ x[66];
  assign t[259] = t[341] ^ x[70];
  assign t[25] = ~(t[105]);
  assign t[260] = t[342] ^ x[69];
  assign t[261] = t[343] ^ x[73];
  assign t[262] = t[344] ^ x[72];
  assign t[263] = t[345] ^ x[76];
  assign t[264] = t[346] ^ x[75];
  assign t[265] = t[347] ^ x[79];
  assign t[266] = t[348] ^ x[78];
  assign t[267] = t[349] ^ x[82];
  assign t[268] = t[350] ^ x[81];
  assign t[269] = t[351] ^ x[85];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[84];
  assign t[271] = t[353] ^ x[88];
  assign t[272] = t[354] ^ x[87];
  assign t[273] = t[355] ^ x[91];
  assign t[274] = t[356] ^ x[90];
  assign t[275] = t[357] ^ x[94];
  assign t[276] = t[358] ^ x[93];
  assign t[277] = t[359] ^ x[97];
  assign t[278] = t[360] ^ x[96];
  assign t[279] = t[361] ^ x[100];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[99];
  assign t[281] = t[363] ^ x[103];
  assign t[282] = t[364] ^ x[102];
  assign t[283] = t[365] ^ x[106];
  assign t[284] = t[366] ^ x[105];
  assign t[285] = t[367] ^ x[109];
  assign t[286] = t[368] ^ x[108];
  assign t[287] = t[369] ^ x[112];
  assign t[288] = t[370] ^ x[111];
  assign t[289] = t[371] ^ x[115];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[114];
  assign t[291] = t[373] ^ x[118];
  assign t[292] = t[374] ^ x[117];
  assign t[293] = t[375] ^ x[121];
  assign t[294] = t[376] ^ x[120];
  assign t[295] = t[377] ^ x[124];
  assign t[296] = t[378] ^ x[123];
  assign t[297] = t[379] ^ x[127];
  assign t[298] = t[380] ^ x[126];
  assign t[299] = t[381] ^ x[130];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[129];
  assign t[301] = t[383] ^ x[133];
  assign t[302] = t[384] ^ x[132];
  assign t[303] = t[385] ^ x[136];
  assign t[304] = t[386] ^ x[135];
  assign t[305] = t[387] ^ x[139];
  assign t[306] = t[388] ^ x[138];
  assign t[307] = (x[0]);
  assign t[308] = (x[0]);
  assign t[309] = (x[8]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[11]);
  assign t[312] = (x[11]);
  assign t[313] = (x[14]);
  assign t[314] = (x[14]);
  assign t[315] = (x[17]);
  assign t[316] = (x[17]);
  assign t[317] = (x[20]);
  assign t[318] = (x[20]);
  assign t[319] = (x[25]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[25]);
  assign t[321] = (x[30]);
  assign t[322] = (x[30]);
  assign t[323] = (x[33]);
  assign t[324] = (x[33]);
  assign t[325] = (x[36]);
  assign t[326] = (x[36]);
  assign t[327] = (x[41]);
  assign t[328] = (x[41]);
  assign t[329] = (x[46]);
  assign t[32] = t[105] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[49]);
  assign t[332] = (x[49]);
  assign t[333] = (x[52]);
  assign t[334] = (x[52]);
  assign t[335] = (x[55]);
  assign t[336] = (x[55]);
  assign t[337] = (x[60]);
  assign t[338] = (x[60]);
  assign t[339] = (x[65]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[68]);
  assign t[342] = (x[68]);
  assign t[343] = (x[71]);
  assign t[344] = (x[71]);
  assign t[345] = (x[74]);
  assign t[346] = (x[74]);
  assign t[347] = (x[77]);
  assign t[348] = (x[77]);
  assign t[349] = (x[80]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[80]);
  assign t[351] = (x[83]);
  assign t[352] = (x[83]);
  assign t[353] = (x[86]);
  assign t[354] = (x[86]);
  assign t[355] = (x[89]);
  assign t[356] = (x[89]);
  assign t[357] = (x[92]);
  assign t[358] = (x[92]);
  assign t[359] = (x[95]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[95]);
  assign t[361] = (x[98]);
  assign t[362] = (x[98]);
  assign t[363] = (x[101]);
  assign t[364] = (x[101]);
  assign t[365] = (x[104]);
  assign t[366] = (x[104]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[54] ^ t[35];
  assign t[370] = (x[110]);
  assign t[371] = (x[113]);
  assign t[372] = (x[113]);
  assign t[373] = (x[116]);
  assign t[374] = (x[116]);
  assign t[375] = (x[119]);
  assign t[376] = (x[119]);
  assign t[377] = (x[122]);
  assign t[378] = (x[122]);
  assign t[379] = (x[125]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[128]);
  assign t[382] = (x[128]);
  assign t[383] = (x[131]);
  assign t[384] = (x[131]);
  assign t[385] = (x[134]);
  assign t[386] = (x[134]);
  assign t[387] = (x[137]);
  assign t[388] = (x[137]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[111];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[105] ? x[40] : x[39];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = t[76] | t[112];
  assign t[54] = t[105] ? x[45] : x[44];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[78] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[80] | t[115];
  assign t[61] = ~(t[81] & t[82]);
  assign t[62] = t[83] | t[116];
  assign t[63] = t[18] ? x[59] : x[58];
  assign t[64] = ~(t[84] & t[85]);
  assign t[65] = t[86] | t[117];
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[87] & t[88]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[89] | t[69]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = t[92] | t[121];
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[93] | t[74]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind251(x, y);
 input [139:0] x;
 output y;

 wire [388:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[2];
  assign t[144] = t[185] ^ x[10];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[27];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[32];
  assign t[151] = t[192] ^ x[35];
  assign t[152] = t[193] ^ x[38];
  assign t[153] = t[194] ^ x[43];
  assign t[154] = t[195] ^ x[48];
  assign t[155] = t[196] ^ x[51];
  assign t[156] = t[197] ^ x[54];
  assign t[157] = t[198] ^ x[57];
  assign t[158] = t[199] ^ x[62];
  assign t[159] = t[200] ^ x[67];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[70];
  assign t[161] = t[202] ^ x[73];
  assign t[162] = t[203] ^ x[76];
  assign t[163] = t[204] ^ x[79];
  assign t[164] = t[205] ^ x[82];
  assign t[165] = t[206] ^ x[85];
  assign t[166] = t[207] ^ x[88];
  assign t[167] = t[208] ^ x[91];
  assign t[168] = t[209] ^ x[94];
  assign t[169] = t[210] ^ x[97];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[100];
  assign t[171] = t[212] ^ x[103];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[109];
  assign t[174] = t[215] ^ x[112];
  assign t[175] = t[216] ^ x[115];
  assign t[176] = t[217] ^ x[118];
  assign t[177] = t[218] ^ x[121];
  assign t[178] = t[219] ^ x[124];
  assign t[179] = t[220] ^ x[127];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[130];
  assign t[181] = t[222] ^ x[133];
  assign t[182] = t[223] ^ x[136];
  assign t[183] = t[224] ^ x[139];
  assign t[184] = (t[225] & ~t[226]);
  assign t[185] = (t[227] & ~t[228]);
  assign t[186] = (t[229] & ~t[230]);
  assign t[187] = (t[231] & ~t[232]);
  assign t[188] = (t[233] & ~t[234]);
  assign t[189] = (t[235] & ~t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[237] & ~t[238]);
  assign t[191] = (t[239] & ~t[240]);
  assign t[192] = (t[241] & ~t[242]);
  assign t[193] = (t[243] & ~t[244]);
  assign t[194] = (t[245] & ~t[246]);
  assign t[195] = (t[247] & ~t[248]);
  assign t[196] = (t[249] & ~t[250]);
  assign t[197] = (t[251] & ~t[252]);
  assign t[198] = (t[253] & ~t[254]);
  assign t[199] = (t[255] & ~t[256]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[257] & ~t[258]);
  assign t[201] = (t[259] & ~t[260]);
  assign t[202] = (t[261] & ~t[262]);
  assign t[203] = (t[263] & ~t[264]);
  assign t[204] = (t[265] & ~t[266]);
  assign t[205] = (t[267] & ~t[268]);
  assign t[206] = (t[269] & ~t[270]);
  assign t[207] = (t[271] & ~t[272]);
  assign t[208] = (t[273] & ~t[274]);
  assign t[209] = (t[275] & ~t[276]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[277] & ~t[278]);
  assign t[211] = (t[279] & ~t[280]);
  assign t[212] = (t[281] & ~t[282]);
  assign t[213] = (t[283] & ~t[284]);
  assign t[214] = (t[285] & ~t[286]);
  assign t[215] = (t[287] & ~t[288]);
  assign t[216] = (t[289] & ~t[290]);
  assign t[217] = (t[291] & ~t[292]);
  assign t[218] = (t[293] & ~t[294]);
  assign t[219] = (t[295] & ~t[296]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[297] & ~t[298]);
  assign t[221] = (t[299] & ~t[300]);
  assign t[222] = (t[301] & ~t[302]);
  assign t[223] = (t[303] & ~t[304]);
  assign t[224] = (t[305] & ~t[306]);
  assign t[225] = t[307] ^ x[2];
  assign t[226] = t[308] ^ x[1];
  assign t[227] = t[309] ^ x[10];
  assign t[228] = t[310] ^ x[9];
  assign t[229] = t[311] ^ x[13];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[312] ^ x[12];
  assign t[231] = t[313] ^ x[16];
  assign t[232] = t[314] ^ x[15];
  assign t[233] = t[315] ^ x[19];
  assign t[234] = t[316] ^ x[18];
  assign t[235] = t[317] ^ x[22];
  assign t[236] = t[318] ^ x[21];
  assign t[237] = t[319] ^ x[27];
  assign t[238] = t[320] ^ x[26];
  assign t[239] = t[321] ^ x[32];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[240] = t[322] ^ x[31];
  assign t[241] = t[323] ^ x[35];
  assign t[242] = t[324] ^ x[34];
  assign t[243] = t[325] ^ x[38];
  assign t[244] = t[326] ^ x[37];
  assign t[245] = t[327] ^ x[43];
  assign t[246] = t[328] ^ x[42];
  assign t[247] = t[329] ^ x[48];
  assign t[248] = t[330] ^ x[47];
  assign t[249] = t[331] ^ x[51];
  assign t[24] = x[4] ? t[36] : t[35];
  assign t[250] = t[332] ^ x[50];
  assign t[251] = t[333] ^ x[54];
  assign t[252] = t[334] ^ x[53];
  assign t[253] = t[335] ^ x[57];
  assign t[254] = t[336] ^ x[56];
  assign t[255] = t[337] ^ x[62];
  assign t[256] = t[338] ^ x[61];
  assign t[257] = t[339] ^ x[67];
  assign t[258] = t[340] ^ x[66];
  assign t[259] = t[341] ^ x[70];
  assign t[25] = ~(t[105]);
  assign t[260] = t[342] ^ x[69];
  assign t[261] = t[343] ^ x[73];
  assign t[262] = t[344] ^ x[72];
  assign t[263] = t[345] ^ x[76];
  assign t[264] = t[346] ^ x[75];
  assign t[265] = t[347] ^ x[79];
  assign t[266] = t[348] ^ x[78];
  assign t[267] = t[349] ^ x[82];
  assign t[268] = t[350] ^ x[81];
  assign t[269] = t[351] ^ x[85];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[352] ^ x[84];
  assign t[271] = t[353] ^ x[88];
  assign t[272] = t[354] ^ x[87];
  assign t[273] = t[355] ^ x[91];
  assign t[274] = t[356] ^ x[90];
  assign t[275] = t[357] ^ x[94];
  assign t[276] = t[358] ^ x[93];
  assign t[277] = t[359] ^ x[97];
  assign t[278] = t[360] ^ x[96];
  assign t[279] = t[361] ^ x[100];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[362] ^ x[99];
  assign t[281] = t[363] ^ x[103];
  assign t[282] = t[364] ^ x[102];
  assign t[283] = t[365] ^ x[106];
  assign t[284] = t[366] ^ x[105];
  assign t[285] = t[367] ^ x[109];
  assign t[286] = t[368] ^ x[108];
  assign t[287] = t[369] ^ x[112];
  assign t[288] = t[370] ^ x[111];
  assign t[289] = t[371] ^ x[115];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[114];
  assign t[291] = t[373] ^ x[118];
  assign t[292] = t[374] ^ x[117];
  assign t[293] = t[375] ^ x[121];
  assign t[294] = t[376] ^ x[120];
  assign t[295] = t[377] ^ x[124];
  assign t[296] = t[378] ^ x[123];
  assign t[297] = t[379] ^ x[127];
  assign t[298] = t[380] ^ x[126];
  assign t[299] = t[381] ^ x[130];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[129];
  assign t[301] = t[383] ^ x[133];
  assign t[302] = t[384] ^ x[132];
  assign t[303] = t[385] ^ x[136];
  assign t[304] = t[386] ^ x[135];
  assign t[305] = t[387] ^ x[139];
  assign t[306] = t[388] ^ x[138];
  assign t[307] = (x[0]);
  assign t[308] = (x[0]);
  assign t[309] = (x[8]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[11]);
  assign t[312] = (x[11]);
  assign t[313] = (x[14]);
  assign t[314] = (x[14]);
  assign t[315] = (x[17]);
  assign t[316] = (x[17]);
  assign t[317] = (x[20]);
  assign t[318] = (x[20]);
  assign t[319] = (x[25]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[25]);
  assign t[321] = (x[30]);
  assign t[322] = (x[30]);
  assign t[323] = (x[33]);
  assign t[324] = (x[33]);
  assign t[325] = (x[36]);
  assign t[326] = (x[36]);
  assign t[327] = (x[41]);
  assign t[328] = (x[41]);
  assign t[329] = (x[46]);
  assign t[32] = t[105] ? x[24] : x[23];
  assign t[330] = (x[46]);
  assign t[331] = (x[49]);
  assign t[332] = (x[49]);
  assign t[333] = (x[52]);
  assign t[334] = (x[52]);
  assign t[335] = (x[55]);
  assign t[336] = (x[55]);
  assign t[337] = (x[60]);
  assign t[338] = (x[60]);
  assign t[339] = (x[65]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[65]);
  assign t[341] = (x[68]);
  assign t[342] = (x[68]);
  assign t[343] = (x[71]);
  assign t[344] = (x[71]);
  assign t[345] = (x[74]);
  assign t[346] = (x[74]);
  assign t[347] = (x[77]);
  assign t[348] = (x[77]);
  assign t[349] = (x[80]);
  assign t[34] = t[50] ^ t[51];
  assign t[350] = (x[80]);
  assign t[351] = (x[83]);
  assign t[352] = (x[83]);
  assign t[353] = (x[86]);
  assign t[354] = (x[86]);
  assign t[355] = (x[89]);
  assign t[356] = (x[89]);
  assign t[357] = (x[92]);
  assign t[358] = (x[92]);
  assign t[359] = (x[95]);
  assign t[35] = ~(t[52] & t[53]);
  assign t[360] = (x[95]);
  assign t[361] = (x[98]);
  assign t[362] = (x[98]);
  assign t[363] = (x[101]);
  assign t[364] = (x[101]);
  assign t[365] = (x[104]);
  assign t[366] = (x[104]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[54] ^ t[35];
  assign t[370] = (x[110]);
  assign t[371] = (x[113]);
  assign t[372] = (x[113]);
  assign t[373] = (x[116]);
  assign t[374] = (x[116]);
  assign t[375] = (x[119]);
  assign t[376] = (x[119]);
  assign t[377] = (x[122]);
  assign t[378] = (x[122]);
  assign t[379] = (x[125]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[380] = (x[125]);
  assign t[381] = (x[128]);
  assign t[382] = (x[128]);
  assign t[383] = (x[131]);
  assign t[384] = (x[131]);
  assign t[385] = (x[134]);
  assign t[386] = (x[134]);
  assign t[387] = (x[137]);
  assign t[388] = (x[137]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[58] ? x[29] : x[28];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[111];
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[105] ? x[40] : x[39];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = t[76] | t[112];
  assign t[54] = t[105] ? x[45] : x[44];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[78] & t[79]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[80] | t[115];
  assign t[61] = ~(t[81] & t[82]);
  assign t[62] = t[83] | t[116];
  assign t[63] = t[18] ? x[59] : x[58];
  assign t[64] = ~(t[84] & t[85]);
  assign t[65] = t[86] | t[117];
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[87] & t[88]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[89] | t[69]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = t[92] | t[121];
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[93] | t[74]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [139:0] x;
 output y;

 wire [484:0] t;
  assign t[0] = t[1] ? t[2] : t[198];
  assign t[100] = ~(t[140] | t[141]);
  assign t[101] = t[137] ? x[81] : x[80];
  assign t[102] = ~(t[142] & t[106]);
  assign t[103] = ~(t[221]);
  assign t[104] = ~(t[210] | t[211]);
  assign t[105] = ~(t[125] | t[50]);
  assign t[106] = ~(t[143] | t[139]);
  assign t[107] = ~(t[222]);
  assign t[108] = ~(t[223]);
  assign t[109] = ~(t[144] | t[145]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[146] | t[147]);
  assign t[111] = ~(t[224] | t[148]);
  assign t[112] = t[30] ? x[95] : x[94];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[225]);
  assign t[115] = ~(t[226]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[227] | t[155]);
  assign t[119] = t[137] ? x[106] : x[105];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[156] & t[157]);
  assign t[121] = ~(t[158] & t[159]);
  assign t[122] = ~(t[160] & t[159]);
  assign t[123] = ~(x[4] & t[161]);
  assign t[124] = ~(t[162] & t[159]);
  assign t[125] = ~(t[79] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[123] & t[166]);
  assign t[128] = t[202] & t[167];
  assign t[129] = t[158] | t[160];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[199] ? t[123] : t[124];
  assign t[131] = ~(t[228]);
  assign t[132] = ~(t[215] | t[216]);
  assign t[133] = ~(t[168] & t[169]);
  assign t[134] = t[139] | t[170];
  assign t[135] = ~(t[229]);
  assign t[136] = ~(t[217] | t[218]);
  assign t[137] = ~(t[48]);
  assign t[138] = ~(t[31] & t[169]);
  assign t[139] = ~(t[164] | t[171]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[230]);
  assign t[141] = ~(t[219] | t[220]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[173]);
  assign t[144] = ~(t[231]);
  assign t[145] = ~(t[222] | t[223]);
  assign t[146] = ~(t[232]);
  assign t[147] = ~(t[233]);
  assign t[148] = ~(t[174] | t[175]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[225] | t[226]);
  assign t[153] = ~(t[235]);
  assign t[154] = ~(t[236]);
  assign t[155] = ~(t[179] | t[180]);
  assign t[156] = ~(t[181] | t[182]);
  assign t[157] = ~(t[183]);
  assign t[158] = ~(x[4] | t[200]);
  assign t[159] = ~(t[202]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[4] & t[200];
  assign t[161] = ~(t[200] | t[202]);
  assign t[162] = ~(x[4] | t[184]);
  assign t[163] = t[199] ? t[121] : t[122];
  assign t[164] = ~(t[79]);
  assign t[165] = t[199] ? t[124] : t[185];
  assign t[166] = ~(t[202] & t[162]);
  assign t[167] = ~(t[79] | t[199]);
  assign t[168] = ~(t[167] & t[186]);
  assign t[169] = ~(t[187] & t[188]);
  assign t[16] = ~(t[199] & t[200]);
  assign t[170] = ~(t[164] | t[189]);
  assign t[171] = t[199] ? t[166] : t[123];
  assign t[172] = ~(t[164] | t[190]);
  assign t[173] = ~(t[181] | t[177]);
  assign t[174] = ~(t[237]);
  assign t[175] = ~(t[232] | t[233]);
  assign t[176] = ~(t[164] | t[191]);
  assign t[177] = ~(t[164] | t[192]);
  assign t[178] = ~(t[31]);
  assign t[179] = ~(t[238]);
  assign t[17] = ~(t[201] & t[202]);
  assign t[180] = ~(t[235] | t[236]);
  assign t[181] = ~(t[164] | t[193]);
  assign t[182] = ~(t[194] & t[31]);
  assign t[183] = ~(t[164] | t[195]);
  assign t[184] = ~(t[200]);
  assign t[185] = ~(x[4] & t[187]);
  assign t[186] = ~(t[166] & t[185]);
  assign t[187] = ~(t[200] | t[159]);
  assign t[188] = t[164] & t[199];
  assign t[189] = t[199] ? t[196] : t[122];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[199] ? t[197] : t[121];
  assign t[191] = t[199] ? t[123] : t[166];
  assign t[192] = t[199] ? t[122] : t[196];
  assign t[193] = t[199] ? t[185] : t[124];
  assign t[194] = ~(t[172] | t[51]);
  assign t[195] = t[199] ? t[121] : t[197];
  assign t[196] = ~(t[158] & t[202]);
  assign t[197] = ~(t[160] & t[202]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = t[280] ^ x[2];
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[281] ^ x[10];
  assign t[241] = t[282] ^ x[13];
  assign t[242] = t[283] ^ x[16];
  assign t[243] = t[284] ^ x[19];
  assign t[244] = t[285] ^ x[22];
  assign t[245] = t[286] ^ x[25];
  assign t[246] = t[287] ^ x[28];
  assign t[247] = t[288] ^ x[31];
  assign t[248] = t[289] ^ x[34];
  assign t[249] = t[290] ^ x[39];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[291] ^ x[42];
  assign t[251] = t[292] ^ x[45];
  assign t[252] = t[293] ^ x[48];
  assign t[253] = t[294] ^ x[53];
  assign t[254] = t[295] ^ x[56];
  assign t[255] = t[296] ^ x[59];
  assign t[256] = t[297] ^ x[62];
  assign t[257] = t[298] ^ x[65];
  assign t[258] = t[299] ^ x[68];
  assign t[259] = t[300] ^ x[71];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[301] ^ x[76];
  assign t[261] = t[302] ^ x[79];
  assign t[262] = t[303] ^ x[84];
  assign t[263] = t[304] ^ x[87];
  assign t[264] = t[305] ^ x[90];
  assign t[265] = t[306] ^ x[93];
  assign t[266] = t[307] ^ x[98];
  assign t[267] = t[308] ^ x[101];
  assign t[268] = t[309] ^ x[104];
  assign t[269] = t[310] ^ x[109];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[311] ^ x[112];
  assign t[271] = t[312] ^ x[115];
  assign t[272] = t[313] ^ x[118];
  assign t[273] = t[314] ^ x[121];
  assign t[274] = t[315] ^ x[124];
  assign t[275] = t[316] ^ x[127];
  assign t[276] = t[317] ^ x[130];
  assign t[277] = t[318] ^ x[133];
  assign t[278] = t[319] ^ x[136];
  assign t[279] = t[320] ^ x[139];
  assign t[27] = ~(t[26] ^ t[43]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = (t[347] & ~t[348]);
  assign t[294] = (t[349] & ~t[350]);
  assign t[295] = (t[351] & ~t[352]);
  assign t[296] = (t[353] & ~t[354]);
  assign t[297] = (t[355] & ~t[356]);
  assign t[298] = (t[357] & ~t[358]);
  assign t[299] = (t[359] & ~t[360]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[361] & ~t[362]);
  assign t[301] = (t[363] & ~t[364]);
  assign t[302] = (t[365] & ~t[366]);
  assign t[303] = (t[367] & ~t[368]);
  assign t[304] = (t[369] & ~t[370]);
  assign t[305] = (t[371] & ~t[372]);
  assign t[306] = (t[373] & ~t[374]);
  assign t[307] = (t[375] & ~t[376]);
  assign t[308] = (t[377] & ~t[378]);
  assign t[309] = (t[379] & ~t[380]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[381] & ~t[382]);
  assign t[311] = (t[383] & ~t[384]);
  assign t[312] = (t[385] & ~t[386]);
  assign t[313] = (t[387] & ~t[388]);
  assign t[314] = (t[389] & ~t[390]);
  assign t[315] = (t[391] & ~t[392]);
  assign t[316] = (t[393] & ~t[394]);
  assign t[317] = (t[395] & ~t[396]);
  assign t[318] = (t[397] & ~t[398]);
  assign t[319] = (t[399] & ~t[400]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[401] & ~t[402]);
  assign t[321] = t[403] ^ x[2];
  assign t[322] = t[404] ^ x[1];
  assign t[323] = t[405] ^ x[10];
  assign t[324] = t[406] ^ x[9];
  assign t[325] = t[407] ^ x[13];
  assign t[326] = t[408] ^ x[12];
  assign t[327] = t[409] ^ x[16];
  assign t[328] = t[410] ^ x[15];
  assign t[329] = t[411] ^ x[19];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[18];
  assign t[331] = t[413] ^ x[22];
  assign t[332] = t[414] ^ x[21];
  assign t[333] = t[415] ^ x[25];
  assign t[334] = t[416] ^ x[24];
  assign t[335] = t[417] ^ x[28];
  assign t[336] = t[418] ^ x[27];
  assign t[337] = t[419] ^ x[31];
  assign t[338] = t[420] ^ x[30];
  assign t[339] = t[421] ^ x[34];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[33];
  assign t[341] = t[423] ^ x[39];
  assign t[342] = t[424] ^ x[38];
  assign t[343] = t[425] ^ x[42];
  assign t[344] = t[426] ^ x[41];
  assign t[345] = t[427] ^ x[45];
  assign t[346] = t[428] ^ x[44];
  assign t[347] = t[429] ^ x[48];
  assign t[348] = t[430] ^ x[47];
  assign t[349] = t[431] ^ x[53];
  assign t[34] = ~(t[203] | t[55]);
  assign t[350] = t[432] ^ x[52];
  assign t[351] = t[433] ^ x[56];
  assign t[352] = t[434] ^ x[55];
  assign t[353] = t[435] ^ x[59];
  assign t[354] = t[436] ^ x[58];
  assign t[355] = t[437] ^ x[62];
  assign t[356] = t[438] ^ x[61];
  assign t[357] = t[439] ^ x[65];
  assign t[358] = t[440] ^ x[64];
  assign t[359] = t[441] ^ x[68];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[442] ^ x[67];
  assign t[361] = t[443] ^ x[71];
  assign t[362] = t[444] ^ x[70];
  assign t[363] = t[445] ^ x[76];
  assign t[364] = t[446] ^ x[75];
  assign t[365] = t[447] ^ x[79];
  assign t[366] = t[448] ^ x[78];
  assign t[367] = t[449] ^ x[84];
  assign t[368] = t[450] ^ x[83];
  assign t[369] = t[451] ^ x[87];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[452] ^ x[86];
  assign t[371] = t[453] ^ x[90];
  assign t[372] = t[454] ^ x[89];
  assign t[373] = t[455] ^ x[93];
  assign t[374] = t[456] ^ x[92];
  assign t[375] = t[457] ^ x[98];
  assign t[376] = t[458] ^ x[97];
  assign t[377] = t[459] ^ x[101];
  assign t[378] = t[460] ^ x[100];
  assign t[379] = t[461] ^ x[104];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[462] ^ x[103];
  assign t[381] = t[463] ^ x[109];
  assign t[382] = t[464] ^ x[108];
  assign t[383] = t[465] ^ x[112];
  assign t[384] = t[466] ^ x[111];
  assign t[385] = t[467] ^ x[115];
  assign t[386] = t[468] ^ x[114];
  assign t[387] = t[469] ^ x[118];
  assign t[388] = t[470] ^ x[117];
  assign t[389] = t[471] ^ x[121];
  assign t[38] = ~(t[39] ^ t[62]);
  assign t[390] = t[472] ^ x[120];
  assign t[391] = t[473] ^ x[124];
  assign t[392] = t[474] ^ x[123];
  assign t[393] = t[475] ^ x[127];
  assign t[394] = t[476] ^ x[126];
  assign t[395] = t[477] ^ x[130];
  assign t[396] = t[478] ^ x[129];
  assign t[397] = t[479] ^ x[133];
  assign t[398] = t[480] ^ x[132];
  assign t[399] = t[481] ^ x[136];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[135];
  assign t[401] = t[483] ^ x[139];
  assign t[402] = t[484] ^ x[138];
  assign t[403] = (x[0]);
  assign t[404] = (x[0]);
  assign t[405] = (x[8]);
  assign t[406] = (x[8]);
  assign t[407] = (x[11]);
  assign t[408] = (x[11]);
  assign t[409] = (x[14]);
  assign t[40] = ~(t[44] ^ t[65]);
  assign t[410] = (x[14]);
  assign t[411] = (x[17]);
  assign t[412] = (x[17]);
  assign t[413] = (x[20]);
  assign t[414] = (x[20]);
  assign t[415] = (x[23]);
  assign t[416] = (x[23]);
  assign t[417] = (x[26]);
  assign t[418] = (x[26]);
  assign t[419] = (x[29]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[29]);
  assign t[421] = (x[32]);
  assign t[422] = (x[32]);
  assign t[423] = (x[37]);
  assign t[424] = (x[37]);
  assign t[425] = (x[40]);
  assign t[426] = (x[40]);
  assign t[427] = (x[43]);
  assign t[428] = (x[43]);
  assign t[429] = (x[46]);
  assign t[42] = ~(t[204] | t[68]);
  assign t[430] = (x[46]);
  assign t[431] = (x[51]);
  assign t[432] = (x[51]);
  assign t[433] = (x[54]);
  assign t[434] = (x[54]);
  assign t[435] = (x[57]);
  assign t[436] = (x[57]);
  assign t[437] = (x[60]);
  assign t[438] = (x[60]);
  assign t[439] = (x[63]);
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[440] = (x[63]);
  assign t[441] = (x[66]);
  assign t[442] = (x[66]);
  assign t[443] = (x[69]);
  assign t[444] = (x[69]);
  assign t[445] = (x[74]);
  assign t[446] = (x[74]);
  assign t[447] = (x[77]);
  assign t[448] = (x[77]);
  assign t[449] = (x[82]);
  assign t[44] = ~(t[71] | t[72]);
  assign t[450] = (x[82]);
  assign t[451] = (x[85]);
  assign t[452] = (x[85]);
  assign t[453] = (x[88]);
  assign t[454] = (x[88]);
  assign t[455] = (x[91]);
  assign t[456] = (x[91]);
  assign t[457] = (x[96]);
  assign t[458] = (x[96]);
  assign t[459] = (x[99]);
  assign t[45] = ~(t[73] ^ t[74]);
  assign t[460] = (x[99]);
  assign t[461] = (x[102]);
  assign t[462] = (x[102]);
  assign t[463] = (x[107]);
  assign t[464] = (x[107]);
  assign t[465] = (x[110]);
  assign t[466] = (x[110]);
  assign t[467] = (x[113]);
  assign t[468] = (x[113]);
  assign t[469] = (x[116]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[116]);
  assign t[471] = (x[119]);
  assign t[472] = (x[119]);
  assign t[473] = (x[122]);
  assign t[474] = (x[122]);
  assign t[475] = (x[125]);
  assign t[476] = (x[125]);
  assign t[477] = (x[128]);
  assign t[478] = (x[128]);
  assign t[479] = (x[131]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[131]);
  assign t[481] = (x[134]);
  assign t[482] = (x[134]);
  assign t[483] = (x[137]);
  assign t[484] = (x[137]);
  assign t[48] = ~(t[201]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = ~(t[82] & t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[205]);
  assign t[54] = ~(t[206]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[207] | t[90]);
  assign t[58] = t[91] ? x[36] : x[35];
  assign t[59] = ~(t[92] & t[84]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[93] | t[94]);
  assign t[61] = ~(t[208] | t[95]);
  assign t[62] = ~(t[96] ^ t[97]);
  assign t[63] = ~(t[98] | t[99]);
  assign t[64] = ~(t[209] | t[100]);
  assign t[65] = ~(t[101] ^ t[102]);
  assign t[66] = ~(t[210]);
  assign t[67] = ~(t[211]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = t[30] ? x[50] : x[49];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[212] | t[109]);
  assign t[73] = ~(t[110] | t[111]);
  assign t[74] = ~(t[112] ^ t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[213] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[201]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[199] ? t[122] : t[121];
  assign t[81] = t[199] ? t[124] : t[123];
  assign t[82] = ~(t[125] | t[126]);
  assign t[83] = ~(t[79] & t[127]);
  assign t[84] = ~(t[128] & t[129]);
  assign t[85] = t[79] | t[130];
  assign t[86] = ~(t[214]);
  assign t[87] = ~(t[205] | t[206]);
  assign t[88] = ~(t[215]);
  assign t[89] = ~(t[216]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[48]);
  assign t[92] = ~(t[133] | t[134]);
  assign t[93] = ~(t[217]);
  assign t[94] = ~(t[218]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = t[137] ? x[73] : x[72];
  assign t[97] = t[138] | t[139];
  assign t[98] = ~(t[219]);
  assign t[99] = ~(t[220]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [139:0] x;
 output y;

 wire [484:0] t;
  assign t[0] = t[1] ? t[2] : t[198];
  assign t[100] = ~(t[140] | t[141]);
  assign t[101] = t[137] ? x[81] : x[80];
  assign t[102] = ~(t[142] & t[106]);
  assign t[103] = ~(t[221]);
  assign t[104] = ~(t[210] | t[211]);
  assign t[105] = ~(t[125] | t[50]);
  assign t[106] = ~(t[143] | t[139]);
  assign t[107] = ~(t[222]);
  assign t[108] = ~(t[223]);
  assign t[109] = ~(t[144] | t[145]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[146] | t[147]);
  assign t[111] = ~(t[224] | t[148]);
  assign t[112] = t[30] ? x[95] : x[94];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[225]);
  assign t[115] = ~(t[226]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[227] | t[155]);
  assign t[119] = t[137] ? x[106] : x[105];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[156] & t[157]);
  assign t[121] = ~(t[158] & t[159]);
  assign t[122] = ~(t[160] & t[159]);
  assign t[123] = ~(x[4] & t[161]);
  assign t[124] = ~(t[162] & t[159]);
  assign t[125] = ~(t[79] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[123] & t[166]);
  assign t[128] = t[202] & t[167];
  assign t[129] = t[158] | t[160];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[199] ? t[123] : t[124];
  assign t[131] = ~(t[228]);
  assign t[132] = ~(t[215] | t[216]);
  assign t[133] = ~(t[168] & t[169]);
  assign t[134] = t[139] | t[170];
  assign t[135] = ~(t[229]);
  assign t[136] = ~(t[217] | t[218]);
  assign t[137] = ~(t[48]);
  assign t[138] = ~(t[31] & t[169]);
  assign t[139] = ~(t[164] | t[171]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[230]);
  assign t[141] = ~(t[219] | t[220]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[173]);
  assign t[144] = ~(t[231]);
  assign t[145] = ~(t[222] | t[223]);
  assign t[146] = ~(t[232]);
  assign t[147] = ~(t[233]);
  assign t[148] = ~(t[174] | t[175]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = x[4] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[225] | t[226]);
  assign t[153] = ~(t[235]);
  assign t[154] = ~(t[236]);
  assign t[155] = ~(t[179] | t[180]);
  assign t[156] = ~(t[181] | t[182]);
  assign t[157] = ~(t[183]);
  assign t[158] = ~(x[4] | t[200]);
  assign t[159] = ~(t[202]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[4] & t[200];
  assign t[161] = ~(t[200] | t[202]);
  assign t[162] = ~(x[4] | t[184]);
  assign t[163] = t[199] ? t[121] : t[122];
  assign t[164] = ~(t[79]);
  assign t[165] = t[199] ? t[124] : t[185];
  assign t[166] = ~(t[202] & t[162]);
  assign t[167] = ~(t[79] | t[199]);
  assign t[168] = ~(t[167] & t[186]);
  assign t[169] = ~(t[187] & t[188]);
  assign t[16] = ~(t[199] & t[200]);
  assign t[170] = ~(t[164] | t[189]);
  assign t[171] = t[199] ? t[166] : t[123];
  assign t[172] = ~(t[164] | t[190]);
  assign t[173] = ~(t[181] | t[177]);
  assign t[174] = ~(t[237]);
  assign t[175] = ~(t[232] | t[233]);
  assign t[176] = ~(t[164] | t[191]);
  assign t[177] = ~(t[164] | t[192]);
  assign t[178] = ~(t[31]);
  assign t[179] = ~(t[238]);
  assign t[17] = ~(t[201] & t[202]);
  assign t[180] = ~(t[235] | t[236]);
  assign t[181] = ~(t[164] | t[193]);
  assign t[182] = ~(t[194] & t[31]);
  assign t[183] = ~(t[164] | t[195]);
  assign t[184] = ~(t[200]);
  assign t[185] = ~(x[4] & t[187]);
  assign t[186] = ~(t[166] & t[185]);
  assign t[187] = ~(t[200] | t[159]);
  assign t[188] = t[164] & t[199];
  assign t[189] = t[199] ? t[196] : t[122];
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = t[199] ? t[197] : t[121];
  assign t[191] = t[199] ? t[123] : t[166];
  assign t[192] = t[199] ? t[122] : t[196];
  assign t[193] = t[199] ? t[185] : t[124];
  assign t[194] = ~(t[172] | t[51]);
  assign t[195] = t[199] ? t[121] : t[197];
  assign t[196] = ~(t[158] & t[202]);
  assign t[197] = ~(t[160] & t[202]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[7] : x[6];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = t[280] ^ x[2];
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[281] ^ x[10];
  assign t[241] = t[282] ^ x[13];
  assign t[242] = t[283] ^ x[16];
  assign t[243] = t[284] ^ x[19];
  assign t[244] = t[285] ^ x[22];
  assign t[245] = t[286] ^ x[25];
  assign t[246] = t[287] ^ x[28];
  assign t[247] = t[288] ^ x[31];
  assign t[248] = t[289] ^ x[34];
  assign t[249] = t[290] ^ x[39];
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = t[291] ^ x[42];
  assign t[251] = t[292] ^ x[45];
  assign t[252] = t[293] ^ x[48];
  assign t[253] = t[294] ^ x[53];
  assign t[254] = t[295] ^ x[56];
  assign t[255] = t[296] ^ x[59];
  assign t[256] = t[297] ^ x[62];
  assign t[257] = t[298] ^ x[65];
  assign t[258] = t[299] ^ x[68];
  assign t[259] = t[300] ^ x[71];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[260] = t[301] ^ x[76];
  assign t[261] = t[302] ^ x[79];
  assign t[262] = t[303] ^ x[84];
  assign t[263] = t[304] ^ x[87];
  assign t[264] = t[305] ^ x[90];
  assign t[265] = t[306] ^ x[93];
  assign t[266] = t[307] ^ x[98];
  assign t[267] = t[308] ^ x[101];
  assign t[268] = t[309] ^ x[104];
  assign t[269] = t[310] ^ x[109];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[311] ^ x[112];
  assign t[271] = t[312] ^ x[115];
  assign t[272] = t[313] ^ x[118];
  assign t[273] = t[314] ^ x[121];
  assign t[274] = t[315] ^ x[124];
  assign t[275] = t[316] ^ x[127];
  assign t[276] = t[317] ^ x[130];
  assign t[277] = t[318] ^ x[133];
  assign t[278] = t[319] ^ x[136];
  assign t[279] = t[320] ^ x[139];
  assign t[27] = ~(t[26] ^ t[43]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = (t[347] & ~t[348]);
  assign t[294] = (t[349] & ~t[350]);
  assign t[295] = (t[351] & ~t[352]);
  assign t[296] = (t[353] & ~t[354]);
  assign t[297] = (t[355] & ~t[356]);
  assign t[298] = (t[357] & ~t[358]);
  assign t[299] = (t[359] & ~t[360]);
  assign t[29] = x[4] ? t[47] : t[46];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (t[361] & ~t[362]);
  assign t[301] = (t[363] & ~t[364]);
  assign t[302] = (t[365] & ~t[366]);
  assign t[303] = (t[367] & ~t[368]);
  assign t[304] = (t[369] & ~t[370]);
  assign t[305] = (t[371] & ~t[372]);
  assign t[306] = (t[373] & ~t[374]);
  assign t[307] = (t[375] & ~t[376]);
  assign t[308] = (t[377] & ~t[378]);
  assign t[309] = (t[379] & ~t[380]);
  assign t[30] = ~(t[48]);
  assign t[310] = (t[381] & ~t[382]);
  assign t[311] = (t[383] & ~t[384]);
  assign t[312] = (t[385] & ~t[386]);
  assign t[313] = (t[387] & ~t[388]);
  assign t[314] = (t[389] & ~t[390]);
  assign t[315] = (t[391] & ~t[392]);
  assign t[316] = (t[393] & ~t[394]);
  assign t[317] = (t[395] & ~t[396]);
  assign t[318] = (t[397] & ~t[398]);
  assign t[319] = (t[399] & ~t[400]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (t[401] & ~t[402]);
  assign t[321] = t[403] ^ x[2];
  assign t[322] = t[404] ^ x[1];
  assign t[323] = t[405] ^ x[10];
  assign t[324] = t[406] ^ x[9];
  assign t[325] = t[407] ^ x[13];
  assign t[326] = t[408] ^ x[12];
  assign t[327] = t[409] ^ x[16];
  assign t[328] = t[410] ^ x[15];
  assign t[329] = t[411] ^ x[19];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[412] ^ x[18];
  assign t[331] = t[413] ^ x[22];
  assign t[332] = t[414] ^ x[21];
  assign t[333] = t[415] ^ x[25];
  assign t[334] = t[416] ^ x[24];
  assign t[335] = t[417] ^ x[28];
  assign t[336] = t[418] ^ x[27];
  assign t[337] = t[419] ^ x[31];
  assign t[338] = t[420] ^ x[30];
  assign t[339] = t[421] ^ x[34];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[422] ^ x[33];
  assign t[341] = t[423] ^ x[39];
  assign t[342] = t[424] ^ x[38];
  assign t[343] = t[425] ^ x[42];
  assign t[344] = t[426] ^ x[41];
  assign t[345] = t[427] ^ x[45];
  assign t[346] = t[428] ^ x[44];
  assign t[347] = t[429] ^ x[48];
  assign t[348] = t[430] ^ x[47];
  assign t[349] = t[431] ^ x[53];
  assign t[34] = ~(t[203] | t[55]);
  assign t[350] = t[432] ^ x[52];
  assign t[351] = t[433] ^ x[56];
  assign t[352] = t[434] ^ x[55];
  assign t[353] = t[435] ^ x[59];
  assign t[354] = t[436] ^ x[58];
  assign t[355] = t[437] ^ x[62];
  assign t[356] = t[438] ^ x[61];
  assign t[357] = t[439] ^ x[65];
  assign t[358] = t[440] ^ x[64];
  assign t[359] = t[441] ^ x[68];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[442] ^ x[67];
  assign t[361] = t[443] ^ x[71];
  assign t[362] = t[444] ^ x[70];
  assign t[363] = t[445] ^ x[76];
  assign t[364] = t[446] ^ x[75];
  assign t[365] = t[447] ^ x[79];
  assign t[366] = t[448] ^ x[78];
  assign t[367] = t[449] ^ x[84];
  assign t[368] = t[450] ^ x[83];
  assign t[369] = t[451] ^ x[87];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[452] ^ x[86];
  assign t[371] = t[453] ^ x[90];
  assign t[372] = t[454] ^ x[89];
  assign t[373] = t[455] ^ x[93];
  assign t[374] = t[456] ^ x[92];
  assign t[375] = t[457] ^ x[98];
  assign t[376] = t[458] ^ x[97];
  assign t[377] = t[459] ^ x[101];
  assign t[378] = t[460] ^ x[100];
  assign t[379] = t[461] ^ x[104];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[462] ^ x[103];
  assign t[381] = t[463] ^ x[109];
  assign t[382] = t[464] ^ x[108];
  assign t[383] = t[465] ^ x[112];
  assign t[384] = t[466] ^ x[111];
  assign t[385] = t[467] ^ x[115];
  assign t[386] = t[468] ^ x[114];
  assign t[387] = t[469] ^ x[118];
  assign t[388] = t[470] ^ x[117];
  assign t[389] = t[471] ^ x[121];
  assign t[38] = ~(t[39] ^ t[62]);
  assign t[390] = t[472] ^ x[120];
  assign t[391] = t[473] ^ x[124];
  assign t[392] = t[474] ^ x[123];
  assign t[393] = t[475] ^ x[127];
  assign t[394] = t[476] ^ x[126];
  assign t[395] = t[477] ^ x[130];
  assign t[396] = t[478] ^ x[129];
  assign t[397] = t[479] ^ x[133];
  assign t[398] = t[480] ^ x[132];
  assign t[399] = t[481] ^ x[136];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[482] ^ x[135];
  assign t[401] = t[483] ^ x[139];
  assign t[402] = t[484] ^ x[138];
  assign t[403] = (x[0]);
  assign t[404] = (x[0]);
  assign t[405] = (x[8]);
  assign t[406] = (x[8]);
  assign t[407] = (x[11]);
  assign t[408] = (x[11]);
  assign t[409] = (x[14]);
  assign t[40] = ~(t[44] ^ t[65]);
  assign t[410] = (x[14]);
  assign t[411] = (x[17]);
  assign t[412] = (x[17]);
  assign t[413] = (x[20]);
  assign t[414] = (x[20]);
  assign t[415] = (x[23]);
  assign t[416] = (x[23]);
  assign t[417] = (x[26]);
  assign t[418] = (x[26]);
  assign t[419] = (x[29]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[29]);
  assign t[421] = (x[32]);
  assign t[422] = (x[32]);
  assign t[423] = (x[37]);
  assign t[424] = (x[37]);
  assign t[425] = (x[40]);
  assign t[426] = (x[40]);
  assign t[427] = (x[43]);
  assign t[428] = (x[43]);
  assign t[429] = (x[46]);
  assign t[42] = ~(t[204] | t[68]);
  assign t[430] = (x[46]);
  assign t[431] = (x[51]);
  assign t[432] = (x[51]);
  assign t[433] = (x[54]);
  assign t[434] = (x[54]);
  assign t[435] = (x[57]);
  assign t[436] = (x[57]);
  assign t[437] = (x[60]);
  assign t[438] = (x[60]);
  assign t[439] = (x[63]);
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[440] = (x[63]);
  assign t[441] = (x[66]);
  assign t[442] = (x[66]);
  assign t[443] = (x[69]);
  assign t[444] = (x[69]);
  assign t[445] = (x[74]);
  assign t[446] = (x[74]);
  assign t[447] = (x[77]);
  assign t[448] = (x[77]);
  assign t[449] = (x[82]);
  assign t[44] = ~(t[71] | t[72]);
  assign t[450] = (x[82]);
  assign t[451] = (x[85]);
  assign t[452] = (x[85]);
  assign t[453] = (x[88]);
  assign t[454] = (x[88]);
  assign t[455] = (x[91]);
  assign t[456] = (x[91]);
  assign t[457] = (x[96]);
  assign t[458] = (x[96]);
  assign t[459] = (x[99]);
  assign t[45] = ~(t[73] ^ t[74]);
  assign t[460] = (x[99]);
  assign t[461] = (x[102]);
  assign t[462] = (x[102]);
  assign t[463] = (x[107]);
  assign t[464] = (x[107]);
  assign t[465] = (x[110]);
  assign t[466] = (x[110]);
  assign t[467] = (x[113]);
  assign t[468] = (x[113]);
  assign t[469] = (x[116]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (x[116]);
  assign t[471] = (x[119]);
  assign t[472] = (x[119]);
  assign t[473] = (x[122]);
  assign t[474] = (x[122]);
  assign t[475] = (x[125]);
  assign t[476] = (x[125]);
  assign t[477] = (x[128]);
  assign t[478] = (x[128]);
  assign t[479] = (x[131]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (x[131]);
  assign t[481] = (x[134]);
  assign t[482] = (x[134]);
  assign t[483] = (x[137]);
  assign t[484] = (x[137]);
  assign t[48] = ~(t[201]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = ~(t[82] & t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[205]);
  assign t[54] = ~(t[206]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[207] | t[90]);
  assign t[58] = t[91] ? x[36] : x[35];
  assign t[59] = ~(t[92] & t[84]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[93] | t[94]);
  assign t[61] = ~(t[208] | t[95]);
  assign t[62] = ~(t[96] ^ t[97]);
  assign t[63] = ~(t[98] | t[99]);
  assign t[64] = ~(t[209] | t[100]);
  assign t[65] = ~(t[101] ^ t[102]);
  assign t[66] = ~(t[210]);
  assign t[67] = ~(t[211]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = t[30] ? x[50] : x[49];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[212] | t[109]);
  assign t[73] = ~(t[110] | t[111]);
  assign t[74] = ~(t[112] ^ t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[213] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[201]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[199] ? t[122] : t[121];
  assign t[81] = t[199] ? t[124] : t[123];
  assign t[82] = ~(t[125] | t[126]);
  assign t[83] = ~(t[79] & t[127]);
  assign t[84] = ~(t[128] & t[129]);
  assign t[85] = t[79] | t[130];
  assign t[86] = ~(t[214]);
  assign t[87] = ~(t[205] | t[206]);
  assign t[88] = ~(t[215]);
  assign t[89] = ~(t[216]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[48]);
  assign t[92] = ~(t[133] | t[134]);
  assign t[93] = ~(t[217]);
  assign t[94] = ~(t[218]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = t[137] ? x[73] : x[72];
  assign t[97] = t[138] | t[139];
  assign t[98] = ~(t[219]);
  assign t[99] = ~(t[220]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[47];
  assign t[139] = t[171] ^ x[50];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[55];
  assign t[141] = t[173] ^ x[58];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[47];
  assign t[215] = t[279] ^ x[46];
  assign t[216] = t[280] ^ x[50];
  assign t[217] = t[281] ^ x[49];
  assign t[218] = t[282] ^ x[55];
  assign t[219] = t[283] ^ x[54];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[58];
  assign t[221] = t[285] ^ x[57];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[45]);
  assign t[279] = (x[45]);
  assign t[27] = t[40] ^ t[26];
  assign t[280] = (x[48]);
  assign t[281] = (x[48]);
  assign t[282] = (x[53]);
  assign t[283] = (x[53]);
  assign t[284] = (x[56]);
  assign t[285] = (x[56]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[27] : x[26];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[43];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[34];
  assign t[38] = ~(t[101] & t[56]);
  assign t[39] = ~(t[102] & t[57]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[35] : x[34];
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[106] & t[69]);
  assign t[51] = ~(t[107] & t[70]);
  assign t[52] = t[71] ? x[52] : x[51];
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = t[71] ? x[60] : x[59];
  assign t[56] = ~(t[110]);
  assign t[57] = ~(t[110] & t[74]);
  assign t[58] = ~(t[111] & t[75]);
  assign t[59] = ~(t[112] & t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[71] ? x[71] : x[70];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[79] : x[78];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[116]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116] & t[84]);
  assign t[71] = ~(t[25]);
  assign t[72] = ~(t[117]);
  assign t[73] = ~(t[117] & t[85]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[118]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[108]);
  assign t[86] = ~(t[111]);
  assign t[87] = ~(t[124]);
  assign t[88] = ~(t[124] & t[92]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [112:0] x;
 output y;

 wire [317:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[2];
  assign t[127] = t[159] ^ x[10];
  assign t[128] = t[160] ^ x[13];
  assign t[129] = t[161] ^ x[16];
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = t[162] ^ x[19];
  assign t[131] = t[163] ^ x[22];
  assign t[132] = t[164] ^ x[25];
  assign t[133] = t[165] ^ x[30];
  assign t[134] = t[166] ^ x[33];
  assign t[135] = t[167] ^ x[38];
  assign t[136] = t[168] ^ x[41];
  assign t[137] = t[169] ^ x[44];
  assign t[138] = t[170] ^ x[47];
  assign t[139] = t[171] ^ x[50];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[55];
  assign t[141] = t[173] ^ x[58];
  assign t[142] = t[174] ^ x[63];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[74];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[91];
  assign t[151] = t[183] ^ x[94];
  assign t[152] = t[184] ^ x[97];
  assign t[153] = t[185] ^ x[100];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = t[188] ^ x[109];
  assign t[157] = t[189] ^ x[112];
  assign t[158] = (t[190] & ~t[191]);
  assign t[159] = (t[192] & ~t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[194] & ~t[195]);
  assign t[161] = (t[196] & ~t[197]);
  assign t[162] = (t[198] & ~t[199]);
  assign t[163] = (t[200] & ~t[201]);
  assign t[164] = (t[202] & ~t[203]);
  assign t[165] = (t[204] & ~t[205]);
  assign t[166] = (t[206] & ~t[207]);
  assign t[167] = (t[208] & ~t[209]);
  assign t[168] = (t[210] & ~t[211]);
  assign t[169] = (t[212] & ~t[213]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (t[214] & ~t[215]);
  assign t[171] = (t[216] & ~t[217]);
  assign t[172] = (t[218] & ~t[219]);
  assign t[173] = (t[220] & ~t[221]);
  assign t[174] = (t[222] & ~t[223]);
  assign t[175] = (t[224] & ~t[225]);
  assign t[176] = (t[226] & ~t[227]);
  assign t[177] = (t[228] & ~t[229]);
  assign t[178] = (t[230] & ~t[231]);
  assign t[179] = (t[232] & ~t[233]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (t[234] & ~t[235]);
  assign t[181] = (t[236] & ~t[237]);
  assign t[182] = (t[238] & ~t[239]);
  assign t[183] = (t[240] & ~t[241]);
  assign t[184] = (t[242] & ~t[243]);
  assign t[185] = (t[244] & ~t[245]);
  assign t[186] = (t[246] & ~t[247]);
  assign t[187] = (t[248] & ~t[249]);
  assign t[188] = (t[250] & ~t[251]);
  assign t[189] = (t[252] & ~t[253]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[254] ^ x[2];
  assign t[191] = t[255] ^ x[1];
  assign t[192] = t[256] ^ x[10];
  assign t[193] = t[257] ^ x[9];
  assign t[194] = t[258] ^ x[13];
  assign t[195] = t[259] ^ x[12];
  assign t[196] = t[260] ^ x[16];
  assign t[197] = t[261] ^ x[15];
  assign t[198] = t[262] ^ x[19];
  assign t[199] = t[263] ^ x[18];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[264] ^ x[22];
  assign t[201] = t[265] ^ x[21];
  assign t[202] = t[266] ^ x[25];
  assign t[203] = t[267] ^ x[24];
  assign t[204] = t[268] ^ x[30];
  assign t[205] = t[269] ^ x[29];
  assign t[206] = t[270] ^ x[33];
  assign t[207] = t[271] ^ x[32];
  assign t[208] = t[272] ^ x[38];
  assign t[209] = t[273] ^ x[37];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[274] ^ x[41];
  assign t[211] = t[275] ^ x[40];
  assign t[212] = t[276] ^ x[44];
  assign t[213] = t[277] ^ x[43];
  assign t[214] = t[278] ^ x[47];
  assign t[215] = t[279] ^ x[46];
  assign t[216] = t[280] ^ x[50];
  assign t[217] = t[281] ^ x[49];
  assign t[218] = t[282] ^ x[55];
  assign t[219] = t[283] ^ x[54];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[284] ^ x[58];
  assign t[221] = t[285] ^ x[57];
  assign t[222] = t[286] ^ x[63];
  assign t[223] = t[287] ^ x[62];
  assign t[224] = t[288] ^ x[66];
  assign t[225] = t[289] ^ x[65];
  assign t[226] = t[290] ^ x[69];
  assign t[227] = t[291] ^ x[68];
  assign t[228] = t[292] ^ x[74];
  assign t[229] = t[293] ^ x[73];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[294] ^ x[77];
  assign t[231] = t[295] ^ x[76];
  assign t[232] = t[296] ^ x[82];
  assign t[233] = t[297] ^ x[81];
  assign t[234] = t[298] ^ x[85];
  assign t[235] = t[299] ^ x[84];
  assign t[236] = t[300] ^ x[88];
  assign t[237] = t[301] ^ x[87];
  assign t[238] = t[302] ^ x[91];
  assign t[239] = t[303] ^ x[90];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[304] ^ x[94];
  assign t[241] = t[305] ^ x[93];
  assign t[242] = t[306] ^ x[97];
  assign t[243] = t[307] ^ x[96];
  assign t[244] = t[308] ^ x[100];
  assign t[245] = t[309] ^ x[99];
  assign t[246] = t[310] ^ x[103];
  assign t[247] = t[311] ^ x[102];
  assign t[248] = t[312] ^ x[106];
  assign t[249] = t[313] ^ x[105];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[314] ^ x[109];
  assign t[251] = t[315] ^ x[108];
  assign t[252] = t[316] ^ x[112];
  assign t[253] = t[317] ^ x[111];
  assign t[254] = (x[0]);
  assign t[255] = (x[0]);
  assign t[256] = (x[8]);
  assign t[257] = (x[8]);
  assign t[258] = (x[11]);
  assign t[259] = (x[11]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[14]);
  assign t[261] = (x[14]);
  assign t[262] = (x[17]);
  assign t[263] = (x[17]);
  assign t[264] = (x[20]);
  assign t[265] = (x[20]);
  assign t[266] = (x[23]);
  assign t[267] = (x[23]);
  assign t[268] = (x[28]);
  assign t[269] = (x[28]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[31]);
  assign t[271] = (x[31]);
  assign t[272] = (x[36]);
  assign t[273] = (x[36]);
  assign t[274] = (x[39]);
  assign t[275] = (x[39]);
  assign t[276] = (x[42]);
  assign t[277] = (x[42]);
  assign t[278] = (x[45]);
  assign t[279] = (x[45]);
  assign t[27] = t[40] ^ t[26];
  assign t[280] = (x[48]);
  assign t[281] = (x[48]);
  assign t[282] = (x[53]);
  assign t[283] = (x[53]);
  assign t[284] = (x[56]);
  assign t[285] = (x[56]);
  assign t[286] = (x[61]);
  assign t[287] = (x[61]);
  assign t[288] = (x[64]);
  assign t[289] = (x[64]);
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = (x[67]);
  assign t[291] = (x[67]);
  assign t[292] = (x[72]);
  assign t[293] = (x[72]);
  assign t[294] = (x[75]);
  assign t[295] = (x[75]);
  assign t[296] = (x[80]);
  assign t[297] = (x[80]);
  assign t[298] = (x[83]);
  assign t[299] = (x[83]);
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[86]);
  assign t[301] = (x[86]);
  assign t[302] = (x[89]);
  assign t[303] = (x[89]);
  assign t[304] = (x[92]);
  assign t[305] = (x[92]);
  assign t[306] = (x[95]);
  assign t[307] = (x[95]);
  assign t[308] = (x[98]);
  assign t[309] = (x[98]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[310] = (x[101]);
  assign t[311] = (x[101]);
  assign t[312] = (x[104]);
  assign t[313] = (x[104]);
  assign t[314] = (x[107]);
  assign t[315] = (x[107]);
  assign t[316] = (x[110]);
  assign t[317] = (x[110]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[27] : x[26];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[43];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[34];
  assign t[38] = ~(t[101] & t[56]);
  assign t[39] = ~(t[102] & t[57]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[35] : x[34];
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[106] & t[69]);
  assign t[51] = ~(t[107] & t[70]);
  assign t[52] = t[71] ? x[52] : x[51];
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = t[71] ? x[60] : x[59];
  assign t[56] = ~(t[110]);
  assign t[57] = ~(t[110] & t[74]);
  assign t[58] = ~(t[111] & t[75]);
  assign t[59] = ~(t[112] & t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = t[71] ? x[71] : x[70];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[79] : x[78];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[116]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116] & t[84]);
  assign t[71] = ~(t[25]);
  assign t[72] = ~(t[117]);
  assign t[73] = ~(t[117] & t[85]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[118]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[108]);
  assign t[86] = ~(t[111]);
  assign t[87] = ~(t[124]);
  assign t[88] = ~(t[124] & t[92]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind256(x, y);
 input [139:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[108] & t[109]);
  assign t[103] = ~(t[140] & t[139]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[150]);
  assign t[107] = ~(t[110] & t[111]);
  assign t[108] = ~(t[147] & t[146]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[2];
  assign t[154] = t[195] ^ x[10];
  assign t[155] = t[196] ^ x[13];
  assign t[156] = t[197] ^ x[16];
  assign t[157] = t[198] ^ x[19];
  assign t[158] = t[199] ^ x[22];
  assign t[159] = t[200] ^ x[27];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[32];
  assign t[161] = t[202] ^ x[35];
  assign t[162] = t[203] ^ x[38];
  assign t[163] = t[204] ^ x[41];
  assign t[164] = t[205] ^ x[46];
  assign t[165] = t[206] ^ x[51];
  assign t[166] = t[207] ^ x[54];
  assign t[167] = t[208] ^ x[57];
  assign t[168] = t[209] ^ x[62];
  assign t[169] = t[210] ^ x[67];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[70];
  assign t[171] = t[212] ^ x[73];
  assign t[172] = t[213] ^ x[76];
  assign t[173] = t[214] ^ x[79];
  assign t[174] = t[215] ^ x[82];
  assign t[175] = t[216] ^ x[85];
  assign t[176] = t[217] ^ x[88];
  assign t[177] = t[218] ^ x[91];
  assign t[178] = t[219] ^ x[94];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[100];
  assign t[181] = t[222] ^ x[103];
  assign t[182] = t[223] ^ x[106];
  assign t[183] = t[224] ^ x[109];
  assign t[184] = t[225] ^ x[112];
  assign t[185] = t[226] ^ x[115];
  assign t[186] = t[227] ^ x[118];
  assign t[187] = t[228] ^ x[121];
  assign t[188] = t[229] ^ x[124];
  assign t[189] = t[230] ^ x[127];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[130];
  assign t[191] = t[232] ^ x[133];
  assign t[192] = t[233] ^ x[136];
  assign t[193] = t[234] ^ x[139];
  assign t[194] = (t[235] & ~t[236]);
  assign t[195] = (t[237] & ~t[238]);
  assign t[196] = (t[239] & ~t[240]);
  assign t[197] = (t[241] & ~t[242]);
  assign t[198] = (t[243] & ~t[244]);
  assign t[199] = (t[245] & ~t[246]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[247] & ~t[248]);
  assign t[201] = (t[249] & ~t[250]);
  assign t[202] = (t[251] & ~t[252]);
  assign t[203] = (t[253] & ~t[254]);
  assign t[204] = (t[255] & ~t[256]);
  assign t[205] = (t[257] & ~t[258]);
  assign t[206] = (t[259] & ~t[260]);
  assign t[207] = (t[261] & ~t[262]);
  assign t[208] = (t[263] & ~t[264]);
  assign t[209] = (t[265] & ~t[266]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[267] & ~t[268]);
  assign t[211] = (t[269] & ~t[270]);
  assign t[212] = (t[271] & ~t[272]);
  assign t[213] = (t[273] & ~t[274]);
  assign t[214] = (t[275] & ~t[276]);
  assign t[215] = (t[277] & ~t[278]);
  assign t[216] = (t[279] & ~t[280]);
  assign t[217] = (t[281] & ~t[282]);
  assign t[218] = (t[283] & ~t[284]);
  assign t[219] = (t[285] & ~t[286]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[287] & ~t[288]);
  assign t[221] = (t[289] & ~t[290]);
  assign t[222] = (t[291] & ~t[292]);
  assign t[223] = (t[293] & ~t[294]);
  assign t[224] = (t[295] & ~t[296]);
  assign t[225] = (t[297] & ~t[298]);
  assign t[226] = (t[299] & ~t[300]);
  assign t[227] = (t[301] & ~t[302]);
  assign t[228] = (t[303] & ~t[304]);
  assign t[229] = (t[305] & ~t[306]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[307] & ~t[308]);
  assign t[231] = (t[309] & ~t[310]);
  assign t[232] = (t[311] & ~t[312]);
  assign t[233] = (t[313] & ~t[314]);
  assign t[234] = (t[315] & ~t[316]);
  assign t[235] = t[317] ^ x[2];
  assign t[236] = t[318] ^ x[1];
  assign t[237] = t[319] ^ x[10];
  assign t[238] = t[320] ^ x[9];
  assign t[239] = t[321] ^ x[13];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[322] ^ x[12];
  assign t[241] = t[323] ^ x[16];
  assign t[242] = t[324] ^ x[15];
  assign t[243] = t[325] ^ x[19];
  assign t[244] = t[326] ^ x[18];
  assign t[245] = t[327] ^ x[22];
  assign t[246] = t[328] ^ x[21];
  assign t[247] = t[329] ^ x[27];
  assign t[248] = t[330] ^ x[26];
  assign t[249] = t[331] ^ x[32];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[332] ^ x[31];
  assign t[251] = t[333] ^ x[35];
  assign t[252] = t[334] ^ x[34];
  assign t[253] = t[335] ^ x[38];
  assign t[254] = t[336] ^ x[37];
  assign t[255] = t[337] ^ x[41];
  assign t[256] = t[338] ^ x[40];
  assign t[257] = t[339] ^ x[46];
  assign t[258] = t[340] ^ x[45];
  assign t[259] = t[341] ^ x[51];
  assign t[25] = ~(t[115]);
  assign t[260] = t[342] ^ x[50];
  assign t[261] = t[343] ^ x[54];
  assign t[262] = t[344] ^ x[53];
  assign t[263] = t[345] ^ x[57];
  assign t[264] = t[346] ^ x[56];
  assign t[265] = t[347] ^ x[62];
  assign t[266] = t[348] ^ x[61];
  assign t[267] = t[349] ^ x[67];
  assign t[268] = t[350] ^ x[66];
  assign t[269] = t[351] ^ x[70];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[352] ^ x[69];
  assign t[271] = t[353] ^ x[73];
  assign t[272] = t[354] ^ x[72];
  assign t[273] = t[355] ^ x[76];
  assign t[274] = t[356] ^ x[75];
  assign t[275] = t[357] ^ x[79];
  assign t[276] = t[358] ^ x[78];
  assign t[277] = t[359] ^ x[82];
  assign t[278] = t[360] ^ x[81];
  assign t[279] = t[361] ^ x[85];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[362] ^ x[84];
  assign t[281] = t[363] ^ x[88];
  assign t[282] = t[364] ^ x[87];
  assign t[283] = t[365] ^ x[91];
  assign t[284] = t[366] ^ x[90];
  assign t[285] = t[367] ^ x[94];
  assign t[286] = t[368] ^ x[93];
  assign t[287] = t[369] ^ x[97];
  assign t[288] = t[370] ^ x[96];
  assign t[289] = t[371] ^ x[100];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[99];
  assign t[291] = t[373] ^ x[103];
  assign t[292] = t[374] ^ x[102];
  assign t[293] = t[375] ^ x[106];
  assign t[294] = t[376] ^ x[105];
  assign t[295] = t[377] ^ x[109];
  assign t[296] = t[378] ^ x[108];
  assign t[297] = t[379] ^ x[112];
  assign t[298] = t[380] ^ x[111];
  assign t[299] = t[381] ^ x[115];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[114];
  assign t[301] = t[383] ^ x[118];
  assign t[302] = t[384] ^ x[117];
  assign t[303] = t[385] ^ x[121];
  assign t[304] = t[386] ^ x[120];
  assign t[305] = t[387] ^ x[124];
  assign t[306] = t[388] ^ x[123];
  assign t[307] = t[389] ^ x[127];
  assign t[308] = t[390] ^ x[126];
  assign t[309] = t[391] ^ x[130];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[129];
  assign t[311] = t[393] ^ x[133];
  assign t[312] = t[394] ^ x[132];
  assign t[313] = t[395] ^ x[136];
  assign t[314] = t[396] ^ x[135];
  assign t[315] = t[397] ^ x[139];
  assign t[316] = t[398] ^ x[138];
  assign t[317] = (x[0]);
  assign t[318] = (x[0]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[8]);
  assign t[321] = (x[11]);
  assign t[322] = (x[11]);
  assign t[323] = (x[14]);
  assign t[324] = (x[14]);
  assign t[325] = (x[17]);
  assign t[326] = (x[17]);
  assign t[327] = (x[20]);
  assign t[328] = (x[20]);
  assign t[329] = (x[25]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[25]);
  assign t[331] = (x[30]);
  assign t[332] = (x[30]);
  assign t[333] = (x[33]);
  assign t[334] = (x[33]);
  assign t[335] = (x[36]);
  assign t[336] = (x[36]);
  assign t[337] = (x[39]);
  assign t[338] = (x[39]);
  assign t[339] = (x[44]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[44]);
  assign t[341] = (x[49]);
  assign t[342] = (x[49]);
  assign t[343] = (x[52]);
  assign t[344] = (x[52]);
  assign t[345] = (x[55]);
  assign t[346] = (x[55]);
  assign t[347] = (x[60]);
  assign t[348] = (x[60]);
  assign t[349] = (x[65]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[65]);
  assign t[351] = (x[68]);
  assign t[352] = (x[68]);
  assign t[353] = (x[71]);
  assign t[354] = (x[71]);
  assign t[355] = (x[74]);
  assign t[356] = (x[74]);
  assign t[357] = (x[77]);
  assign t[358] = (x[77]);
  assign t[359] = (x[80]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[80]);
  assign t[361] = (x[83]);
  assign t[362] = (x[83]);
  assign t[363] = (x[86]);
  assign t[364] = (x[86]);
  assign t[365] = (x[89]);
  assign t[366] = (x[89]);
  assign t[367] = (x[92]);
  assign t[368] = (x[92]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[95]);
  assign t[371] = (x[98]);
  assign t[372] = (x[98]);
  assign t[373] = (x[101]);
  assign t[374] = (x[101]);
  assign t[375] = (x[104]);
  assign t[376] = (x[104]);
  assign t[377] = (x[107]);
  assign t[378] = (x[107]);
  assign t[379] = (x[110]);
  assign t[37] = t[56] ^ t[43];
  assign t[380] = (x[110]);
  assign t[381] = (x[113]);
  assign t[382] = (x[113]);
  assign t[383] = (x[116]);
  assign t[384] = (x[116]);
  assign t[385] = (x[119]);
  assign t[386] = (x[119]);
  assign t[387] = (x[122]);
  assign t[388] = (x[122]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[125]);
  assign t[391] = (x[128]);
  assign t[392] = (x[128]);
  assign t[393] = (x[131]);
  assign t[394] = (x[131]);
  assign t[395] = (x[134]);
  assign t[396] = (x[134]);
  assign t[397] = (x[137]);
  assign t[398] = (x[137]);
  assign t[39] = ~(t[59] & t[118]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[70] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[121]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[122]);
  assign t[53] = t[76] ? x[43] : x[42];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = ~(t[79] & t[123]);
  assign t[56] = t[76] ? x[48] : x[47];
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[125]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[126]);
  assign t[62] = t[76] ? x[59] : x[58];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = ~(t[89] & t[127]);
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = ~(t[120] & t[119]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[130]);
  assign t[72] = ~(t[92] & t[93]);
  assign t[73] = ~(t[131]);
  assign t[74] = ~(t[132]);
  assign t[75] = ~(t[94] & t[95]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[133]);
  assign t[78] = ~(t[134]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[125] & t[124]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[98] & t[99]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[140]);
  assign t[89] = ~(t[103] & t[104]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[107] & t[141]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[134] & t[133]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[137] & t[136]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [139:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[108] & t[109]);
  assign t[103] = ~(t[140] & t[139]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[150]);
  assign t[107] = ~(t[110] & t[111]);
  assign t[108] = ~(t[147] & t[146]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[2];
  assign t[154] = t[195] ^ x[10];
  assign t[155] = t[196] ^ x[13];
  assign t[156] = t[197] ^ x[16];
  assign t[157] = t[198] ^ x[19];
  assign t[158] = t[199] ^ x[22];
  assign t[159] = t[200] ^ x[27];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[32];
  assign t[161] = t[202] ^ x[35];
  assign t[162] = t[203] ^ x[38];
  assign t[163] = t[204] ^ x[41];
  assign t[164] = t[205] ^ x[46];
  assign t[165] = t[206] ^ x[51];
  assign t[166] = t[207] ^ x[54];
  assign t[167] = t[208] ^ x[57];
  assign t[168] = t[209] ^ x[62];
  assign t[169] = t[210] ^ x[67];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[70];
  assign t[171] = t[212] ^ x[73];
  assign t[172] = t[213] ^ x[76];
  assign t[173] = t[214] ^ x[79];
  assign t[174] = t[215] ^ x[82];
  assign t[175] = t[216] ^ x[85];
  assign t[176] = t[217] ^ x[88];
  assign t[177] = t[218] ^ x[91];
  assign t[178] = t[219] ^ x[94];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[100];
  assign t[181] = t[222] ^ x[103];
  assign t[182] = t[223] ^ x[106];
  assign t[183] = t[224] ^ x[109];
  assign t[184] = t[225] ^ x[112];
  assign t[185] = t[226] ^ x[115];
  assign t[186] = t[227] ^ x[118];
  assign t[187] = t[228] ^ x[121];
  assign t[188] = t[229] ^ x[124];
  assign t[189] = t[230] ^ x[127];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[130];
  assign t[191] = t[232] ^ x[133];
  assign t[192] = t[233] ^ x[136];
  assign t[193] = t[234] ^ x[139];
  assign t[194] = (t[235] & ~t[236]);
  assign t[195] = (t[237] & ~t[238]);
  assign t[196] = (t[239] & ~t[240]);
  assign t[197] = (t[241] & ~t[242]);
  assign t[198] = (t[243] & ~t[244]);
  assign t[199] = (t[245] & ~t[246]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[247] & ~t[248]);
  assign t[201] = (t[249] & ~t[250]);
  assign t[202] = (t[251] & ~t[252]);
  assign t[203] = (t[253] & ~t[254]);
  assign t[204] = (t[255] & ~t[256]);
  assign t[205] = (t[257] & ~t[258]);
  assign t[206] = (t[259] & ~t[260]);
  assign t[207] = (t[261] & ~t[262]);
  assign t[208] = (t[263] & ~t[264]);
  assign t[209] = (t[265] & ~t[266]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[267] & ~t[268]);
  assign t[211] = (t[269] & ~t[270]);
  assign t[212] = (t[271] & ~t[272]);
  assign t[213] = (t[273] & ~t[274]);
  assign t[214] = (t[275] & ~t[276]);
  assign t[215] = (t[277] & ~t[278]);
  assign t[216] = (t[279] & ~t[280]);
  assign t[217] = (t[281] & ~t[282]);
  assign t[218] = (t[283] & ~t[284]);
  assign t[219] = (t[285] & ~t[286]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[287] & ~t[288]);
  assign t[221] = (t[289] & ~t[290]);
  assign t[222] = (t[291] & ~t[292]);
  assign t[223] = (t[293] & ~t[294]);
  assign t[224] = (t[295] & ~t[296]);
  assign t[225] = (t[297] & ~t[298]);
  assign t[226] = (t[299] & ~t[300]);
  assign t[227] = (t[301] & ~t[302]);
  assign t[228] = (t[303] & ~t[304]);
  assign t[229] = (t[305] & ~t[306]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (t[307] & ~t[308]);
  assign t[231] = (t[309] & ~t[310]);
  assign t[232] = (t[311] & ~t[312]);
  assign t[233] = (t[313] & ~t[314]);
  assign t[234] = (t[315] & ~t[316]);
  assign t[235] = t[317] ^ x[2];
  assign t[236] = t[318] ^ x[1];
  assign t[237] = t[319] ^ x[10];
  assign t[238] = t[320] ^ x[9];
  assign t[239] = t[321] ^ x[13];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[322] ^ x[12];
  assign t[241] = t[323] ^ x[16];
  assign t[242] = t[324] ^ x[15];
  assign t[243] = t[325] ^ x[19];
  assign t[244] = t[326] ^ x[18];
  assign t[245] = t[327] ^ x[22];
  assign t[246] = t[328] ^ x[21];
  assign t[247] = t[329] ^ x[27];
  assign t[248] = t[330] ^ x[26];
  assign t[249] = t[331] ^ x[32];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[332] ^ x[31];
  assign t[251] = t[333] ^ x[35];
  assign t[252] = t[334] ^ x[34];
  assign t[253] = t[335] ^ x[38];
  assign t[254] = t[336] ^ x[37];
  assign t[255] = t[337] ^ x[41];
  assign t[256] = t[338] ^ x[40];
  assign t[257] = t[339] ^ x[46];
  assign t[258] = t[340] ^ x[45];
  assign t[259] = t[341] ^ x[51];
  assign t[25] = ~(t[115]);
  assign t[260] = t[342] ^ x[50];
  assign t[261] = t[343] ^ x[54];
  assign t[262] = t[344] ^ x[53];
  assign t[263] = t[345] ^ x[57];
  assign t[264] = t[346] ^ x[56];
  assign t[265] = t[347] ^ x[62];
  assign t[266] = t[348] ^ x[61];
  assign t[267] = t[349] ^ x[67];
  assign t[268] = t[350] ^ x[66];
  assign t[269] = t[351] ^ x[70];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[352] ^ x[69];
  assign t[271] = t[353] ^ x[73];
  assign t[272] = t[354] ^ x[72];
  assign t[273] = t[355] ^ x[76];
  assign t[274] = t[356] ^ x[75];
  assign t[275] = t[357] ^ x[79];
  assign t[276] = t[358] ^ x[78];
  assign t[277] = t[359] ^ x[82];
  assign t[278] = t[360] ^ x[81];
  assign t[279] = t[361] ^ x[85];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[362] ^ x[84];
  assign t[281] = t[363] ^ x[88];
  assign t[282] = t[364] ^ x[87];
  assign t[283] = t[365] ^ x[91];
  assign t[284] = t[366] ^ x[90];
  assign t[285] = t[367] ^ x[94];
  assign t[286] = t[368] ^ x[93];
  assign t[287] = t[369] ^ x[97];
  assign t[288] = t[370] ^ x[96];
  assign t[289] = t[371] ^ x[100];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[99];
  assign t[291] = t[373] ^ x[103];
  assign t[292] = t[374] ^ x[102];
  assign t[293] = t[375] ^ x[106];
  assign t[294] = t[376] ^ x[105];
  assign t[295] = t[377] ^ x[109];
  assign t[296] = t[378] ^ x[108];
  assign t[297] = t[379] ^ x[112];
  assign t[298] = t[380] ^ x[111];
  assign t[299] = t[381] ^ x[115];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[114];
  assign t[301] = t[383] ^ x[118];
  assign t[302] = t[384] ^ x[117];
  assign t[303] = t[385] ^ x[121];
  assign t[304] = t[386] ^ x[120];
  assign t[305] = t[387] ^ x[124];
  assign t[306] = t[388] ^ x[123];
  assign t[307] = t[389] ^ x[127];
  assign t[308] = t[390] ^ x[126];
  assign t[309] = t[391] ^ x[130];
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = t[392] ^ x[129];
  assign t[311] = t[393] ^ x[133];
  assign t[312] = t[394] ^ x[132];
  assign t[313] = t[395] ^ x[136];
  assign t[314] = t[396] ^ x[135];
  assign t[315] = t[397] ^ x[139];
  assign t[316] = t[398] ^ x[138];
  assign t[317] = (x[0]);
  assign t[318] = (x[0]);
  assign t[319] = (x[8]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[8]);
  assign t[321] = (x[11]);
  assign t[322] = (x[11]);
  assign t[323] = (x[14]);
  assign t[324] = (x[14]);
  assign t[325] = (x[17]);
  assign t[326] = (x[17]);
  assign t[327] = (x[20]);
  assign t[328] = (x[20]);
  assign t[329] = (x[25]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[25]);
  assign t[331] = (x[30]);
  assign t[332] = (x[30]);
  assign t[333] = (x[33]);
  assign t[334] = (x[33]);
  assign t[335] = (x[36]);
  assign t[336] = (x[36]);
  assign t[337] = (x[39]);
  assign t[338] = (x[39]);
  assign t[339] = (x[44]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[44]);
  assign t[341] = (x[49]);
  assign t[342] = (x[49]);
  assign t[343] = (x[52]);
  assign t[344] = (x[52]);
  assign t[345] = (x[55]);
  assign t[346] = (x[55]);
  assign t[347] = (x[60]);
  assign t[348] = (x[60]);
  assign t[349] = (x[65]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[65]);
  assign t[351] = (x[68]);
  assign t[352] = (x[68]);
  assign t[353] = (x[71]);
  assign t[354] = (x[71]);
  assign t[355] = (x[74]);
  assign t[356] = (x[74]);
  assign t[357] = (x[77]);
  assign t[358] = (x[77]);
  assign t[359] = (x[80]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[80]);
  assign t[361] = (x[83]);
  assign t[362] = (x[83]);
  assign t[363] = (x[86]);
  assign t[364] = (x[86]);
  assign t[365] = (x[89]);
  assign t[366] = (x[89]);
  assign t[367] = (x[92]);
  assign t[368] = (x[92]);
  assign t[369] = (x[95]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[95]);
  assign t[371] = (x[98]);
  assign t[372] = (x[98]);
  assign t[373] = (x[101]);
  assign t[374] = (x[101]);
  assign t[375] = (x[104]);
  assign t[376] = (x[104]);
  assign t[377] = (x[107]);
  assign t[378] = (x[107]);
  assign t[379] = (x[110]);
  assign t[37] = t[56] ^ t[43];
  assign t[380] = (x[110]);
  assign t[381] = (x[113]);
  assign t[382] = (x[113]);
  assign t[383] = (x[116]);
  assign t[384] = (x[116]);
  assign t[385] = (x[119]);
  assign t[386] = (x[119]);
  assign t[387] = (x[122]);
  assign t[388] = (x[122]);
  assign t[389] = (x[125]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[390] = (x[125]);
  assign t[391] = (x[128]);
  assign t[392] = (x[128]);
  assign t[393] = (x[131]);
  assign t[394] = (x[131]);
  assign t[395] = (x[134]);
  assign t[396] = (x[134]);
  assign t[397] = (x[137]);
  assign t[398] = (x[137]);
  assign t[39] = ~(t[59] & t[118]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[70] & t[71]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[121]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[122]);
  assign t[53] = t[76] ? x[43] : x[42];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = ~(t[79] & t[123]);
  assign t[56] = t[76] ? x[48] : x[47];
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[125]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[126]);
  assign t[62] = t[76] ? x[59] : x[58];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = ~(t[89] & t[127]);
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = ~(t[120] & t[119]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[130]);
  assign t[72] = ~(t[92] & t[93]);
  assign t[73] = ~(t[131]);
  assign t[74] = ~(t[132]);
  assign t[75] = ~(t[94] & t[95]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[133]);
  assign t[78] = ~(t[134]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[125] & t[124]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[98] & t[99]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[140]);
  assign t[89] = ~(t[103] & t[104]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[107] & t[141]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[134] & t[133]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[137] & t[136]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [139:0] x;
 output y;

 wire [389:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[102] | t[98]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[2];
  assign t[145] = t[186] ^ x[10];
  assign t[146] = t[187] ^ x[13];
  assign t[147] = t[188] ^ x[16];
  assign t[148] = t[189] ^ x[19];
  assign t[149] = t[190] ^ x[22];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[27];
  assign t[151] = t[192] ^ x[32];
  assign t[152] = t[193] ^ x[35];
  assign t[153] = t[194] ^ x[38];
  assign t[154] = t[195] ^ x[41];
  assign t[155] = t[196] ^ x[46];
  assign t[156] = t[197] ^ x[51];
  assign t[157] = t[198] ^ x[54];
  assign t[158] = t[199] ^ x[57];
  assign t[159] = t[200] ^ x[62];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[67];
  assign t[161] = t[202] ^ x[70];
  assign t[162] = t[203] ^ x[73];
  assign t[163] = t[204] ^ x[76];
  assign t[164] = t[205] ^ x[79];
  assign t[165] = t[206] ^ x[82];
  assign t[166] = t[207] ^ x[85];
  assign t[167] = t[208] ^ x[88];
  assign t[168] = t[209] ^ x[91];
  assign t[169] = t[210] ^ x[94];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[100];
  assign t[172] = t[213] ^ x[103];
  assign t[173] = t[214] ^ x[106];
  assign t[174] = t[215] ^ x[109];
  assign t[175] = t[216] ^ x[112];
  assign t[176] = t[217] ^ x[115];
  assign t[177] = t[218] ^ x[118];
  assign t[178] = t[219] ^ x[121];
  assign t[179] = t[220] ^ x[124];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[127];
  assign t[181] = t[222] ^ x[130];
  assign t[182] = t[223] ^ x[133];
  assign t[183] = t[224] ^ x[136];
  assign t[184] = t[225] ^ x[139];
  assign t[185] = (t[226] & ~t[227]);
  assign t[186] = (t[228] & ~t[229]);
  assign t[187] = (t[230] & ~t[231]);
  assign t[188] = (t[232] & ~t[233]);
  assign t[189] = (t[234] & ~t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[236] & ~t[237]);
  assign t[191] = (t[238] & ~t[239]);
  assign t[192] = (t[240] & ~t[241]);
  assign t[193] = (t[242] & ~t[243]);
  assign t[194] = (t[244] & ~t[245]);
  assign t[195] = (t[246] & ~t[247]);
  assign t[196] = (t[248] & ~t[249]);
  assign t[197] = (t[250] & ~t[251]);
  assign t[198] = (t[252] & ~t[253]);
  assign t[199] = (t[254] & ~t[255]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[256] & ~t[257]);
  assign t[201] = (t[258] & ~t[259]);
  assign t[202] = (t[260] & ~t[261]);
  assign t[203] = (t[262] & ~t[263]);
  assign t[204] = (t[264] & ~t[265]);
  assign t[205] = (t[266] & ~t[267]);
  assign t[206] = (t[268] & ~t[269]);
  assign t[207] = (t[270] & ~t[271]);
  assign t[208] = (t[272] & ~t[273]);
  assign t[209] = (t[274] & ~t[275]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[276] & ~t[277]);
  assign t[211] = (t[278] & ~t[279]);
  assign t[212] = (t[280] & ~t[281]);
  assign t[213] = (t[282] & ~t[283]);
  assign t[214] = (t[284] & ~t[285]);
  assign t[215] = (t[286] & ~t[287]);
  assign t[216] = (t[288] & ~t[289]);
  assign t[217] = (t[290] & ~t[291]);
  assign t[218] = (t[292] & ~t[293]);
  assign t[219] = (t[294] & ~t[295]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[296] & ~t[297]);
  assign t[221] = (t[298] & ~t[299]);
  assign t[222] = (t[300] & ~t[301]);
  assign t[223] = (t[302] & ~t[303]);
  assign t[224] = (t[304] & ~t[305]);
  assign t[225] = (t[306] & ~t[307]);
  assign t[226] = t[308] ^ x[2];
  assign t[227] = t[309] ^ x[1];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[9];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[12];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[15];
  assign t[234] = t[316] ^ x[19];
  assign t[235] = t[317] ^ x[18];
  assign t[236] = t[318] ^ x[22];
  assign t[237] = t[319] ^ x[21];
  assign t[238] = t[320] ^ x[27];
  assign t[239] = t[321] ^ x[26];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[322] ^ x[32];
  assign t[241] = t[323] ^ x[31];
  assign t[242] = t[324] ^ x[35];
  assign t[243] = t[325] ^ x[34];
  assign t[244] = t[326] ^ x[38];
  assign t[245] = t[327] ^ x[37];
  assign t[246] = t[328] ^ x[41];
  assign t[247] = t[329] ^ x[40];
  assign t[248] = t[330] ^ x[46];
  assign t[249] = t[331] ^ x[45];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[332] ^ x[51];
  assign t[251] = t[333] ^ x[50];
  assign t[252] = t[334] ^ x[54];
  assign t[253] = t[335] ^ x[53];
  assign t[254] = t[336] ^ x[57];
  assign t[255] = t[337] ^ x[56];
  assign t[256] = t[338] ^ x[62];
  assign t[257] = t[339] ^ x[61];
  assign t[258] = t[340] ^ x[67];
  assign t[259] = t[341] ^ x[66];
  assign t[25] = ~(t[106]);
  assign t[260] = t[342] ^ x[70];
  assign t[261] = t[343] ^ x[69];
  assign t[262] = t[344] ^ x[73];
  assign t[263] = t[345] ^ x[72];
  assign t[264] = t[346] ^ x[76];
  assign t[265] = t[347] ^ x[75];
  assign t[266] = t[348] ^ x[79];
  assign t[267] = t[349] ^ x[78];
  assign t[268] = t[350] ^ x[82];
  assign t[269] = t[351] ^ x[81];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[352] ^ x[85];
  assign t[271] = t[353] ^ x[84];
  assign t[272] = t[354] ^ x[88];
  assign t[273] = t[355] ^ x[87];
  assign t[274] = t[356] ^ x[91];
  assign t[275] = t[357] ^ x[90];
  assign t[276] = t[358] ^ x[94];
  assign t[277] = t[359] ^ x[93];
  assign t[278] = t[360] ^ x[97];
  assign t[279] = t[361] ^ x[96];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[362] ^ x[100];
  assign t[281] = t[363] ^ x[99];
  assign t[282] = t[364] ^ x[103];
  assign t[283] = t[365] ^ x[102];
  assign t[284] = t[366] ^ x[106];
  assign t[285] = t[367] ^ x[105];
  assign t[286] = t[368] ^ x[109];
  assign t[287] = t[369] ^ x[108];
  assign t[288] = t[370] ^ x[112];
  assign t[289] = t[371] ^ x[111];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[115];
  assign t[291] = t[373] ^ x[114];
  assign t[292] = t[374] ^ x[118];
  assign t[293] = t[375] ^ x[117];
  assign t[294] = t[376] ^ x[121];
  assign t[295] = t[377] ^ x[120];
  assign t[296] = t[378] ^ x[124];
  assign t[297] = t[379] ^ x[123];
  assign t[298] = t[380] ^ x[127];
  assign t[299] = t[381] ^ x[126];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[130];
  assign t[301] = t[383] ^ x[129];
  assign t[302] = t[384] ^ x[133];
  assign t[303] = t[385] ^ x[132];
  assign t[304] = t[386] ^ x[136];
  assign t[305] = t[387] ^ x[135];
  assign t[306] = t[388] ^ x[139];
  assign t[307] = t[389] ^ x[138];
  assign t[308] = (x[0]);
  assign t[309] = (x[0]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[8]);
  assign t[312] = (x[11]);
  assign t[313] = (x[11]);
  assign t[314] = (x[14]);
  assign t[315] = (x[14]);
  assign t[316] = (x[17]);
  assign t[317] = (x[17]);
  assign t[318] = (x[20]);
  assign t[319] = (x[20]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[25]);
  assign t[321] = (x[25]);
  assign t[322] = (x[30]);
  assign t[323] = (x[30]);
  assign t[324] = (x[33]);
  assign t[325] = (x[33]);
  assign t[326] = (x[36]);
  assign t[327] = (x[36]);
  assign t[328] = (x[39]);
  assign t[329] = (x[39]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[44]);
  assign t[331] = (x[44]);
  assign t[332] = (x[49]);
  assign t[333] = (x[49]);
  assign t[334] = (x[52]);
  assign t[335] = (x[52]);
  assign t[336] = (x[55]);
  assign t[337] = (x[55]);
  assign t[338] = (x[60]);
  assign t[339] = (x[60]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[65]);
  assign t[341] = (x[65]);
  assign t[342] = (x[68]);
  assign t[343] = (x[68]);
  assign t[344] = (x[71]);
  assign t[345] = (x[71]);
  assign t[346] = (x[74]);
  assign t[347] = (x[74]);
  assign t[348] = (x[77]);
  assign t[349] = (x[77]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[80]);
  assign t[351] = (x[80]);
  assign t[352] = (x[83]);
  assign t[353] = (x[83]);
  assign t[354] = (x[86]);
  assign t[355] = (x[86]);
  assign t[356] = (x[89]);
  assign t[357] = (x[89]);
  assign t[358] = (x[92]);
  assign t[359] = (x[92]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[95]);
  assign t[361] = (x[95]);
  assign t[362] = (x[98]);
  assign t[363] = (x[98]);
  assign t[364] = (x[101]);
  assign t[365] = (x[101]);
  assign t[366] = (x[104]);
  assign t[367] = (x[104]);
  assign t[368] = (x[107]);
  assign t[369] = (x[107]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[110]);
  assign t[371] = (x[110]);
  assign t[372] = (x[113]);
  assign t[373] = (x[113]);
  assign t[374] = (x[116]);
  assign t[375] = (x[116]);
  assign t[376] = (x[119]);
  assign t[377] = (x[119]);
  assign t[378] = (x[122]);
  assign t[379] = (x[122]);
  assign t[37] = t[56] ^ t[43];
  assign t[380] = (x[125]);
  assign t[381] = (x[125]);
  assign t[382] = (x[128]);
  assign t[383] = (x[128]);
  assign t[384] = (x[131]);
  assign t[385] = (x[131]);
  assign t[386] = (x[134]);
  assign t[387] = (x[134]);
  assign t[388] = (x[137]);
  assign t[389] = (x[137]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] | t[109];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[69] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[71] | t[112];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = t[74] | t[113];
  assign t[53] = t[75] ? x[43] : x[42];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = t[78] | t[114];
  assign t[56] = t[75] ? x[48] : x[47];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[79] | t[57]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[80] & t[81]);
  assign t[61] = t[82] | t[117];
  assign t[62] = t[75] ? x[59] : x[58];
  assign t[63] = ~(t[83] & t[84]);
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = t[87] | t[118];
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[88] & t[89]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[91] | t[72]);
  assign t[75] = ~(t[25]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[93] | t[80]);
  assign t[83] = ~(t[94] & t[95]);
  assign t[84] = t[96] | t[129];
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[131]);
  assign t[87] = ~(t[97] | t[85]);
  assign t[88] = ~(t[98] & t[99]);
  assign t[89] = t[100] | t[132];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[137]);
  assign t[95] = ~(t[138]);
  assign t[96] = ~(t[101] | t[94]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [139:0] x;
 output y;

 wire [389:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[102] | t[98]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[7] : x[6];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[2];
  assign t[145] = t[186] ^ x[10];
  assign t[146] = t[187] ^ x[13];
  assign t[147] = t[188] ^ x[16];
  assign t[148] = t[189] ^ x[19];
  assign t[149] = t[190] ^ x[22];
  assign t[14] = x[4] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[27];
  assign t[151] = t[192] ^ x[32];
  assign t[152] = t[193] ^ x[35];
  assign t[153] = t[194] ^ x[38];
  assign t[154] = t[195] ^ x[41];
  assign t[155] = t[196] ^ x[46];
  assign t[156] = t[197] ^ x[51];
  assign t[157] = t[198] ^ x[54];
  assign t[158] = t[199] ^ x[57];
  assign t[159] = t[200] ^ x[62];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[67];
  assign t[161] = t[202] ^ x[70];
  assign t[162] = t[203] ^ x[73];
  assign t[163] = t[204] ^ x[76];
  assign t[164] = t[205] ^ x[79];
  assign t[165] = t[206] ^ x[82];
  assign t[166] = t[207] ^ x[85];
  assign t[167] = t[208] ^ x[88];
  assign t[168] = t[209] ^ x[91];
  assign t[169] = t[210] ^ x[94];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[100];
  assign t[172] = t[213] ^ x[103];
  assign t[173] = t[214] ^ x[106];
  assign t[174] = t[215] ^ x[109];
  assign t[175] = t[216] ^ x[112];
  assign t[176] = t[217] ^ x[115];
  assign t[177] = t[218] ^ x[118];
  assign t[178] = t[219] ^ x[121];
  assign t[179] = t[220] ^ x[124];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[127];
  assign t[181] = t[222] ^ x[130];
  assign t[182] = t[223] ^ x[133];
  assign t[183] = t[224] ^ x[136];
  assign t[184] = t[225] ^ x[139];
  assign t[185] = (t[226] & ~t[227]);
  assign t[186] = (t[228] & ~t[229]);
  assign t[187] = (t[230] & ~t[231]);
  assign t[188] = (t[232] & ~t[233]);
  assign t[189] = (t[234] & ~t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[236] & ~t[237]);
  assign t[191] = (t[238] & ~t[239]);
  assign t[192] = (t[240] & ~t[241]);
  assign t[193] = (t[242] & ~t[243]);
  assign t[194] = (t[244] & ~t[245]);
  assign t[195] = (t[246] & ~t[247]);
  assign t[196] = (t[248] & ~t[249]);
  assign t[197] = (t[250] & ~t[251]);
  assign t[198] = (t[252] & ~t[253]);
  assign t[199] = (t[254] & ~t[255]);
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (t[256] & ~t[257]);
  assign t[201] = (t[258] & ~t[259]);
  assign t[202] = (t[260] & ~t[261]);
  assign t[203] = (t[262] & ~t[263]);
  assign t[204] = (t[264] & ~t[265]);
  assign t[205] = (t[266] & ~t[267]);
  assign t[206] = (t[268] & ~t[269]);
  assign t[207] = (t[270] & ~t[271]);
  assign t[208] = (t[272] & ~t[273]);
  assign t[209] = (t[274] & ~t[275]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[276] & ~t[277]);
  assign t[211] = (t[278] & ~t[279]);
  assign t[212] = (t[280] & ~t[281]);
  assign t[213] = (t[282] & ~t[283]);
  assign t[214] = (t[284] & ~t[285]);
  assign t[215] = (t[286] & ~t[287]);
  assign t[216] = (t[288] & ~t[289]);
  assign t[217] = (t[290] & ~t[291]);
  assign t[218] = (t[292] & ~t[293]);
  assign t[219] = (t[294] & ~t[295]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[296] & ~t[297]);
  assign t[221] = (t[298] & ~t[299]);
  assign t[222] = (t[300] & ~t[301]);
  assign t[223] = (t[302] & ~t[303]);
  assign t[224] = (t[304] & ~t[305]);
  assign t[225] = (t[306] & ~t[307]);
  assign t[226] = t[308] ^ x[2];
  assign t[227] = t[309] ^ x[1];
  assign t[228] = t[310] ^ x[10];
  assign t[229] = t[311] ^ x[9];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[312] ^ x[13];
  assign t[231] = t[313] ^ x[12];
  assign t[232] = t[314] ^ x[16];
  assign t[233] = t[315] ^ x[15];
  assign t[234] = t[316] ^ x[19];
  assign t[235] = t[317] ^ x[18];
  assign t[236] = t[318] ^ x[22];
  assign t[237] = t[319] ^ x[21];
  assign t[238] = t[320] ^ x[27];
  assign t[239] = t[321] ^ x[26];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[322] ^ x[32];
  assign t[241] = t[323] ^ x[31];
  assign t[242] = t[324] ^ x[35];
  assign t[243] = t[325] ^ x[34];
  assign t[244] = t[326] ^ x[38];
  assign t[245] = t[327] ^ x[37];
  assign t[246] = t[328] ^ x[41];
  assign t[247] = t[329] ^ x[40];
  assign t[248] = t[330] ^ x[46];
  assign t[249] = t[331] ^ x[45];
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = t[332] ^ x[51];
  assign t[251] = t[333] ^ x[50];
  assign t[252] = t[334] ^ x[54];
  assign t[253] = t[335] ^ x[53];
  assign t[254] = t[336] ^ x[57];
  assign t[255] = t[337] ^ x[56];
  assign t[256] = t[338] ^ x[62];
  assign t[257] = t[339] ^ x[61];
  assign t[258] = t[340] ^ x[67];
  assign t[259] = t[341] ^ x[66];
  assign t[25] = ~(t[106]);
  assign t[260] = t[342] ^ x[70];
  assign t[261] = t[343] ^ x[69];
  assign t[262] = t[344] ^ x[73];
  assign t[263] = t[345] ^ x[72];
  assign t[264] = t[346] ^ x[76];
  assign t[265] = t[347] ^ x[75];
  assign t[266] = t[348] ^ x[79];
  assign t[267] = t[349] ^ x[78];
  assign t[268] = t[350] ^ x[82];
  assign t[269] = t[351] ^ x[81];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[352] ^ x[85];
  assign t[271] = t[353] ^ x[84];
  assign t[272] = t[354] ^ x[88];
  assign t[273] = t[355] ^ x[87];
  assign t[274] = t[356] ^ x[91];
  assign t[275] = t[357] ^ x[90];
  assign t[276] = t[358] ^ x[94];
  assign t[277] = t[359] ^ x[93];
  assign t[278] = t[360] ^ x[97];
  assign t[279] = t[361] ^ x[96];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[362] ^ x[100];
  assign t[281] = t[363] ^ x[99];
  assign t[282] = t[364] ^ x[103];
  assign t[283] = t[365] ^ x[102];
  assign t[284] = t[366] ^ x[106];
  assign t[285] = t[367] ^ x[105];
  assign t[286] = t[368] ^ x[109];
  assign t[287] = t[369] ^ x[108];
  assign t[288] = t[370] ^ x[112];
  assign t[289] = t[371] ^ x[111];
  assign t[28] = x[4] ? t[42] : t[41];
  assign t[290] = t[372] ^ x[115];
  assign t[291] = t[373] ^ x[114];
  assign t[292] = t[374] ^ x[118];
  assign t[293] = t[375] ^ x[117];
  assign t[294] = t[376] ^ x[121];
  assign t[295] = t[377] ^ x[120];
  assign t[296] = t[378] ^ x[124];
  assign t[297] = t[379] ^ x[123];
  assign t[298] = t[380] ^ x[127];
  assign t[299] = t[381] ^ x[126];
  assign t[29] = x[4] ? t[44] : t[43];
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = t[382] ^ x[130];
  assign t[301] = t[383] ^ x[129];
  assign t[302] = t[384] ^ x[133];
  assign t[303] = t[385] ^ x[132];
  assign t[304] = t[386] ^ x[136];
  assign t[305] = t[387] ^ x[135];
  assign t[306] = t[388] ^ x[139];
  assign t[307] = t[389] ^ x[138];
  assign t[308] = (x[0]);
  assign t[309] = (x[0]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[8]);
  assign t[311] = (x[8]);
  assign t[312] = (x[11]);
  assign t[313] = (x[11]);
  assign t[314] = (x[14]);
  assign t[315] = (x[14]);
  assign t[316] = (x[17]);
  assign t[317] = (x[17]);
  assign t[318] = (x[20]);
  assign t[319] = (x[20]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[25]);
  assign t[321] = (x[25]);
  assign t[322] = (x[30]);
  assign t[323] = (x[30]);
  assign t[324] = (x[33]);
  assign t[325] = (x[33]);
  assign t[326] = (x[36]);
  assign t[327] = (x[36]);
  assign t[328] = (x[39]);
  assign t[329] = (x[39]);
  assign t[32] = t[48] ? x[24] : x[23];
  assign t[330] = (x[44]);
  assign t[331] = (x[44]);
  assign t[332] = (x[49]);
  assign t[333] = (x[49]);
  assign t[334] = (x[52]);
  assign t[335] = (x[52]);
  assign t[336] = (x[55]);
  assign t[337] = (x[55]);
  assign t[338] = (x[60]);
  assign t[339] = (x[60]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[65]);
  assign t[341] = (x[65]);
  assign t[342] = (x[68]);
  assign t[343] = (x[68]);
  assign t[344] = (x[71]);
  assign t[345] = (x[71]);
  assign t[346] = (x[74]);
  assign t[347] = (x[74]);
  assign t[348] = (x[77]);
  assign t[349] = (x[77]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[80]);
  assign t[351] = (x[80]);
  assign t[352] = (x[83]);
  assign t[353] = (x[83]);
  assign t[354] = (x[86]);
  assign t[355] = (x[86]);
  assign t[356] = (x[89]);
  assign t[357] = (x[89]);
  assign t[358] = (x[92]);
  assign t[359] = (x[92]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[95]);
  assign t[361] = (x[95]);
  assign t[362] = (x[98]);
  assign t[363] = (x[98]);
  assign t[364] = (x[101]);
  assign t[365] = (x[101]);
  assign t[366] = (x[104]);
  assign t[367] = (x[104]);
  assign t[368] = (x[107]);
  assign t[369] = (x[107]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[110]);
  assign t[371] = (x[110]);
  assign t[372] = (x[113]);
  assign t[373] = (x[113]);
  assign t[374] = (x[116]);
  assign t[375] = (x[116]);
  assign t[376] = (x[119]);
  assign t[377] = (x[119]);
  assign t[378] = (x[122]);
  assign t[379] = (x[122]);
  assign t[37] = t[56] ^ t[43];
  assign t[380] = (x[125]);
  assign t[381] = (x[125]);
  assign t[382] = (x[128]);
  assign t[383] = (x[128]);
  assign t[384] = (x[131]);
  assign t[385] = (x[131]);
  assign t[386] = (x[134]);
  assign t[387] = (x[134]);
  assign t[388] = (x[137]);
  assign t[389] = (x[137]);
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] | t[109];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[29] : x[28];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[69] & t[70]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = t[71] | t[112];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = t[74] | t[113];
  assign t[53] = t[75] ? x[43] : x[42];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = t[78] | t[114];
  assign t[56] = t[75] ? x[48] : x[47];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[79] | t[57]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[80] & t[81]);
  assign t[61] = t[82] | t[117];
  assign t[62] = t[75] ? x[59] : x[58];
  assign t[63] = ~(t[83] & t[84]);
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = t[87] | t[118];
  assign t[66] = t[18] ? x[64] : x[63];
  assign t[67] = ~(t[88] & t[89]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[91] | t[72]);
  assign t[75] = ~(t[25]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[93] | t[80]);
  assign t[83] = ~(t[94] & t[95]);
  assign t[84] = t[96] | t[129];
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[131]);
  assign t[87] = ~(t[97] | t[85]);
  assign t[88] = ~(t[98] & t[99]);
  assign t[89] = t[100] | t[132];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[137]);
  assign t[95] = ~(t[138]);
  assign t[96] = ~(t[101] | t[94]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[141]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [97:0] x;
 output y;

 wire [347:0] t;
  assign t[0] = t[1] ? t[2] : t[145];
  assign t[100] = ~(t[169]);
  assign t[101] = ~(t[162] | t[163]);
  assign t[102] = ~(t[170]);
  assign t[103] = ~(t[171]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[34]);
  assign t[106] = ~(t[85] | t[127]);
  assign t[107] = ~(t[128]);
  assign t[108] = x[4] & t[147];
  assign t[109] = ~(t[149]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = ~(x[4] | t[147]);
  assign t[111] = ~(t[147] | t[149]);
  assign t[112] = ~(x[4] | t[129]);
  assign t[113] = t[146] ? t[130] : t[84];
  assign t[114] = t[146] ? t[81] : t[131];
  assign t[115] = t[146] ? t[81] : t[82];
  assign t[116] = ~(t[35] | t[132]);
  assign t[117] = ~(t[54] & t[133]);
  assign t[118] = ~(t[123] & t[134]);
  assign t[119] = t[54] | t[135];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[172]);
  assign t[121] = ~(t[167] | t[168]);
  assign t[122] = ~(t[58] | t[136]);
  assign t[123] = t[149] & t[137];
  assign t[124] = ~(t[65]);
  assign t[125] = ~(t[173]);
  assign t[126] = ~(t[170] | t[171]);
  assign t[127] = ~(t[138] & t[65]);
  assign t[128] = ~(t[58] | t[139]);
  assign t[129] = ~(t[147]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(x[4] & t[140]);
  assign t[131] = ~(t[110] & t[149]);
  assign t[132] = ~(t[58] | t[141]);
  assign t[133] = ~(t[83] & t[87]);
  assign t[134] = t[110] | t[108];
  assign t[135] = t[146] ? t[83] : t[84];
  assign t[136] = t[146] ? t[83] : t[87];
  assign t[137] = ~(t[54] | t[146]);
  assign t[138] = ~(t[142] | t[91]);
  assign t[139] = t[146] ? t[82] : t[143];
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = ~(t[147] | t[109]);
  assign t[141] = t[146] ? t[84] : t[130];
  assign t[142] = ~(t[58] | t[144]);
  assign t[143] = ~(t[108] & t[149]);
  assign t[144] = t[146] ? t[143] : t[82];
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = ~(t[146] & t[147]);
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = (t[195]);
  assign t[167] = (t[196]);
  assign t[168] = (t[197]);
  assign t[169] = (t[198]);
  assign t[16] = ~(t[148] & t[149]);
  assign t[170] = (t[199]);
  assign t[171] = (t[200]);
  assign t[172] = (t[201]);
  assign t[173] = (t[202]);
  assign t[174] = t[203] ^ x[2];
  assign t[175] = t[204] ^ x[10];
  assign t[176] = t[205] ^ x[13];
  assign t[177] = t[206] ^ x[16];
  assign t[178] = t[207] ^ x[19];
  assign t[179] = t[208] ^ x[22];
  assign t[17] = t[23] ? x[7] : x[6];
  assign t[180] = t[209] ^ x[25];
  assign t[181] = t[210] ^ x[28];
  assign t[182] = t[211] ^ x[31];
  assign t[183] = t[212] ^ x[36];
  assign t[184] = t[213] ^ x[39];
  assign t[185] = t[214] ^ x[42];
  assign t[186] = t[215] ^ x[45];
  assign t[187] = t[216] ^ x[48];
  assign t[188] = t[217] ^ x[51];
  assign t[189] = t[218] ^ x[54];
  assign t[18] = ~(t[24] & t[25]);
  assign t[190] = t[219] ^ x[57];
  assign t[191] = t[220] ^ x[62];
  assign t[192] = t[221] ^ x[65];
  assign t[193] = t[222] ^ x[68];
  assign t[194] = t[223] ^ x[73];
  assign t[195] = t[224] ^ x[76];
  assign t[196] = t[225] ^ x[79];
  assign t[197] = t[226] ^ x[82];
  assign t[198] = t[227] ^ x[85];
  assign t[199] = t[228] ^ x[88];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[229] ^ x[91];
  assign t[201] = t[230] ^ x[94];
  assign t[202] = t[231] ^ x[97];
  assign t[203] = (t[232] & ~t[233]);
  assign t[204] = (t[234] & ~t[235]);
  assign t[205] = (t[236] & ~t[237]);
  assign t[206] = (t[238] & ~t[239]);
  assign t[207] = (t[240] & ~t[241]);
  assign t[208] = (t[242] & ~t[243]);
  assign t[209] = (t[244] & ~t[245]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[246] & ~t[247]);
  assign t[211] = (t[248] & ~t[249]);
  assign t[212] = (t[250] & ~t[251]);
  assign t[213] = (t[252] & ~t[253]);
  assign t[214] = (t[254] & ~t[255]);
  assign t[215] = (t[256] & ~t[257]);
  assign t[216] = (t[258] & ~t[259]);
  assign t[217] = (t[260] & ~t[261]);
  assign t[218] = (t[262] & ~t[263]);
  assign t[219] = (t[264] & ~t[265]);
  assign t[21] = x[4] ? t[31] : t[30];
  assign t[220] = (t[266] & ~t[267]);
  assign t[221] = (t[268] & ~t[269]);
  assign t[222] = (t[270] & ~t[271]);
  assign t[223] = (t[272] & ~t[273]);
  assign t[224] = (t[274] & ~t[275]);
  assign t[225] = (t[276] & ~t[277]);
  assign t[226] = (t[278] & ~t[279]);
  assign t[227] = (t[280] & ~t[281]);
  assign t[228] = (t[282] & ~t[283]);
  assign t[229] = (t[284] & ~t[285]);
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[230] = (t[286] & ~t[287]);
  assign t[231] = (t[288] & ~t[289]);
  assign t[232] = t[290] ^ x[2];
  assign t[233] = t[291] ^ x[1];
  assign t[234] = t[292] ^ x[10];
  assign t[235] = t[293] ^ x[9];
  assign t[236] = t[294] ^ x[13];
  assign t[237] = t[295] ^ x[12];
  assign t[238] = t[296] ^ x[16];
  assign t[239] = t[297] ^ x[15];
  assign t[23] = ~(t[34]);
  assign t[240] = t[298] ^ x[19];
  assign t[241] = t[299] ^ x[18];
  assign t[242] = t[300] ^ x[22];
  assign t[243] = t[301] ^ x[21];
  assign t[244] = t[302] ^ x[25];
  assign t[245] = t[303] ^ x[24];
  assign t[246] = t[304] ^ x[28];
  assign t[247] = t[305] ^ x[27];
  assign t[248] = t[306] ^ x[31];
  assign t[249] = t[307] ^ x[30];
  assign t[24] = ~(t[35] | t[36]);
  assign t[250] = t[308] ^ x[36];
  assign t[251] = t[309] ^ x[35];
  assign t[252] = t[310] ^ x[39];
  assign t[253] = t[311] ^ x[38];
  assign t[254] = t[312] ^ x[42];
  assign t[255] = t[313] ^ x[41];
  assign t[256] = t[314] ^ x[45];
  assign t[257] = t[315] ^ x[44];
  assign t[258] = t[316] ^ x[48];
  assign t[259] = t[317] ^ x[47];
  assign t[25] = ~(t[37] | t[38]);
  assign t[260] = t[318] ^ x[51];
  assign t[261] = t[319] ^ x[50];
  assign t[262] = t[320] ^ x[54];
  assign t[263] = t[321] ^ x[53];
  assign t[264] = t[322] ^ x[57];
  assign t[265] = t[323] ^ x[56];
  assign t[266] = t[324] ^ x[62];
  assign t[267] = t[325] ^ x[61];
  assign t[268] = t[326] ^ x[65];
  assign t[269] = t[327] ^ x[64];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[328] ^ x[68];
  assign t[271] = t[329] ^ x[67];
  assign t[272] = t[330] ^ x[73];
  assign t[273] = t[331] ^ x[72];
  assign t[274] = t[332] ^ x[76];
  assign t[275] = t[333] ^ x[75];
  assign t[276] = t[334] ^ x[79];
  assign t[277] = t[335] ^ x[78];
  assign t[278] = t[336] ^ x[82];
  assign t[279] = t[337] ^ x[81];
  assign t[27] = ~(t[150] | t[41]);
  assign t[280] = t[338] ^ x[85];
  assign t[281] = t[339] ^ x[84];
  assign t[282] = t[340] ^ x[88];
  assign t[283] = t[341] ^ x[87];
  assign t[284] = t[342] ^ x[91];
  assign t[285] = t[343] ^ x[90];
  assign t[286] = t[344] ^ x[94];
  assign t[287] = t[345] ^ x[93];
  assign t[288] = t[346] ^ x[97];
  assign t[289] = t[347] ^ x[96];
  assign t[28] = ~(t[42] | t[43]);
  assign t[290] = (x[0]);
  assign t[291] = (x[0]);
  assign t[292] = (x[8]);
  assign t[293] = (x[8]);
  assign t[294] = (x[11]);
  assign t[295] = (x[11]);
  assign t[296] = (x[14]);
  assign t[297] = (x[14]);
  assign t[298] = (x[17]);
  assign t[299] = (x[17]);
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[20]);
  assign t[301] = (x[20]);
  assign t[302] = (x[23]);
  assign t[303] = (x[23]);
  assign t[304] = (x[26]);
  assign t[305] = (x[26]);
  assign t[306] = (x[29]);
  assign t[307] = (x[29]);
  assign t[308] = (x[34]);
  assign t[309] = (x[34]);
  assign t[30] = ~(t[46] | t[47]);
  assign t[310] = (x[37]);
  assign t[311] = (x[37]);
  assign t[312] = (x[40]);
  assign t[313] = (x[40]);
  assign t[314] = (x[43]);
  assign t[315] = (x[43]);
  assign t[316] = (x[46]);
  assign t[317] = (x[46]);
  assign t[318] = (x[49]);
  assign t[319] = (x[49]);
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[320] = (x[52]);
  assign t[321] = (x[52]);
  assign t[322] = (x[55]);
  assign t[323] = (x[55]);
  assign t[324] = (x[60]);
  assign t[325] = (x[60]);
  assign t[326] = (x[63]);
  assign t[327] = (x[63]);
  assign t[328] = (x[66]);
  assign t[329] = (x[66]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[71]);
  assign t[331] = (x[71]);
  assign t[332] = (x[74]);
  assign t[333] = (x[74]);
  assign t[334] = (x[77]);
  assign t[335] = (x[77]);
  assign t[336] = (x[80]);
  assign t[337] = (x[80]);
  assign t[338] = (x[83]);
  assign t[339] = (x[83]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = (x[86]);
  assign t[341] = (x[86]);
  assign t[342] = (x[89]);
  assign t[343] = (x[89]);
  assign t[344] = (x[92]);
  assign t[345] = (x[92]);
  assign t[346] = (x[95]);
  assign t[347] = (x[95]);
  assign t[34] = ~(t[148]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[54] | t[56]);
  assign t[37] = ~(t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = ~(t[151]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[152]);
  assign t[41] = ~(t[60] | t[61]);
  assign t[42] = ~(t[62] | t[63]);
  assign t[43] = ~(t[153] | t[64]);
  assign t[44] = t[23] ? x[33] : x[32];
  assign t[45] = ~(t[65] & t[66]);
  assign t[46] = ~(t[67] | t[68]);
  assign t[47] = ~(t[154] | t[69]);
  assign t[48] = ~(t[70] | t[71]);
  assign t[49] = ~(t[72] ^ t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] | t[75]);
  assign t[51] = ~(t[155] | t[76]);
  assign t[52] = ~(t[77] | t[78]);
  assign t[53] = ~(t[79] ^ t[80]);
  assign t[54] = ~(t[148]);
  assign t[55] = t[146] ? t[82] : t[81];
  assign t[56] = t[146] ? t[84] : t[83];
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[54]);
  assign t[59] = t[146] ? t[87] : t[83];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[156]);
  assign t[61] = ~(t[151] | t[152]);
  assign t[62] = ~(t[157]);
  assign t[63] = ~(t[158]);
  assign t[64] = ~(t[88] | t[89]);
  assign t[65] = ~(t[90] | t[36]);
  assign t[66] = ~(t[91] | t[92]);
  assign t[67] = ~(t[159]);
  assign t[68] = ~(t[160]);
  assign t[69] = ~(t[93] | t[94]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] | t[96]);
  assign t[71] = ~(t[161] | t[97]);
  assign t[72] = t[23] ? x[59] : x[58];
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[162]);
  assign t[75] = ~(t[163]);
  assign t[76] = ~(t[100] | t[101]);
  assign t[77] = ~(t[102] | t[103]);
  assign t[78] = ~(t[164] | t[104]);
  assign t[79] = t[105] ? x[70] : x[69];
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = ~(t[106] & t[107]);
  assign t[81] = ~(t[108] & t[109]);
  assign t[82] = ~(t[110] & t[109]);
  assign t[83] = ~(x[4] & t[111]);
  assign t[84] = ~(t[112] & t[109]);
  assign t[85] = ~(t[58] | t[113]);
  assign t[86] = ~(t[58] | t[114]);
  assign t[87] = ~(t[149] & t[112]);
  assign t[88] = ~(t[165]);
  assign t[89] = ~(t[157] | t[158]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = ~(t[54] | t[115]);
  assign t[91] = ~(t[116] & t[117]);
  assign t[92] = ~(t[118] & t[119]);
  assign t[93] = ~(t[166]);
  assign t[94] = ~(t[159] | t[160]);
  assign t[95] = ~(t[167]);
  assign t[96] = ~(t[168]);
  assign t[97] = ~(t[120] | t[121]);
  assign t[98] = ~(t[122] | t[86]);
  assign t[99] = ~(t[123] | t[124]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind261(x, y);
 input [97:0] x;
 output y;

 wire [347:0] t;
  assign t[0] = t[1] ? t[2] : t[145];
  assign t[100] = ~(t[169]);
  assign t[101] = ~(t[162] | t[163]);
  assign t[102] = ~(t[170]);
  assign t[103] = ~(t[171]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[34]);
  assign t[106] = ~(t[85] | t[127]);
  assign t[107] = ~(t[128]);
  assign t[108] = x[4] & t[147];
  assign t[109] = ~(t[149]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = ~(x[4] | t[147]);
  assign t[111] = ~(t[147] | t[149]);
  assign t[112] = ~(x[4] | t[129]);
  assign t[113] = t[146] ? t[130] : t[84];
  assign t[114] = t[146] ? t[81] : t[131];
  assign t[115] = t[146] ? t[81] : t[82];
  assign t[116] = ~(t[35] | t[132]);
  assign t[117] = ~(t[54] & t[133]);
  assign t[118] = ~(t[123] & t[134]);
  assign t[119] = t[54] | t[135];
  assign t[11] = ~(x[3]);
  assign t[120] = ~(t[172]);
  assign t[121] = ~(t[167] | t[168]);
  assign t[122] = ~(t[58] | t[136]);
  assign t[123] = t[149] & t[137];
  assign t[124] = ~(t[65]);
  assign t[125] = ~(t[173]);
  assign t[126] = ~(t[170] | t[171]);
  assign t[127] = ~(t[138] & t[65]);
  assign t[128] = ~(t[58] | t[139]);
  assign t[129] = ~(t[147]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(x[4] & t[140]);
  assign t[131] = ~(t[110] & t[149]);
  assign t[132] = ~(t[58] | t[141]);
  assign t[133] = ~(t[83] & t[87]);
  assign t[134] = t[110] | t[108];
  assign t[135] = t[146] ? t[83] : t[84];
  assign t[136] = t[146] ? t[83] : t[87];
  assign t[137] = ~(t[54] | t[146]);
  assign t[138] = ~(t[142] | t[91]);
  assign t[139] = t[146] ? t[82] : t[143];
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = ~(t[147] | t[109]);
  assign t[141] = t[146] ? t[84] : t[130];
  assign t[142] = ~(t[58] | t[144]);
  assign t[143] = ~(t[108] & t[149]);
  assign t[144] = t[146] ? t[143] : t[82];
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = ~(t[146] & t[147]);
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = (t[195]);
  assign t[167] = (t[196]);
  assign t[168] = (t[197]);
  assign t[169] = (t[198]);
  assign t[16] = ~(t[148] & t[149]);
  assign t[170] = (t[199]);
  assign t[171] = (t[200]);
  assign t[172] = (t[201]);
  assign t[173] = (t[202]);
  assign t[174] = t[203] ^ x[2];
  assign t[175] = t[204] ^ x[10];
  assign t[176] = t[205] ^ x[13];
  assign t[177] = t[206] ^ x[16];
  assign t[178] = t[207] ^ x[19];
  assign t[179] = t[208] ^ x[22];
  assign t[17] = t[23] ? x[7] : x[6];
  assign t[180] = t[209] ^ x[25];
  assign t[181] = t[210] ^ x[28];
  assign t[182] = t[211] ^ x[31];
  assign t[183] = t[212] ^ x[36];
  assign t[184] = t[213] ^ x[39];
  assign t[185] = t[214] ^ x[42];
  assign t[186] = t[215] ^ x[45];
  assign t[187] = t[216] ^ x[48];
  assign t[188] = t[217] ^ x[51];
  assign t[189] = t[218] ^ x[54];
  assign t[18] = ~(t[24] & t[25]);
  assign t[190] = t[219] ^ x[57];
  assign t[191] = t[220] ^ x[62];
  assign t[192] = t[221] ^ x[65];
  assign t[193] = t[222] ^ x[68];
  assign t[194] = t[223] ^ x[73];
  assign t[195] = t[224] ^ x[76];
  assign t[196] = t[225] ^ x[79];
  assign t[197] = t[226] ^ x[82];
  assign t[198] = t[227] ^ x[85];
  assign t[199] = t[228] ^ x[88];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[229] ^ x[91];
  assign t[201] = t[230] ^ x[94];
  assign t[202] = t[231] ^ x[97];
  assign t[203] = (t[232] & ~t[233]);
  assign t[204] = (t[234] & ~t[235]);
  assign t[205] = (t[236] & ~t[237]);
  assign t[206] = (t[238] & ~t[239]);
  assign t[207] = (t[240] & ~t[241]);
  assign t[208] = (t[242] & ~t[243]);
  assign t[209] = (t[244] & ~t[245]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (t[246] & ~t[247]);
  assign t[211] = (t[248] & ~t[249]);
  assign t[212] = (t[250] & ~t[251]);
  assign t[213] = (t[252] & ~t[253]);
  assign t[214] = (t[254] & ~t[255]);
  assign t[215] = (t[256] & ~t[257]);
  assign t[216] = (t[258] & ~t[259]);
  assign t[217] = (t[260] & ~t[261]);
  assign t[218] = (t[262] & ~t[263]);
  assign t[219] = (t[264] & ~t[265]);
  assign t[21] = x[4] ? t[31] : t[30];
  assign t[220] = (t[266] & ~t[267]);
  assign t[221] = (t[268] & ~t[269]);
  assign t[222] = (t[270] & ~t[271]);
  assign t[223] = (t[272] & ~t[273]);
  assign t[224] = (t[274] & ~t[275]);
  assign t[225] = (t[276] & ~t[277]);
  assign t[226] = (t[278] & ~t[279]);
  assign t[227] = (t[280] & ~t[281]);
  assign t[228] = (t[282] & ~t[283]);
  assign t[229] = (t[284] & ~t[285]);
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[230] = (t[286] & ~t[287]);
  assign t[231] = (t[288] & ~t[289]);
  assign t[232] = t[290] ^ x[2];
  assign t[233] = t[291] ^ x[1];
  assign t[234] = t[292] ^ x[10];
  assign t[235] = t[293] ^ x[9];
  assign t[236] = t[294] ^ x[13];
  assign t[237] = t[295] ^ x[12];
  assign t[238] = t[296] ^ x[16];
  assign t[239] = t[297] ^ x[15];
  assign t[23] = ~(t[34]);
  assign t[240] = t[298] ^ x[19];
  assign t[241] = t[299] ^ x[18];
  assign t[242] = t[300] ^ x[22];
  assign t[243] = t[301] ^ x[21];
  assign t[244] = t[302] ^ x[25];
  assign t[245] = t[303] ^ x[24];
  assign t[246] = t[304] ^ x[28];
  assign t[247] = t[305] ^ x[27];
  assign t[248] = t[306] ^ x[31];
  assign t[249] = t[307] ^ x[30];
  assign t[24] = ~(t[35] | t[36]);
  assign t[250] = t[308] ^ x[36];
  assign t[251] = t[309] ^ x[35];
  assign t[252] = t[310] ^ x[39];
  assign t[253] = t[311] ^ x[38];
  assign t[254] = t[312] ^ x[42];
  assign t[255] = t[313] ^ x[41];
  assign t[256] = t[314] ^ x[45];
  assign t[257] = t[315] ^ x[44];
  assign t[258] = t[316] ^ x[48];
  assign t[259] = t[317] ^ x[47];
  assign t[25] = ~(t[37] | t[38]);
  assign t[260] = t[318] ^ x[51];
  assign t[261] = t[319] ^ x[50];
  assign t[262] = t[320] ^ x[54];
  assign t[263] = t[321] ^ x[53];
  assign t[264] = t[322] ^ x[57];
  assign t[265] = t[323] ^ x[56];
  assign t[266] = t[324] ^ x[62];
  assign t[267] = t[325] ^ x[61];
  assign t[268] = t[326] ^ x[65];
  assign t[269] = t[327] ^ x[64];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[328] ^ x[68];
  assign t[271] = t[329] ^ x[67];
  assign t[272] = t[330] ^ x[73];
  assign t[273] = t[331] ^ x[72];
  assign t[274] = t[332] ^ x[76];
  assign t[275] = t[333] ^ x[75];
  assign t[276] = t[334] ^ x[79];
  assign t[277] = t[335] ^ x[78];
  assign t[278] = t[336] ^ x[82];
  assign t[279] = t[337] ^ x[81];
  assign t[27] = ~(t[150] | t[41]);
  assign t[280] = t[338] ^ x[85];
  assign t[281] = t[339] ^ x[84];
  assign t[282] = t[340] ^ x[88];
  assign t[283] = t[341] ^ x[87];
  assign t[284] = t[342] ^ x[91];
  assign t[285] = t[343] ^ x[90];
  assign t[286] = t[344] ^ x[94];
  assign t[287] = t[345] ^ x[93];
  assign t[288] = t[346] ^ x[97];
  assign t[289] = t[347] ^ x[96];
  assign t[28] = ~(t[42] | t[43]);
  assign t[290] = (x[0]);
  assign t[291] = (x[0]);
  assign t[292] = (x[8]);
  assign t[293] = (x[8]);
  assign t[294] = (x[11]);
  assign t[295] = (x[11]);
  assign t[296] = (x[14]);
  assign t[297] = (x[14]);
  assign t[298] = (x[17]);
  assign t[299] = (x[17]);
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[300] = (x[20]);
  assign t[301] = (x[20]);
  assign t[302] = (x[23]);
  assign t[303] = (x[23]);
  assign t[304] = (x[26]);
  assign t[305] = (x[26]);
  assign t[306] = (x[29]);
  assign t[307] = (x[29]);
  assign t[308] = (x[34]);
  assign t[309] = (x[34]);
  assign t[30] = ~(t[46] | t[47]);
  assign t[310] = (x[37]);
  assign t[311] = (x[37]);
  assign t[312] = (x[40]);
  assign t[313] = (x[40]);
  assign t[314] = (x[43]);
  assign t[315] = (x[43]);
  assign t[316] = (x[46]);
  assign t[317] = (x[46]);
  assign t[318] = (x[49]);
  assign t[319] = (x[49]);
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[320] = (x[52]);
  assign t[321] = (x[52]);
  assign t[322] = (x[55]);
  assign t[323] = (x[55]);
  assign t[324] = (x[60]);
  assign t[325] = (x[60]);
  assign t[326] = (x[63]);
  assign t[327] = (x[63]);
  assign t[328] = (x[66]);
  assign t[329] = (x[66]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[71]);
  assign t[331] = (x[71]);
  assign t[332] = (x[74]);
  assign t[333] = (x[74]);
  assign t[334] = (x[77]);
  assign t[335] = (x[77]);
  assign t[336] = (x[80]);
  assign t[337] = (x[80]);
  assign t[338] = (x[83]);
  assign t[339] = (x[83]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = (x[86]);
  assign t[341] = (x[86]);
  assign t[342] = (x[89]);
  assign t[343] = (x[89]);
  assign t[344] = (x[92]);
  assign t[345] = (x[92]);
  assign t[346] = (x[95]);
  assign t[347] = (x[95]);
  assign t[34] = ~(t[148]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[54] | t[56]);
  assign t[37] = ~(t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = ~(t[151]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[152]);
  assign t[41] = ~(t[60] | t[61]);
  assign t[42] = ~(t[62] | t[63]);
  assign t[43] = ~(t[153] | t[64]);
  assign t[44] = t[23] ? x[33] : x[32];
  assign t[45] = ~(t[65] & t[66]);
  assign t[46] = ~(t[67] | t[68]);
  assign t[47] = ~(t[154] | t[69]);
  assign t[48] = ~(t[70] | t[71]);
  assign t[49] = ~(t[72] ^ t[73]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[74] | t[75]);
  assign t[51] = ~(t[155] | t[76]);
  assign t[52] = ~(t[77] | t[78]);
  assign t[53] = ~(t[79] ^ t[80]);
  assign t[54] = ~(t[148]);
  assign t[55] = t[146] ? t[82] : t[81];
  assign t[56] = t[146] ? t[84] : t[83];
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[54]);
  assign t[59] = t[146] ? t[87] : t[83];
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[156]);
  assign t[61] = ~(t[151] | t[152]);
  assign t[62] = ~(t[157]);
  assign t[63] = ~(t[158]);
  assign t[64] = ~(t[88] | t[89]);
  assign t[65] = ~(t[90] | t[36]);
  assign t[66] = ~(t[91] | t[92]);
  assign t[67] = ~(t[159]);
  assign t[68] = ~(t[160]);
  assign t[69] = ~(t[93] | t[94]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] | t[96]);
  assign t[71] = ~(t[161] | t[97]);
  assign t[72] = t[23] ? x[59] : x[58];
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[162]);
  assign t[75] = ~(t[163]);
  assign t[76] = ~(t[100] | t[101]);
  assign t[77] = ~(t[102] | t[103]);
  assign t[78] = ~(t[164] | t[104]);
  assign t[79] = t[105] ? x[70] : x[69];
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = ~(t[106] & t[107]);
  assign t[81] = ~(t[108] & t[109]);
  assign t[82] = ~(t[110] & t[109]);
  assign t[83] = ~(x[4] & t[111]);
  assign t[84] = ~(t[112] & t[109]);
  assign t[85] = ~(t[58] | t[113]);
  assign t[86] = ~(t[58] | t[114]);
  assign t[87] = ~(t[149] & t[112]);
  assign t[88] = ~(t[165]);
  assign t[89] = ~(t[157] | t[158]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = ~(t[54] | t[115]);
  assign t[91] = ~(t[116] & t[117]);
  assign t[92] = ~(t[118] & t[119]);
  assign t[93] = ~(t[166]);
  assign t[94] = ~(t[159] | t[160]);
  assign t[95] = ~(t[167]);
  assign t[96] = ~(t[168]);
  assign t[97] = ~(t[120] | t[121]);
  assign t[98] = ~(t[122] | t[86]);
  assign t[99] = ~(t[123] | t[124]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [79:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[2] : t[64];
  assign t[100] = t[123] ^ x[50];
  assign t[101] = t[124] ^ x[55];
  assign t[102] = t[125] ^ x[58];
  assign t[103] = t[126] ^ x[61];
  assign t[104] = t[127] ^ x[64];
  assign t[105] = t[128] ^ x[67];
  assign t[106] = t[129] ^ x[70];
  assign t[107] = t[130] ^ x[73];
  assign t[108] = t[131] ^ x[76];
  assign t[109] = t[132] ^ x[79];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[133] & ~t[134]);
  assign t[111] = (t[135] & ~t[136]);
  assign t[112] = (t[137] & ~t[138]);
  assign t[113] = (t[139] & ~t[140]);
  assign t[114] = (t[141] & ~t[142]);
  assign t[115] = (t[143] & ~t[144]);
  assign t[116] = (t[145] & ~t[146]);
  assign t[117] = (t[147] & ~t[148]);
  assign t[118] = (t[149] & ~t[150]);
  assign t[119] = (t[151] & ~t[152]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[153] & ~t[154]);
  assign t[121] = (t[155] & ~t[156]);
  assign t[122] = (t[157] & ~t[158]);
  assign t[123] = (t[159] & ~t[160]);
  assign t[124] = (t[161] & ~t[162]);
  assign t[125] = (t[163] & ~t[164]);
  assign t[126] = (t[165] & ~t[166]);
  assign t[127] = (t[167] & ~t[168]);
  assign t[128] = (t[169] & ~t[170]);
  assign t[129] = (t[171] & ~t[172]);
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = (t[173] & ~t[174]);
  assign t[131] = (t[175] & ~t[176]);
  assign t[132] = (t[177] & ~t[178]);
  assign t[133] = t[179] ^ x[2];
  assign t[134] = t[180] ^ x[1];
  assign t[135] = t[181] ^ x[10];
  assign t[136] = t[182] ^ x[9];
  assign t[137] = t[183] ^ x[13];
  assign t[138] = t[184] ^ x[12];
  assign t[139] = t[185] ^ x[16];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[186] ^ x[15];
  assign t[141] = t[187] ^ x[19];
  assign t[142] = t[188] ^ x[18];
  assign t[143] = t[189] ^ x[22];
  assign t[144] = t[190] ^ x[21];
  assign t[145] = t[191] ^ x[25];
  assign t[146] = t[192] ^ x[24];
  assign t[147] = t[193] ^ x[30];
  assign t[148] = t[194] ^ x[29];
  assign t[149] = t[195] ^ x[33];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[196] ^ x[32];
  assign t[151] = t[197] ^ x[36];
  assign t[152] = t[198] ^ x[35];
  assign t[153] = t[199] ^ x[39];
  assign t[154] = t[200] ^ x[38];
  assign t[155] = t[201] ^ x[42];
  assign t[156] = t[202] ^ x[41];
  assign t[157] = t[203] ^ x[47];
  assign t[158] = t[204] ^ x[46];
  assign t[159] = t[205] ^ x[50];
  assign t[15] = ~(t[65] & t[66]);
  assign t[160] = t[206] ^ x[49];
  assign t[161] = t[207] ^ x[55];
  assign t[162] = t[208] ^ x[54];
  assign t[163] = t[209] ^ x[58];
  assign t[164] = t[210] ^ x[57];
  assign t[165] = t[211] ^ x[61];
  assign t[166] = t[212] ^ x[60];
  assign t[167] = t[213] ^ x[64];
  assign t[168] = t[214] ^ x[63];
  assign t[169] = t[215] ^ x[67];
  assign t[16] = ~(t[67] & t[68]);
  assign t[170] = t[216] ^ x[66];
  assign t[171] = t[217] ^ x[70];
  assign t[172] = t[218] ^ x[69];
  assign t[173] = t[219] ^ x[73];
  assign t[174] = t[220] ^ x[72];
  assign t[175] = t[221] ^ x[76];
  assign t[176] = t[222] ^ x[75];
  assign t[177] = t[223] ^ x[79];
  assign t[178] = t[224] ^ x[78];
  assign t[179] = (x[0]);
  assign t[17] = ~(t[22]);
  assign t[180] = (x[0]);
  assign t[181] = (x[8]);
  assign t[182] = (x[8]);
  assign t[183] = (x[11]);
  assign t[184] = (x[11]);
  assign t[185] = (x[14]);
  assign t[186] = (x[14]);
  assign t[187] = (x[17]);
  assign t[188] = (x[17]);
  assign t[189] = (x[20]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = (x[20]);
  assign t[191] = (x[23]);
  assign t[192] = (x[23]);
  assign t[193] = (x[28]);
  assign t[194] = (x[28]);
  assign t[195] = (x[31]);
  assign t[196] = (x[31]);
  assign t[197] = (x[34]);
  assign t[198] = (x[34]);
  assign t[199] = (x[37]);
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[37]);
  assign t[201] = (x[40]);
  assign t[202] = (x[40]);
  assign t[203] = (x[45]);
  assign t[204] = (x[45]);
  assign t[205] = (x[48]);
  assign t[206] = (x[48]);
  assign t[207] = (x[53]);
  assign t[208] = (x[53]);
  assign t[209] = (x[56]);
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = (x[56]);
  assign t[211] = (x[59]);
  assign t[212] = (x[59]);
  assign t[213] = (x[62]);
  assign t[214] = (x[62]);
  assign t[215] = (x[65]);
  assign t[216] = (x[65]);
  assign t[217] = (x[68]);
  assign t[218] = (x[68]);
  assign t[219] = (x[71]);
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = (x[71]);
  assign t[221] = (x[74]);
  assign t[222] = (x[74]);
  assign t[223] = (x[77]);
  assign t[224] = (x[77]);
  assign t[22] = ~(t[67]);
  assign t[23] = ~(t[69] & t[31]);
  assign t[24] = ~(t[70] & t[32]);
  assign t[25] = t[17] ? x[27] : x[26];
  assign t[26] = ~(t[33] & t[34]);
  assign t[27] = ~(t[35] & t[36]);
  assign t[28] = t[37] ^ t[38];
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[71]);
  assign t[32] = ~(t[71] & t[43]);
  assign t[33] = ~(t[72] & t[44]);
  assign t[34] = ~(t[73] & t[45]);
  assign t[35] = ~(t[74] & t[46]);
  assign t[36] = ~(t[75] & t[47]);
  assign t[37] = t[48] ? x[44] : x[43];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[76] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[77] & t[52]);
  assign t[41] = t[17] ? x[52] : x[51];
  assign t[42] = ~(t[53] & t[54]);
  assign t[43] = ~(t[69]);
  assign t[44] = ~(t[78]);
  assign t[45] = ~(t[78] & t[55]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[56]);
  assign t[48] = ~(t[22]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[82]);
  assign t[52] = ~(t[82] & t[59]);
  assign t[53] = ~(t[83] & t[60]);
  assign t[54] = ~(t[84] & t[61]);
  assign t[55] = ~(t[72]);
  assign t[56] = ~(t[74]);
  assign t[57] = ~(t[85]);
  assign t[58] = ~(t[85] & t[62]);
  assign t[59] = ~(t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[86]);
  assign t[61] = ~(t[86] & t[63]);
  assign t[62] = ~(t[80]);
  assign t[63] = ~(t[83]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = (t[107]);
  assign t[85] = (t[108]);
  assign t[86] = (t[109]);
  assign t[87] = t[110] ^ x[2];
  assign t[88] = t[111] ^ x[10];
  assign t[89] = t[112] ^ x[13];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = t[113] ^ x[16];
  assign t[91] = t[114] ^ x[19];
  assign t[92] = t[115] ^ x[22];
  assign t[93] = t[116] ^ x[25];
  assign t[94] = t[117] ^ x[30];
  assign t[95] = t[118] ^ x[33];
  assign t[96] = t[119] ^ x[36];
  assign t[97] = t[120] ^ x[39];
  assign t[98] = t[121] ^ x[42];
  assign t[99] = t[122] ^ x[47];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [79:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[2] : t[64];
  assign t[100] = t[123] ^ x[50];
  assign t[101] = t[124] ^ x[55];
  assign t[102] = t[125] ^ x[58];
  assign t[103] = t[126] ^ x[61];
  assign t[104] = t[127] ^ x[64];
  assign t[105] = t[128] ^ x[67];
  assign t[106] = t[129] ^ x[70];
  assign t[107] = t[130] ^ x[73];
  assign t[108] = t[131] ^ x[76];
  assign t[109] = t[132] ^ x[79];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[133] & ~t[134]);
  assign t[111] = (t[135] & ~t[136]);
  assign t[112] = (t[137] & ~t[138]);
  assign t[113] = (t[139] & ~t[140]);
  assign t[114] = (t[141] & ~t[142]);
  assign t[115] = (t[143] & ~t[144]);
  assign t[116] = (t[145] & ~t[146]);
  assign t[117] = (t[147] & ~t[148]);
  assign t[118] = (t[149] & ~t[150]);
  assign t[119] = (t[151] & ~t[152]);
  assign t[11] = ~(x[3]);
  assign t[120] = (t[153] & ~t[154]);
  assign t[121] = (t[155] & ~t[156]);
  assign t[122] = (t[157] & ~t[158]);
  assign t[123] = (t[159] & ~t[160]);
  assign t[124] = (t[161] & ~t[162]);
  assign t[125] = (t[163] & ~t[164]);
  assign t[126] = (t[165] & ~t[166]);
  assign t[127] = (t[167] & ~t[168]);
  assign t[128] = (t[169] & ~t[170]);
  assign t[129] = (t[171] & ~t[172]);
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = (t[173] & ~t[174]);
  assign t[131] = (t[175] & ~t[176]);
  assign t[132] = (t[177] & ~t[178]);
  assign t[133] = t[179] ^ x[2];
  assign t[134] = t[180] ^ x[1];
  assign t[135] = t[181] ^ x[10];
  assign t[136] = t[182] ^ x[9];
  assign t[137] = t[183] ^ x[13];
  assign t[138] = t[184] ^ x[12];
  assign t[139] = t[185] ^ x[16];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[186] ^ x[15];
  assign t[141] = t[187] ^ x[19];
  assign t[142] = t[188] ^ x[18];
  assign t[143] = t[189] ^ x[22];
  assign t[144] = t[190] ^ x[21];
  assign t[145] = t[191] ^ x[25];
  assign t[146] = t[192] ^ x[24];
  assign t[147] = t[193] ^ x[30];
  assign t[148] = t[194] ^ x[29];
  assign t[149] = t[195] ^ x[33];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[196] ^ x[32];
  assign t[151] = t[197] ^ x[36];
  assign t[152] = t[198] ^ x[35];
  assign t[153] = t[199] ^ x[39];
  assign t[154] = t[200] ^ x[38];
  assign t[155] = t[201] ^ x[42];
  assign t[156] = t[202] ^ x[41];
  assign t[157] = t[203] ^ x[47];
  assign t[158] = t[204] ^ x[46];
  assign t[159] = t[205] ^ x[50];
  assign t[15] = ~(t[65] & t[66]);
  assign t[160] = t[206] ^ x[49];
  assign t[161] = t[207] ^ x[55];
  assign t[162] = t[208] ^ x[54];
  assign t[163] = t[209] ^ x[58];
  assign t[164] = t[210] ^ x[57];
  assign t[165] = t[211] ^ x[61];
  assign t[166] = t[212] ^ x[60];
  assign t[167] = t[213] ^ x[64];
  assign t[168] = t[214] ^ x[63];
  assign t[169] = t[215] ^ x[67];
  assign t[16] = ~(t[67] & t[68]);
  assign t[170] = t[216] ^ x[66];
  assign t[171] = t[217] ^ x[70];
  assign t[172] = t[218] ^ x[69];
  assign t[173] = t[219] ^ x[73];
  assign t[174] = t[220] ^ x[72];
  assign t[175] = t[221] ^ x[76];
  assign t[176] = t[222] ^ x[75];
  assign t[177] = t[223] ^ x[79];
  assign t[178] = t[224] ^ x[78];
  assign t[179] = (x[0]);
  assign t[17] = ~(t[22]);
  assign t[180] = (x[0]);
  assign t[181] = (x[8]);
  assign t[182] = (x[8]);
  assign t[183] = (x[11]);
  assign t[184] = (x[11]);
  assign t[185] = (x[14]);
  assign t[186] = (x[14]);
  assign t[187] = (x[17]);
  assign t[188] = (x[17]);
  assign t[189] = (x[20]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = (x[20]);
  assign t[191] = (x[23]);
  assign t[192] = (x[23]);
  assign t[193] = (x[28]);
  assign t[194] = (x[28]);
  assign t[195] = (x[31]);
  assign t[196] = (x[31]);
  assign t[197] = (x[34]);
  assign t[198] = (x[34]);
  assign t[199] = (x[37]);
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[37]);
  assign t[201] = (x[40]);
  assign t[202] = (x[40]);
  assign t[203] = (x[45]);
  assign t[204] = (x[45]);
  assign t[205] = (x[48]);
  assign t[206] = (x[48]);
  assign t[207] = (x[53]);
  assign t[208] = (x[53]);
  assign t[209] = (x[56]);
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = (x[56]);
  assign t[211] = (x[59]);
  assign t[212] = (x[59]);
  assign t[213] = (x[62]);
  assign t[214] = (x[62]);
  assign t[215] = (x[65]);
  assign t[216] = (x[65]);
  assign t[217] = (x[68]);
  assign t[218] = (x[68]);
  assign t[219] = (x[71]);
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = (x[71]);
  assign t[221] = (x[74]);
  assign t[222] = (x[74]);
  assign t[223] = (x[77]);
  assign t[224] = (x[77]);
  assign t[22] = ~(t[67]);
  assign t[23] = ~(t[69] & t[31]);
  assign t[24] = ~(t[70] & t[32]);
  assign t[25] = t[17] ? x[27] : x[26];
  assign t[26] = ~(t[33] & t[34]);
  assign t[27] = ~(t[35] & t[36]);
  assign t[28] = t[37] ^ t[38];
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[71]);
  assign t[32] = ~(t[71] & t[43]);
  assign t[33] = ~(t[72] & t[44]);
  assign t[34] = ~(t[73] & t[45]);
  assign t[35] = ~(t[74] & t[46]);
  assign t[36] = ~(t[75] & t[47]);
  assign t[37] = t[48] ? x[44] : x[43];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[76] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[77] & t[52]);
  assign t[41] = t[17] ? x[52] : x[51];
  assign t[42] = ~(t[53] & t[54]);
  assign t[43] = ~(t[69]);
  assign t[44] = ~(t[78]);
  assign t[45] = ~(t[78] & t[55]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[56]);
  assign t[48] = ~(t[22]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[82]);
  assign t[52] = ~(t[82] & t[59]);
  assign t[53] = ~(t[83] & t[60]);
  assign t[54] = ~(t[84] & t[61]);
  assign t[55] = ~(t[72]);
  assign t[56] = ~(t[74]);
  assign t[57] = ~(t[85]);
  assign t[58] = ~(t[85] & t[62]);
  assign t[59] = ~(t[76]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[86]);
  assign t[61] = ~(t[86] & t[63]);
  assign t[62] = ~(t[80]);
  assign t[63] = ~(t[83]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = (t[107]);
  assign t[85] = (t[108]);
  assign t[86] = (t[109]);
  assign t[87] = t[110] ^ x[2];
  assign t[88] = t[111] ^ x[10];
  assign t[89] = t[112] ^ x[13];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = t[113] ^ x[16];
  assign t[91] = t[114] ^ x[19];
  assign t[92] = t[115] ^ x[22];
  assign t[93] = t[116] ^ x[25];
  assign t[94] = t[117] ^ x[30];
  assign t[95] = t[118] ^ x[33];
  assign t[96] = t[119] ^ x[36];
  assign t[97] = t[120] ^ x[39];
  assign t[98] = t[121] ^ x[42];
  assign t[99] = t[122] ^ x[47];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [97:0] x;
 output y;

 wire [278:0] t;
  assign t[0] = t[1] ? t[2] : t[76];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = (t[131]);
  assign t[103] = (t[132]);
  assign t[104] = (t[133]);
  assign t[105] = t[134] ^ x[2];
  assign t[106] = t[135] ^ x[10];
  assign t[107] = t[136] ^ x[13];
  assign t[108] = t[137] ^ x[16];
  assign t[109] = t[138] ^ x[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[22];
  assign t[111] = t[140] ^ x[27];
  assign t[112] = t[141] ^ x[30];
  assign t[113] = t[142] ^ x[33];
  assign t[114] = t[143] ^ x[36];
  assign t[115] = t[144] ^ x[41];
  assign t[116] = t[145] ^ x[46];
  assign t[117] = t[146] ^ x[49];
  assign t[118] = t[147] ^ x[52];
  assign t[119] = t[148] ^ x[55];
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ^ x[58];
  assign t[121] = t[150] ^ x[61];
  assign t[122] = t[151] ^ x[64];
  assign t[123] = t[152] ^ x[67];
  assign t[124] = t[153] ^ x[70];
  assign t[125] = t[154] ^ x[73];
  assign t[126] = t[155] ^ x[76];
  assign t[127] = t[156] ^ x[79];
  assign t[128] = t[157] ^ x[82];
  assign t[129] = t[158] ^ x[85];
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = t[159] ^ x[88];
  assign t[131] = t[160] ^ x[91];
  assign t[132] = t[161] ^ x[94];
  assign t[133] = t[162] ^ x[97];
  assign t[134] = (t[163] & ~t[164]);
  assign t[135] = (t[165] & ~t[166]);
  assign t[136] = (t[167] & ~t[168]);
  assign t[137] = (t[169] & ~t[170]);
  assign t[138] = (t[171] & ~t[172]);
  assign t[139] = (t[173] & ~t[174]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (t[175] & ~t[176]);
  assign t[141] = (t[177] & ~t[178]);
  assign t[142] = (t[179] & ~t[180]);
  assign t[143] = (t[181] & ~t[182]);
  assign t[144] = (t[183] & ~t[184]);
  assign t[145] = (t[185] & ~t[186]);
  assign t[146] = (t[187] & ~t[188]);
  assign t[147] = (t[189] & ~t[190]);
  assign t[148] = (t[191] & ~t[192]);
  assign t[149] = (t[193] & ~t[194]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (t[195] & ~t[196]);
  assign t[151] = (t[197] & ~t[198]);
  assign t[152] = (t[199] & ~t[200]);
  assign t[153] = (t[201] & ~t[202]);
  assign t[154] = (t[203] & ~t[204]);
  assign t[155] = (t[205] & ~t[206]);
  assign t[156] = (t[207] & ~t[208]);
  assign t[157] = (t[209] & ~t[210]);
  assign t[158] = (t[211] & ~t[212]);
  assign t[159] = (t[213] & ~t[214]);
  assign t[15] = ~(t[77] & t[78]);
  assign t[160] = (t[215] & ~t[216]);
  assign t[161] = (t[217] & ~t[218]);
  assign t[162] = (t[219] & ~t[220]);
  assign t[163] = t[221] ^ x[2];
  assign t[164] = t[222] ^ x[1];
  assign t[165] = t[223] ^ x[10];
  assign t[166] = t[224] ^ x[9];
  assign t[167] = t[225] ^ x[13];
  assign t[168] = t[226] ^ x[12];
  assign t[169] = t[227] ^ x[16];
  assign t[16] = ~(t[79] & t[80]);
  assign t[170] = t[228] ^ x[15];
  assign t[171] = t[229] ^ x[19];
  assign t[172] = t[230] ^ x[18];
  assign t[173] = t[231] ^ x[22];
  assign t[174] = t[232] ^ x[21];
  assign t[175] = t[233] ^ x[27];
  assign t[176] = t[234] ^ x[26];
  assign t[177] = t[235] ^ x[30];
  assign t[178] = t[236] ^ x[29];
  assign t[179] = t[237] ^ x[33];
  assign t[17] = ~(t[22]);
  assign t[180] = t[238] ^ x[32];
  assign t[181] = t[239] ^ x[36];
  assign t[182] = t[240] ^ x[35];
  assign t[183] = t[241] ^ x[41];
  assign t[184] = t[242] ^ x[40];
  assign t[185] = t[243] ^ x[46];
  assign t[186] = t[244] ^ x[45];
  assign t[187] = t[245] ^ x[49];
  assign t[188] = t[246] ^ x[48];
  assign t[189] = t[247] ^ x[52];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[248] ^ x[51];
  assign t[191] = t[249] ^ x[55];
  assign t[192] = t[250] ^ x[54];
  assign t[193] = t[251] ^ x[58];
  assign t[194] = t[252] ^ x[57];
  assign t[195] = t[253] ^ x[61];
  assign t[196] = t[254] ^ x[60];
  assign t[197] = t[255] ^ x[64];
  assign t[198] = t[256] ^ x[63];
  assign t[199] = t[257] ^ x[67];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[258] ^ x[66];
  assign t[201] = t[259] ^ x[70];
  assign t[202] = t[260] ^ x[69];
  assign t[203] = t[261] ^ x[73];
  assign t[204] = t[262] ^ x[72];
  assign t[205] = t[263] ^ x[76];
  assign t[206] = t[264] ^ x[75];
  assign t[207] = t[265] ^ x[79];
  assign t[208] = t[266] ^ x[78];
  assign t[209] = t[267] ^ x[82];
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = t[268] ^ x[81];
  assign t[211] = t[269] ^ x[85];
  assign t[212] = t[270] ^ x[84];
  assign t[213] = t[271] ^ x[88];
  assign t[214] = t[272] ^ x[87];
  assign t[215] = t[273] ^ x[91];
  assign t[216] = t[274] ^ x[90];
  assign t[217] = t[275] ^ x[94];
  assign t[218] = t[276] ^ x[93];
  assign t[219] = t[277] ^ x[97];
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = t[278] ^ x[96];
  assign t[221] = (x[0]);
  assign t[222] = (x[0]);
  assign t[223] = (x[8]);
  assign t[224] = (x[8]);
  assign t[225] = (x[11]);
  assign t[226] = (x[11]);
  assign t[227] = (x[14]);
  assign t[228] = (x[14]);
  assign t[229] = (x[17]);
  assign t[22] = ~(t[79]);
  assign t[230] = (x[17]);
  assign t[231] = (x[20]);
  assign t[232] = (x[20]);
  assign t[233] = (x[25]);
  assign t[234] = (x[25]);
  assign t[235] = (x[28]);
  assign t[236] = (x[28]);
  assign t[237] = (x[31]);
  assign t[238] = (x[31]);
  assign t[239] = (x[34]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[34]);
  assign t[241] = (x[39]);
  assign t[242] = (x[39]);
  assign t[243] = (x[44]);
  assign t[244] = (x[44]);
  assign t[245] = (x[47]);
  assign t[246] = (x[47]);
  assign t[247] = (x[50]);
  assign t[248] = (x[50]);
  assign t[249] = (x[53]);
  assign t[24] = ~(t[33] & t[81]);
  assign t[250] = (x[53]);
  assign t[251] = (x[56]);
  assign t[252] = (x[56]);
  assign t[253] = (x[59]);
  assign t[254] = (x[59]);
  assign t[255] = (x[62]);
  assign t[256] = (x[62]);
  assign t[257] = (x[65]);
  assign t[258] = (x[65]);
  assign t[259] = (x[68]);
  assign t[25] = t[17] ? x[24] : x[23];
  assign t[260] = (x[68]);
  assign t[261] = (x[71]);
  assign t[262] = (x[71]);
  assign t[263] = (x[74]);
  assign t[264] = (x[74]);
  assign t[265] = (x[77]);
  assign t[266] = (x[77]);
  assign t[267] = (x[80]);
  assign t[268] = (x[80]);
  assign t[269] = (x[83]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[270] = (x[83]);
  assign t[271] = (x[86]);
  assign t[272] = (x[86]);
  assign t[273] = (x[89]);
  assign t[274] = (x[89]);
  assign t[275] = (x[92]);
  assign t[276] = (x[92]);
  assign t[277] = (x[95]);
  assign t[278] = (x[95]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[82]);
  assign t[32] = ~(t[83]);
  assign t[33] = ~(t[44] & t[45]);
  assign t[34] = ~(t[46] & t[47]);
  assign t[35] = ~(t[48] & t[84]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[51] & t[85]);
  assign t[38] = t[52] ? x[38] : x[37];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[86]);
  assign t[42] = t[17] ? x[43] : x[42];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[83] & t[82]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[89]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[90]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[91]);
  assign t[51] = ~(t[62] & t[63]);
  assign t[52] = ~(t[22]);
  assign t[53] = ~(t[64] & t[65]);
  assign t[54] = ~(t[66] & t[92]);
  assign t[55] = ~(t[93]);
  assign t[56] = ~(t[94]);
  assign t[57] = ~(t[67] & t[68]);
  assign t[58] = ~(t[69] & t[70]);
  assign t[59] = ~(t[71] & t[95]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[89] & t[88]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[91] & t[90]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[72] & t[73]);
  assign t[67] = ~(t[94] & t[93]);
  assign t[68] = ~(t[100]);
  assign t[69] = ~(t[101]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[102]);
  assign t[71] = ~(t[74] & t[75]);
  assign t[72] = ~(t[99] & t[98]);
  assign t[73] = ~(t[103]);
  assign t[74] = ~(t[102] & t[101]);
  assign t[75] = ~(t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [97:0] x;
 output y;

 wire [278:0] t;
  assign t[0] = t[1] ? t[2] : t[76];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = (t[131]);
  assign t[103] = (t[132]);
  assign t[104] = (t[133]);
  assign t[105] = t[134] ^ x[2];
  assign t[106] = t[135] ^ x[10];
  assign t[107] = t[136] ^ x[13];
  assign t[108] = t[137] ^ x[16];
  assign t[109] = t[138] ^ x[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[22];
  assign t[111] = t[140] ^ x[27];
  assign t[112] = t[141] ^ x[30];
  assign t[113] = t[142] ^ x[33];
  assign t[114] = t[143] ^ x[36];
  assign t[115] = t[144] ^ x[41];
  assign t[116] = t[145] ^ x[46];
  assign t[117] = t[146] ^ x[49];
  assign t[118] = t[147] ^ x[52];
  assign t[119] = t[148] ^ x[55];
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ^ x[58];
  assign t[121] = t[150] ^ x[61];
  assign t[122] = t[151] ^ x[64];
  assign t[123] = t[152] ^ x[67];
  assign t[124] = t[153] ^ x[70];
  assign t[125] = t[154] ^ x[73];
  assign t[126] = t[155] ^ x[76];
  assign t[127] = t[156] ^ x[79];
  assign t[128] = t[157] ^ x[82];
  assign t[129] = t[158] ^ x[85];
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = t[159] ^ x[88];
  assign t[131] = t[160] ^ x[91];
  assign t[132] = t[161] ^ x[94];
  assign t[133] = t[162] ^ x[97];
  assign t[134] = (t[163] & ~t[164]);
  assign t[135] = (t[165] & ~t[166]);
  assign t[136] = (t[167] & ~t[168]);
  assign t[137] = (t[169] & ~t[170]);
  assign t[138] = (t[171] & ~t[172]);
  assign t[139] = (t[173] & ~t[174]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (t[175] & ~t[176]);
  assign t[141] = (t[177] & ~t[178]);
  assign t[142] = (t[179] & ~t[180]);
  assign t[143] = (t[181] & ~t[182]);
  assign t[144] = (t[183] & ~t[184]);
  assign t[145] = (t[185] & ~t[186]);
  assign t[146] = (t[187] & ~t[188]);
  assign t[147] = (t[189] & ~t[190]);
  assign t[148] = (t[191] & ~t[192]);
  assign t[149] = (t[193] & ~t[194]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (t[195] & ~t[196]);
  assign t[151] = (t[197] & ~t[198]);
  assign t[152] = (t[199] & ~t[200]);
  assign t[153] = (t[201] & ~t[202]);
  assign t[154] = (t[203] & ~t[204]);
  assign t[155] = (t[205] & ~t[206]);
  assign t[156] = (t[207] & ~t[208]);
  assign t[157] = (t[209] & ~t[210]);
  assign t[158] = (t[211] & ~t[212]);
  assign t[159] = (t[213] & ~t[214]);
  assign t[15] = ~(t[77] & t[78]);
  assign t[160] = (t[215] & ~t[216]);
  assign t[161] = (t[217] & ~t[218]);
  assign t[162] = (t[219] & ~t[220]);
  assign t[163] = t[221] ^ x[2];
  assign t[164] = t[222] ^ x[1];
  assign t[165] = t[223] ^ x[10];
  assign t[166] = t[224] ^ x[9];
  assign t[167] = t[225] ^ x[13];
  assign t[168] = t[226] ^ x[12];
  assign t[169] = t[227] ^ x[16];
  assign t[16] = ~(t[79] & t[80]);
  assign t[170] = t[228] ^ x[15];
  assign t[171] = t[229] ^ x[19];
  assign t[172] = t[230] ^ x[18];
  assign t[173] = t[231] ^ x[22];
  assign t[174] = t[232] ^ x[21];
  assign t[175] = t[233] ^ x[27];
  assign t[176] = t[234] ^ x[26];
  assign t[177] = t[235] ^ x[30];
  assign t[178] = t[236] ^ x[29];
  assign t[179] = t[237] ^ x[33];
  assign t[17] = ~(t[22]);
  assign t[180] = t[238] ^ x[32];
  assign t[181] = t[239] ^ x[36];
  assign t[182] = t[240] ^ x[35];
  assign t[183] = t[241] ^ x[41];
  assign t[184] = t[242] ^ x[40];
  assign t[185] = t[243] ^ x[46];
  assign t[186] = t[244] ^ x[45];
  assign t[187] = t[245] ^ x[49];
  assign t[188] = t[246] ^ x[48];
  assign t[189] = t[247] ^ x[52];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[248] ^ x[51];
  assign t[191] = t[249] ^ x[55];
  assign t[192] = t[250] ^ x[54];
  assign t[193] = t[251] ^ x[58];
  assign t[194] = t[252] ^ x[57];
  assign t[195] = t[253] ^ x[61];
  assign t[196] = t[254] ^ x[60];
  assign t[197] = t[255] ^ x[64];
  assign t[198] = t[256] ^ x[63];
  assign t[199] = t[257] ^ x[67];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[258] ^ x[66];
  assign t[201] = t[259] ^ x[70];
  assign t[202] = t[260] ^ x[69];
  assign t[203] = t[261] ^ x[73];
  assign t[204] = t[262] ^ x[72];
  assign t[205] = t[263] ^ x[76];
  assign t[206] = t[264] ^ x[75];
  assign t[207] = t[265] ^ x[79];
  assign t[208] = t[266] ^ x[78];
  assign t[209] = t[267] ^ x[82];
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = t[268] ^ x[81];
  assign t[211] = t[269] ^ x[85];
  assign t[212] = t[270] ^ x[84];
  assign t[213] = t[271] ^ x[88];
  assign t[214] = t[272] ^ x[87];
  assign t[215] = t[273] ^ x[91];
  assign t[216] = t[274] ^ x[90];
  assign t[217] = t[275] ^ x[94];
  assign t[218] = t[276] ^ x[93];
  assign t[219] = t[277] ^ x[97];
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = t[278] ^ x[96];
  assign t[221] = (x[0]);
  assign t[222] = (x[0]);
  assign t[223] = (x[8]);
  assign t[224] = (x[8]);
  assign t[225] = (x[11]);
  assign t[226] = (x[11]);
  assign t[227] = (x[14]);
  assign t[228] = (x[14]);
  assign t[229] = (x[17]);
  assign t[22] = ~(t[79]);
  assign t[230] = (x[17]);
  assign t[231] = (x[20]);
  assign t[232] = (x[20]);
  assign t[233] = (x[25]);
  assign t[234] = (x[25]);
  assign t[235] = (x[28]);
  assign t[236] = (x[28]);
  assign t[237] = (x[31]);
  assign t[238] = (x[31]);
  assign t[239] = (x[34]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[34]);
  assign t[241] = (x[39]);
  assign t[242] = (x[39]);
  assign t[243] = (x[44]);
  assign t[244] = (x[44]);
  assign t[245] = (x[47]);
  assign t[246] = (x[47]);
  assign t[247] = (x[50]);
  assign t[248] = (x[50]);
  assign t[249] = (x[53]);
  assign t[24] = ~(t[33] & t[81]);
  assign t[250] = (x[53]);
  assign t[251] = (x[56]);
  assign t[252] = (x[56]);
  assign t[253] = (x[59]);
  assign t[254] = (x[59]);
  assign t[255] = (x[62]);
  assign t[256] = (x[62]);
  assign t[257] = (x[65]);
  assign t[258] = (x[65]);
  assign t[259] = (x[68]);
  assign t[25] = t[17] ? x[24] : x[23];
  assign t[260] = (x[68]);
  assign t[261] = (x[71]);
  assign t[262] = (x[71]);
  assign t[263] = (x[74]);
  assign t[264] = (x[74]);
  assign t[265] = (x[77]);
  assign t[266] = (x[77]);
  assign t[267] = (x[80]);
  assign t[268] = (x[80]);
  assign t[269] = (x[83]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[270] = (x[83]);
  assign t[271] = (x[86]);
  assign t[272] = (x[86]);
  assign t[273] = (x[89]);
  assign t[274] = (x[89]);
  assign t[275] = (x[92]);
  assign t[276] = (x[92]);
  assign t[277] = (x[95]);
  assign t[278] = (x[95]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[82]);
  assign t[32] = ~(t[83]);
  assign t[33] = ~(t[44] & t[45]);
  assign t[34] = ~(t[46] & t[47]);
  assign t[35] = ~(t[48] & t[84]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[51] & t[85]);
  assign t[38] = t[52] ? x[38] : x[37];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[86]);
  assign t[42] = t[17] ? x[43] : x[42];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[83] & t[82]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[89]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[90]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[91]);
  assign t[51] = ~(t[62] & t[63]);
  assign t[52] = ~(t[22]);
  assign t[53] = ~(t[64] & t[65]);
  assign t[54] = ~(t[66] & t[92]);
  assign t[55] = ~(t[93]);
  assign t[56] = ~(t[94]);
  assign t[57] = ~(t[67] & t[68]);
  assign t[58] = ~(t[69] & t[70]);
  assign t[59] = ~(t[71] & t[95]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[89] & t[88]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[91] & t[90]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[72] & t[73]);
  assign t[67] = ~(t[94] & t[93]);
  assign t[68] = ~(t[100]);
  assign t[69] = ~(t[101]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[102]);
  assign t[71] = ~(t[74] & t[75]);
  assign t[72] = ~(t[99] & t[98]);
  assign t[73] = ~(t[103]);
  assign t[74] = ~(t[102] & t[101]);
  assign t[75] = ~(t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind266(x, y);
 input [97:0] x;
 output y;

 wire [272:0] t;
  assign t[0] = t[1] ? t[2] : t[70];
  assign t[100] = t[129] ^ x[10];
  assign t[101] = t[130] ^ x[13];
  assign t[102] = t[131] ^ x[16];
  assign t[103] = t[132] ^ x[19];
  assign t[104] = t[133] ^ x[22];
  assign t[105] = t[134] ^ x[27];
  assign t[106] = t[135] ^ x[30];
  assign t[107] = t[136] ^ x[33];
  assign t[108] = t[137] ^ x[36];
  assign t[109] = t[138] ^ x[41];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[46];
  assign t[111] = t[140] ^ x[49];
  assign t[112] = t[141] ^ x[52];
  assign t[113] = t[142] ^ x[55];
  assign t[114] = t[143] ^ x[58];
  assign t[115] = t[144] ^ x[61];
  assign t[116] = t[145] ^ x[64];
  assign t[117] = t[146] ^ x[67];
  assign t[118] = t[147] ^ x[70];
  assign t[119] = t[148] ^ x[73];
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ^ x[76];
  assign t[121] = t[150] ^ x[79];
  assign t[122] = t[151] ^ x[82];
  assign t[123] = t[152] ^ x[85];
  assign t[124] = t[153] ^ x[88];
  assign t[125] = t[154] ^ x[91];
  assign t[126] = t[155] ^ x[94];
  assign t[127] = t[156] ^ x[97];
  assign t[128] = (t[157] & ~t[158]);
  assign t[129] = (t[159] & ~t[160]);
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = (t[161] & ~t[162]);
  assign t[131] = (t[163] & ~t[164]);
  assign t[132] = (t[165] & ~t[166]);
  assign t[133] = (t[167] & ~t[168]);
  assign t[134] = (t[169] & ~t[170]);
  assign t[135] = (t[171] & ~t[172]);
  assign t[136] = (t[173] & ~t[174]);
  assign t[137] = (t[175] & ~t[176]);
  assign t[138] = (t[177] & ~t[178]);
  assign t[139] = (t[179] & ~t[180]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (t[181] & ~t[182]);
  assign t[141] = (t[183] & ~t[184]);
  assign t[142] = (t[185] & ~t[186]);
  assign t[143] = (t[187] & ~t[188]);
  assign t[144] = (t[189] & ~t[190]);
  assign t[145] = (t[191] & ~t[192]);
  assign t[146] = (t[193] & ~t[194]);
  assign t[147] = (t[195] & ~t[196]);
  assign t[148] = (t[197] & ~t[198]);
  assign t[149] = (t[199] & ~t[200]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (t[201] & ~t[202]);
  assign t[151] = (t[203] & ~t[204]);
  assign t[152] = (t[205] & ~t[206]);
  assign t[153] = (t[207] & ~t[208]);
  assign t[154] = (t[209] & ~t[210]);
  assign t[155] = (t[211] & ~t[212]);
  assign t[156] = (t[213] & ~t[214]);
  assign t[157] = t[215] ^ x[2];
  assign t[158] = t[216] ^ x[1];
  assign t[159] = t[217] ^ x[10];
  assign t[15] = ~(t[71] & t[72]);
  assign t[160] = t[218] ^ x[9];
  assign t[161] = t[219] ^ x[13];
  assign t[162] = t[220] ^ x[12];
  assign t[163] = t[221] ^ x[16];
  assign t[164] = t[222] ^ x[15];
  assign t[165] = t[223] ^ x[19];
  assign t[166] = t[224] ^ x[18];
  assign t[167] = t[225] ^ x[22];
  assign t[168] = t[226] ^ x[21];
  assign t[169] = t[227] ^ x[27];
  assign t[16] = ~(t[73] & t[74]);
  assign t[170] = t[228] ^ x[26];
  assign t[171] = t[229] ^ x[30];
  assign t[172] = t[230] ^ x[29];
  assign t[173] = t[231] ^ x[33];
  assign t[174] = t[232] ^ x[32];
  assign t[175] = t[233] ^ x[36];
  assign t[176] = t[234] ^ x[35];
  assign t[177] = t[235] ^ x[41];
  assign t[178] = t[236] ^ x[40];
  assign t[179] = t[237] ^ x[46];
  assign t[17] = ~(t[22]);
  assign t[180] = t[238] ^ x[45];
  assign t[181] = t[239] ^ x[49];
  assign t[182] = t[240] ^ x[48];
  assign t[183] = t[241] ^ x[52];
  assign t[184] = t[242] ^ x[51];
  assign t[185] = t[243] ^ x[55];
  assign t[186] = t[244] ^ x[54];
  assign t[187] = t[245] ^ x[58];
  assign t[188] = t[246] ^ x[57];
  assign t[189] = t[247] ^ x[61];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[248] ^ x[60];
  assign t[191] = t[249] ^ x[64];
  assign t[192] = t[250] ^ x[63];
  assign t[193] = t[251] ^ x[67];
  assign t[194] = t[252] ^ x[66];
  assign t[195] = t[253] ^ x[70];
  assign t[196] = t[254] ^ x[69];
  assign t[197] = t[255] ^ x[73];
  assign t[198] = t[256] ^ x[72];
  assign t[199] = t[257] ^ x[76];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[258] ^ x[75];
  assign t[201] = t[259] ^ x[79];
  assign t[202] = t[260] ^ x[78];
  assign t[203] = t[261] ^ x[82];
  assign t[204] = t[262] ^ x[81];
  assign t[205] = t[263] ^ x[85];
  assign t[206] = t[264] ^ x[84];
  assign t[207] = t[265] ^ x[88];
  assign t[208] = t[266] ^ x[87];
  assign t[209] = t[267] ^ x[91];
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = t[268] ^ x[90];
  assign t[211] = t[269] ^ x[94];
  assign t[212] = t[270] ^ x[93];
  assign t[213] = t[271] ^ x[97];
  assign t[214] = t[272] ^ x[96];
  assign t[215] = (x[0]);
  assign t[216] = (x[0]);
  assign t[217] = (x[8]);
  assign t[218] = (x[8]);
  assign t[219] = (x[11]);
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = (x[11]);
  assign t[221] = (x[14]);
  assign t[222] = (x[14]);
  assign t[223] = (x[17]);
  assign t[224] = (x[17]);
  assign t[225] = (x[20]);
  assign t[226] = (x[20]);
  assign t[227] = (x[25]);
  assign t[228] = (x[25]);
  assign t[229] = (x[28]);
  assign t[22] = ~(t[73]);
  assign t[230] = (x[28]);
  assign t[231] = (x[31]);
  assign t[232] = (x[31]);
  assign t[233] = (x[34]);
  assign t[234] = (x[34]);
  assign t[235] = (x[39]);
  assign t[236] = (x[39]);
  assign t[237] = (x[44]);
  assign t[238] = (x[44]);
  assign t[239] = (x[47]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[47]);
  assign t[241] = (x[50]);
  assign t[242] = (x[50]);
  assign t[243] = (x[53]);
  assign t[244] = (x[53]);
  assign t[245] = (x[56]);
  assign t[246] = (x[56]);
  assign t[247] = (x[59]);
  assign t[248] = (x[59]);
  assign t[249] = (x[62]);
  assign t[24] = t[33] | t[75];
  assign t[250] = (x[62]);
  assign t[251] = (x[65]);
  assign t[252] = (x[65]);
  assign t[253] = (x[68]);
  assign t[254] = (x[68]);
  assign t[255] = (x[71]);
  assign t[256] = (x[71]);
  assign t[257] = (x[74]);
  assign t[258] = (x[74]);
  assign t[259] = (x[77]);
  assign t[25] = t[17] ? x[24] : x[23];
  assign t[260] = (x[77]);
  assign t[261] = (x[80]);
  assign t[262] = (x[80]);
  assign t[263] = (x[83]);
  assign t[264] = (x[83]);
  assign t[265] = (x[86]);
  assign t[266] = (x[86]);
  assign t[267] = (x[89]);
  assign t[268] = (x[89]);
  assign t[269] = (x[92]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[270] = (x[92]);
  assign t[271] = (x[95]);
  assign t[272] = (x[95]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[76]);
  assign t[32] = ~(t[77]);
  assign t[33] = ~(t[44] | t[31]);
  assign t[34] = ~(t[45] & t[46]);
  assign t[35] = t[47] | t[78];
  assign t[36] = ~(t[48] & t[49]);
  assign t[37] = t[50] | t[79];
  assign t[38] = t[51] ? x[38] : x[37];
  assign t[39] = ~(t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[80];
  assign t[42] = t[17] ? x[43] : x[42];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[83]);
  assign t[47] = ~(t[59] | t[45]);
  assign t[48] = ~(t[84]);
  assign t[49] = ~(t[85]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[60] | t[48]);
  assign t[51] = ~(t[22]);
  assign t[52] = ~(t[61] & t[62]);
  assign t[53] = t[63] | t[86];
  assign t[54] = ~(t[87]);
  assign t[55] = ~(t[88]);
  assign t[56] = ~(t[64] | t[54]);
  assign t[57] = ~(t[65] & t[66]);
  assign t[58] = t[67] | t[89];
  assign t[59] = ~(t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[92]);
  assign t[62] = ~(t[93]);
  assign t[63] = ~(t[68] | t[61]);
  assign t[64] = ~(t[94]);
  assign t[65] = ~(t[95]);
  assign t[66] = ~(t[96]);
  assign t[67] = ~(t[69] | t[65]);
  assign t[68] = ~(t[97]);
  assign t[69] = ~(t[98]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = t[128] ^ x[2];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [97:0] x;
 output y;

 wire [272:0] t;
  assign t[0] = t[1] ? t[2] : t[70];
  assign t[100] = t[129] ^ x[10];
  assign t[101] = t[130] ^ x[13];
  assign t[102] = t[131] ^ x[16];
  assign t[103] = t[132] ^ x[19];
  assign t[104] = t[133] ^ x[22];
  assign t[105] = t[134] ^ x[27];
  assign t[106] = t[135] ^ x[30];
  assign t[107] = t[136] ^ x[33];
  assign t[108] = t[137] ^ x[36];
  assign t[109] = t[138] ^ x[41];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[46];
  assign t[111] = t[140] ^ x[49];
  assign t[112] = t[141] ^ x[52];
  assign t[113] = t[142] ^ x[55];
  assign t[114] = t[143] ^ x[58];
  assign t[115] = t[144] ^ x[61];
  assign t[116] = t[145] ^ x[64];
  assign t[117] = t[146] ^ x[67];
  assign t[118] = t[147] ^ x[70];
  assign t[119] = t[148] ^ x[73];
  assign t[11] = ~(x[3]);
  assign t[120] = t[149] ^ x[76];
  assign t[121] = t[150] ^ x[79];
  assign t[122] = t[151] ^ x[82];
  assign t[123] = t[152] ^ x[85];
  assign t[124] = t[153] ^ x[88];
  assign t[125] = t[154] ^ x[91];
  assign t[126] = t[155] ^ x[94];
  assign t[127] = t[156] ^ x[97];
  assign t[128] = (t[157] & ~t[158]);
  assign t[129] = (t[159] & ~t[160]);
  assign t[12] = t[17] ? x[7] : x[6];
  assign t[130] = (t[161] & ~t[162]);
  assign t[131] = (t[163] & ~t[164]);
  assign t[132] = (t[165] & ~t[166]);
  assign t[133] = (t[167] & ~t[168]);
  assign t[134] = (t[169] & ~t[170]);
  assign t[135] = (t[171] & ~t[172]);
  assign t[136] = (t[173] & ~t[174]);
  assign t[137] = (t[175] & ~t[176]);
  assign t[138] = (t[177] & ~t[178]);
  assign t[139] = (t[179] & ~t[180]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (t[181] & ~t[182]);
  assign t[141] = (t[183] & ~t[184]);
  assign t[142] = (t[185] & ~t[186]);
  assign t[143] = (t[187] & ~t[188]);
  assign t[144] = (t[189] & ~t[190]);
  assign t[145] = (t[191] & ~t[192]);
  assign t[146] = (t[193] & ~t[194]);
  assign t[147] = (t[195] & ~t[196]);
  assign t[148] = (t[197] & ~t[198]);
  assign t[149] = (t[199] & ~t[200]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (t[201] & ~t[202]);
  assign t[151] = (t[203] & ~t[204]);
  assign t[152] = (t[205] & ~t[206]);
  assign t[153] = (t[207] & ~t[208]);
  assign t[154] = (t[209] & ~t[210]);
  assign t[155] = (t[211] & ~t[212]);
  assign t[156] = (t[213] & ~t[214]);
  assign t[157] = t[215] ^ x[2];
  assign t[158] = t[216] ^ x[1];
  assign t[159] = t[217] ^ x[10];
  assign t[15] = ~(t[71] & t[72]);
  assign t[160] = t[218] ^ x[9];
  assign t[161] = t[219] ^ x[13];
  assign t[162] = t[220] ^ x[12];
  assign t[163] = t[221] ^ x[16];
  assign t[164] = t[222] ^ x[15];
  assign t[165] = t[223] ^ x[19];
  assign t[166] = t[224] ^ x[18];
  assign t[167] = t[225] ^ x[22];
  assign t[168] = t[226] ^ x[21];
  assign t[169] = t[227] ^ x[27];
  assign t[16] = ~(t[73] & t[74]);
  assign t[170] = t[228] ^ x[26];
  assign t[171] = t[229] ^ x[30];
  assign t[172] = t[230] ^ x[29];
  assign t[173] = t[231] ^ x[33];
  assign t[174] = t[232] ^ x[32];
  assign t[175] = t[233] ^ x[36];
  assign t[176] = t[234] ^ x[35];
  assign t[177] = t[235] ^ x[41];
  assign t[178] = t[236] ^ x[40];
  assign t[179] = t[237] ^ x[46];
  assign t[17] = ~(t[22]);
  assign t[180] = t[238] ^ x[45];
  assign t[181] = t[239] ^ x[49];
  assign t[182] = t[240] ^ x[48];
  assign t[183] = t[241] ^ x[52];
  assign t[184] = t[242] ^ x[51];
  assign t[185] = t[243] ^ x[55];
  assign t[186] = t[244] ^ x[54];
  assign t[187] = t[245] ^ x[58];
  assign t[188] = t[246] ^ x[57];
  assign t[189] = t[247] ^ x[61];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[248] ^ x[60];
  assign t[191] = t[249] ^ x[64];
  assign t[192] = t[250] ^ x[63];
  assign t[193] = t[251] ^ x[67];
  assign t[194] = t[252] ^ x[66];
  assign t[195] = t[253] ^ x[70];
  assign t[196] = t[254] ^ x[69];
  assign t[197] = t[255] ^ x[73];
  assign t[198] = t[256] ^ x[72];
  assign t[199] = t[257] ^ x[76];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[258] ^ x[75];
  assign t[201] = t[259] ^ x[79];
  assign t[202] = t[260] ^ x[78];
  assign t[203] = t[261] ^ x[82];
  assign t[204] = t[262] ^ x[81];
  assign t[205] = t[263] ^ x[85];
  assign t[206] = t[264] ^ x[84];
  assign t[207] = t[265] ^ x[88];
  assign t[208] = t[266] ^ x[87];
  assign t[209] = t[267] ^ x[91];
  assign t[20] = x[4] ? t[28] : t[27];
  assign t[210] = t[268] ^ x[90];
  assign t[211] = t[269] ^ x[94];
  assign t[212] = t[270] ^ x[93];
  assign t[213] = t[271] ^ x[97];
  assign t[214] = t[272] ^ x[96];
  assign t[215] = (x[0]);
  assign t[216] = (x[0]);
  assign t[217] = (x[8]);
  assign t[218] = (x[8]);
  assign t[219] = (x[11]);
  assign t[21] = x[4] ? t[30] : t[29];
  assign t[220] = (x[11]);
  assign t[221] = (x[14]);
  assign t[222] = (x[14]);
  assign t[223] = (x[17]);
  assign t[224] = (x[17]);
  assign t[225] = (x[20]);
  assign t[226] = (x[20]);
  assign t[227] = (x[25]);
  assign t[228] = (x[25]);
  assign t[229] = (x[28]);
  assign t[22] = ~(t[73]);
  assign t[230] = (x[28]);
  assign t[231] = (x[31]);
  assign t[232] = (x[31]);
  assign t[233] = (x[34]);
  assign t[234] = (x[34]);
  assign t[235] = (x[39]);
  assign t[236] = (x[39]);
  assign t[237] = (x[44]);
  assign t[238] = (x[44]);
  assign t[239] = (x[47]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[47]);
  assign t[241] = (x[50]);
  assign t[242] = (x[50]);
  assign t[243] = (x[53]);
  assign t[244] = (x[53]);
  assign t[245] = (x[56]);
  assign t[246] = (x[56]);
  assign t[247] = (x[59]);
  assign t[248] = (x[59]);
  assign t[249] = (x[62]);
  assign t[24] = t[33] | t[75];
  assign t[250] = (x[62]);
  assign t[251] = (x[65]);
  assign t[252] = (x[65]);
  assign t[253] = (x[68]);
  assign t[254] = (x[68]);
  assign t[255] = (x[71]);
  assign t[256] = (x[71]);
  assign t[257] = (x[74]);
  assign t[258] = (x[74]);
  assign t[259] = (x[77]);
  assign t[25] = t[17] ? x[24] : x[23];
  assign t[260] = (x[77]);
  assign t[261] = (x[80]);
  assign t[262] = (x[80]);
  assign t[263] = (x[83]);
  assign t[264] = (x[83]);
  assign t[265] = (x[86]);
  assign t[266] = (x[86]);
  assign t[267] = (x[89]);
  assign t[268] = (x[89]);
  assign t[269] = (x[92]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[270] = (x[92]);
  assign t[271] = (x[95]);
  assign t[272] = (x[95]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[3] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[76]);
  assign t[32] = ~(t[77]);
  assign t[33] = ~(t[44] | t[31]);
  assign t[34] = ~(t[45] & t[46]);
  assign t[35] = t[47] | t[78];
  assign t[36] = ~(t[48] & t[49]);
  assign t[37] = t[50] | t[79];
  assign t[38] = t[51] ? x[38] : x[37];
  assign t[39] = ~(t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[80];
  assign t[42] = t[17] ? x[43] : x[42];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[83]);
  assign t[47] = ~(t[59] | t[45]);
  assign t[48] = ~(t[84]);
  assign t[49] = ~(t[85]);
  assign t[4] = x[4] ? t[8] : t[7];
  assign t[50] = ~(t[60] | t[48]);
  assign t[51] = ~(t[22]);
  assign t[52] = ~(t[61] & t[62]);
  assign t[53] = t[63] | t[86];
  assign t[54] = ~(t[87]);
  assign t[55] = ~(t[88]);
  assign t[56] = ~(t[64] | t[54]);
  assign t[57] = ~(t[65] & t[66]);
  assign t[58] = t[67] | t[89];
  assign t[59] = ~(t[90]);
  assign t[5] = t[9] ^ x[5];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[92]);
  assign t[62] = ~(t[93]);
  assign t[63] = ~(t[68] | t[61]);
  assign t[64] = ~(t[94]);
  assign t[65] = ~(t[95]);
  assign t[66] = ~(t[96]);
  assign t[67] = ~(t[69] | t[65]);
  assign t[68] = ~(t[97]);
  assign t[69] = ~(t[98]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = t[128] ^ x[2];
  assign t[9] = x[6] ^ x[7];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [400:0] x;
 output [267:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[5], x[4], x[3], x[8], x[7], x[6], x[15]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[5], x[4], x[3], x[8], x[7], x[6], x[15]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[5], x[4], x[3], x[15]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[5], x[4], x[3], x[15]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[14], x[13], x[12], x[15]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[14], x[13], x[12], x[15]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[15]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[15]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[26], x[25], x[24], x[29], x[28], x[27], x[23], x[22], x[21], x[31], x[30]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[26], x[25], x[24], x[29], x[28], x[27], x[23], x[22], x[21], x[31], x[30]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[23], x[22], x[21], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[33], x[32]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[23], x[22], x[21], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[33], x[32]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[23], x[22], x[21], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[35], x[34]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[23], x[22], x[21], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[35], x[34]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[46], x[45], x[44], x[49], x[48], x[47], x[43], x[42], x[41], x[51], x[50]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[46], x[45], x[44], x[49], x[48], x[47], x[43], x[42], x[41], x[51], x[50]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[43], x[42], x[41], x[49], x[48], x[47], x[46], x[45], x[44], x[40], x[39], x[38], x[53], x[52]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[43], x[42], x[41], x[49], x[48], x[47], x[46], x[45], x[44], x[40], x[39], x[38], x[53], x[52]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[43], x[42], x[41], x[49], x[48], x[47], x[46], x[45], x[44], x[40], x[39], x[38], x[55], x[54]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[43], x[42], x[41], x[49], x[48], x[47], x[46], x[45], x[44], x[40], x[39], x[38], x[55], x[54]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[66], x[65], x[64], x[69], x[68], x[67], x[63], x[62], x[61], x[71], x[70]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[66], x[65], x[64], x[69], x[68], x[67], x[63], x[62], x[61], x[71], x[70]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[60], x[59], x[58], x[73], x[72]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[60], x[59], x[58], x[73], x[72]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[60], x[59], x[58], x[75], x[74]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[60], x[59], x[58], x[75], x[74]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[86], x[85], x[84], x[89], x[88], x[87], x[83], x[82], x[81], x[91], x[90]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[86], x[85], x[84], x[89], x[88], x[87], x[83], x[82], x[81], x[91], x[90]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[83], x[82], x[81], x[89], x[88], x[87], x[86], x[85], x[84], x[80], x[79], x[78], x[93], x[92]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[83], x[82], x[81], x[89], x[88], x[87], x[86], x[85], x[84], x[80], x[79], x[78], x[93], x[92]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[83], x[82], x[81], x[89], x[88], x[87], x[86], x[85], x[84], x[80], x[79], x[78], x[95], x[94]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[83], x[82], x[81], x[89], x[88], x[87], x[86], x[85], x[84], x[80], x[79], x[78], x[95], x[94]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[106], x[105], x[104], x[109], x[108], x[107], x[103], x[102], x[101], x[111], x[110]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[106], x[105], x[104], x[109], x[108], x[107], x[103], x[102], x[101], x[111], x[110]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[103], x[102], x[101], x[109], x[108], x[107], x[106], x[105], x[104], x[100], x[99], x[98], x[113], x[112]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[103], x[102], x[101], x[109], x[108], x[107], x[106], x[105], x[104], x[100], x[99], x[98], x[113], x[112]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[103], x[102], x[101], x[109], x[108], x[107], x[106], x[105], x[104], x[100], x[99], x[98], x[115], x[114]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[103], x[102], x[101], x[109], x[108], x[107], x[106], x[105], x[104], x[100], x[99], x[98], x[115], x[114]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[126], x[125], x[124], x[129], x[128], x[127], x[123], x[122], x[121], x[131], x[130]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[126], x[125], x[124], x[129], x[128], x[127], x[123], x[122], x[121], x[131], x[130]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[123], x[122], x[121], x[129], x[128], x[127], x[126], x[125], x[124], x[120], x[119], x[118], x[133], x[132]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[123], x[122], x[121], x[129], x[128], x[127], x[126], x[125], x[124], x[120], x[119], x[118], x[133], x[132]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[123], x[122], x[121], x[129], x[128], x[127], x[126], x[125], x[124], x[120], x[119], x[118], x[135], x[134]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[123], x[122], x[121], x[129], x[128], x[127], x[126], x[125], x[124], x[120], x[119], x[118], x[135], x[134]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[146], x[145], x[144], x[149], x[148], x[147], x[143], x[142], x[141], x[151], x[150]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[146], x[145], x[144], x[149], x[148], x[147], x[143], x[142], x[141], x[151], x[150]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[143], x[142], x[141], x[149], x[148], x[147], x[146], x[145], x[144], x[140], x[139], x[138], x[153], x[152]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[143], x[142], x[141], x[149], x[148], x[147], x[146], x[145], x[144], x[140], x[139], x[138], x[153], x[152]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[143], x[142], x[141], x[149], x[148], x[147], x[146], x[145], x[144], x[140], x[139], x[138], x[155], x[154]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[143], x[142], x[141], x[149], x[148], x[147], x[146], x[145], x[144], x[140], x[139], x[138], x[155], x[154]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[166], x[165], x[164], x[169], x[168], x[167], x[163], x[162], x[161], x[171], x[170]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[166], x[165], x[164], x[169], x[168], x[167], x[163], x[162], x[161], x[171], x[170]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[163], x[162], x[161], x[169], x[168], x[167], x[166], x[165], x[164], x[160], x[159], x[158], x[173], x[172]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[163], x[162], x[161], x[169], x[168], x[167], x[166], x[165], x[164], x[160], x[159], x[158], x[173], x[172]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[163], x[162], x[161], x[169], x[168], x[167], x[166], x[165], x[164], x[160], x[159], x[158], x[175], x[174]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[163], x[162], x[161], x[169], x[168], x[167], x[166], x[165], x[164], x[160], x[159], x[158], x[175], x[174]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[186], x[185], x[184], x[189], x[188], x[187], x[183], x[182], x[181], x[191], x[190]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[186], x[185], x[184], x[189], x[188], x[187], x[183], x[182], x[181], x[191], x[190]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[193], x[192]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[193], x[192]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[195], x[194]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[195], x[194]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[206], x[205], x[204], x[209], x[208], x[207], x[203], x[202], x[201], x[211], x[210]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[206], x[205], x[204], x[209], x[208], x[207], x[203], x[202], x[201], x[211], x[210]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[203], x[202], x[201], x[209], x[208], x[207], x[206], x[205], x[204], x[200], x[199], x[198], x[213], x[212]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[203], x[202], x[201], x[209], x[208], x[207], x[206], x[205], x[204], x[200], x[199], x[198], x[213], x[212]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[203], x[202], x[201], x[209], x[208], x[207], x[206], x[205], x[204], x[200], x[199], x[198], x[215], x[214]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[203], x[202], x[201], x[209], x[208], x[207], x[206], x[205], x[204], x[200], x[199], x[198], x[215], x[214]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[226], x[225], x[224], x[229], x[228], x[227], x[223], x[222], x[221], x[231], x[230]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[226], x[225], x[224], x[229], x[228], x[227], x[223], x[222], x[221], x[231], x[230]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[223], x[222], x[221], x[229], x[228], x[227], x[226], x[225], x[224], x[220], x[219], x[218], x[233], x[232]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[223], x[222], x[221], x[229], x[228], x[227], x[226], x[225], x[224], x[220], x[219], x[218], x[233], x[232]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[223], x[222], x[221], x[229], x[228], x[227], x[226], x[225], x[224], x[220], x[219], x[218], x[235], x[234]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[223], x[222], x[221], x[229], x[228], x[227], x[226], x[225], x[224], x[220], x[219], x[218], x[235], x[234]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[246], x[245], x[244], x[249], x[248], x[247], x[243], x[242], x[241], x[251], x[250]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[246], x[245], x[244], x[249], x[248], x[247], x[243], x[242], x[241], x[251], x[250]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[243], x[242], x[241], x[249], x[248], x[247], x[246], x[245], x[244], x[240], x[239], x[238], x[253], x[252]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[243], x[242], x[241], x[249], x[248], x[247], x[246], x[245], x[244], x[240], x[239], x[238], x[253], x[252]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[243], x[242], x[241], x[249], x[248], x[247], x[246], x[245], x[244], x[240], x[239], x[238], x[255], x[254]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[243], x[242], x[241], x[249], x[248], x[247], x[246], x[245], x[244], x[240], x[239], x[238], x[255], x[254]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[266], x[265], x[264], x[269], x[268], x[267], x[263], x[262], x[261], x[271], x[270]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[266], x[265], x[264], x[269], x[268], x[267], x[263], x[262], x[261], x[271], x[270]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[263], x[262], x[261], x[269], x[268], x[267], x[266], x[265], x[264], x[260], x[259], x[258], x[273], x[272]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[263], x[262], x[261], x[269], x[268], x[267], x[266], x[265], x[264], x[260], x[259], x[258], x[273], x[272]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[263], x[262], x[261], x[269], x[268], x[267], x[266], x[265], x[264], x[260], x[259], x[258], x[275], x[274]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[263], x[262], x[261], x[269], x[268], x[267], x[266], x[265], x[264], x[260], x[259], x[258], x[275], x[274]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[286], x[285], x[284], x[289], x[288], x[287], x[283], x[282], x[281], x[291], x[290]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[286], x[285], x[284], x[289], x[288], x[287], x[283], x[282], x[281], x[291], x[290]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[283], x[282], x[281], x[289], x[288], x[287], x[286], x[285], x[284], x[280], x[279], x[278], x[293], x[292]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[283], x[282], x[281], x[289], x[288], x[287], x[286], x[285], x[284], x[280], x[279], x[278], x[293], x[292]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[283], x[282], x[281], x[289], x[288], x[287], x[286], x[285], x[284], x[280], x[279], x[278], x[295], x[294]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[283], x[282], x[281], x[289], x[288], x[287], x[286], x[285], x[284], x[280], x[279], x[278], x[295], x[294]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[306], x[305], x[304], x[309], x[308], x[307], x[303], x[302], x[301], x[311], x[310]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[306], x[305], x[304], x[309], x[308], x[307], x[303], x[302], x[301], x[311], x[310]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[303], x[302], x[301], x[309], x[308], x[307], x[306], x[305], x[304], x[300], x[299], x[298], x[313], x[312]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[303], x[302], x[301], x[309], x[308], x[307], x[306], x[305], x[304], x[300], x[299], x[298], x[313], x[312]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[303], x[302], x[301], x[309], x[308], x[307], x[306], x[305], x[304], x[300], x[299], x[298], x[315], x[314]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[303], x[302], x[301], x[309], x[308], x[307], x[306], x[305], x[304], x[300], x[299], x[298], x[315], x[314]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[326], x[325], x[324], x[329], x[328], x[327], x[323], x[322], x[321], x[331], x[330]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[326], x[325], x[324], x[329], x[328], x[327], x[323], x[322], x[321], x[331], x[330]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[323], x[322], x[321], x[329], x[328], x[327], x[326], x[325], x[324], x[320], x[319], x[318], x[333], x[332]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[323], x[322], x[321], x[329], x[328], x[327], x[326], x[325], x[324], x[320], x[319], x[318], x[333], x[332]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[323], x[322], x[321], x[329], x[328], x[327], x[326], x[325], x[324], x[320], x[319], x[318], x[335], x[334]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[323], x[322], x[321], x[329], x[328], x[327], x[326], x[325], x[324], x[320], x[319], x[318], x[335], x[334]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[89], x[88], x[87], x[309], x[308], x[307], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[49], x[48], x[47], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[229], x[228], x[227], x[60], x[59], x[58], x[180], x[179], x[178], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[120], x[119], x[118], x[320], x[319], x[318], x[277], x[276], x[226], x[225], x[224], x[223], x[222], x[221], x[280], x[279], x[278], x[220], x[219], x[218], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[17], x[16], x[337], x[336], x[15], x[29], x[28], x[27]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[89], x[88], x[87], x[309], x[308], x[307], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[49], x[48], x[47], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[229], x[228], x[227], x[60], x[59], x[58], x[180], x[179], x[178], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[120], x[119], x[118], x[320], x[319], x[318], x[277], x[276], x[226], x[225], x[224], x[223], x[222], x[221], x[280], x[279], x[278], x[220], x[219], x[218], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[17], x[16], x[337], x[336], x[15], x[29], x[28], x[27]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[86], x[85], x[84], x[306], x[305], x[304], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[46], x[45], x[44], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[226], x[225], x[224], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[338], x[336], x[15], x[20], x[19], x[18]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[86], x[85], x[84], x[306], x[305], x[304], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[46], x[45], x[44], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[226], x[225], x[224], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[338], x[336], x[15], x[20], x[19], x[18]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[83], x[82], x[81], x[303], x[302], x[301], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[43], x[42], x[41], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[223], x[222], x[221], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[229], x[228], x[227], x[226], x[225], x[224], x[52], x[53], x[280], x[279], x[278], x[293], x[292], x[220], x[219], x[218], x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[33], x[32], x[339], x[336], x[15], x[23], x[22], x[21]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[83], x[82], x[81], x[303], x[302], x[301], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[43], x[42], x[41], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[223], x[222], x[221], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[229], x[228], x[227], x[226], x[225], x[224], x[52], x[53], x[280], x[279], x[278], x[293], x[292], x[220], x[219], x[218], x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[33], x[32], x[339], x[336], x[15], x[23], x[22], x[21]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[83], x[82], x[81], x[303], x[302], x[301], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[43], x[42], x[41], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[223], x[222], x[221], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[229], x[228], x[227], x[226], x[225], x[224], x[55], x[54], x[280], x[279], x[278], x[295], x[294], x[220], x[219], x[218], x[35], x[34], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[340], x[336], x[15], x[26], x[25], x[24]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[83], x[82], x[81], x[303], x[302], x[301], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[43], x[42], x[41], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[223], x[222], x[221], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[229], x[228], x[227], x[226], x[225], x[224], x[55], x[54], x[280], x[279], x[278], x[295], x[294], x[220], x[219], x[218], x[35], x[34], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[340], x[336], x[15], x[26], x[25], x[24]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[89], x[88], x[87], x[209], x[208], x[207], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[29], x[28], x[27], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[229], x[228], x[227], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[176], x[177], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[60], x[59], x[58], x[180], x[179], x[178], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[300], x[299], x[298], x[100], x[99], x[98], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[160], x[159], x[158], x[240], x[239], x[238], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[37], x[36], x[341], x[336], x[15], x[49], x[48], x[47]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[89], x[88], x[87], x[209], x[208], x[207], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[29], x[28], x[27], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[229], x[228], x[227], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[176], x[177], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[60], x[59], x[58], x[180], x[179], x[178], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[300], x[299], x[298], x[100], x[99], x[98], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[160], x[159], x[158], x[240], x[239], x[238], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[37], x[36], x[341], x[336], x[15], x[49], x[48], x[47]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[86], x[85], x[84], x[206], x[205], x[204], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[26], x[25], x[24], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[306], x[305], x[304], x[226], x[225], x[224], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[51], x[50], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[342], x[336], x[15], x[40], x[39], x[38]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[86], x[85], x[84], x[206], x[205], x[204], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[26], x[25], x[24], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[306], x[305], x[304], x[226], x[225], x[224], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[51], x[50], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[342], x[336], x[15], x[40], x[39], x[38]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[83], x[82], x[81], x[203], x[202], x[201], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[23], x[22], x[21], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[303], x[302], x[301], x[223], x[222], x[221], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[309], x[308], x[307], x[306], x[305], x[304], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[32], x[33], x[160], x[159], x[158], x[233], x[232], x[240], x[239], x[238], x[53], x[52], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[343], x[336], x[15], x[43], x[42], x[41]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[83], x[82], x[81], x[203], x[202], x[201], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[23], x[22], x[21], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[303], x[302], x[301], x[223], x[222], x[221], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[309], x[308], x[307], x[306], x[305], x[304], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[32], x[33], x[160], x[159], x[158], x[233], x[232], x[240], x[239], x[238], x[53], x[52], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[343], x[336], x[15], x[43], x[42], x[41]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[83], x[82], x[81], x[203], x[202], x[201], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[23], x[22], x[21], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[303], x[302], x[301], x[223], x[222], x[221], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[309], x[308], x[307], x[306], x[305], x[304], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[34], x[35], x[160], x[159], x[158], x[235], x[234], x[240], x[239], x[238], x[55], x[54], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[344], x[336], x[15], x[46], x[45], x[44]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[83], x[82], x[81], x[203], x[202], x[201], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[23], x[22], x[21], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[303], x[302], x[301], x[223], x[222], x[221], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[309], x[308], x[307], x[306], x[305], x[304], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[34], x[35], x[160], x[159], x[158], x[235], x[234], x[240], x[239], x[238], x[55], x[54], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[344], x[336], x[15], x[46], x[45], x[44]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[29], x[28], x[27], x[49], x[48], x[47], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[89], x[88], x[87], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[160], x[159], x[158], x[280], x[279], x[278], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[57], x[56], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[345], x[336], x[15], x[69], x[68], x[67]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[29], x[28], x[27], x[49], x[48], x[47], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[89], x[88], x[87], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[160], x[159], x[158], x[280], x[279], x[278], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[57], x[56], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[345], x[336], x[15], x[69], x[68], x[67]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[46], x[45], x[44], x[26], x[25], x[24], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[86], x[85], x[84], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[346], x[336], x[15], x[60], x[59], x[58]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[46], x[45], x[44], x[26], x[25], x[24], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[86], x[85], x[84], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[346], x[336], x[15], x[60], x[59], x[58]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[83], x[82], x[81], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[92], x[93], x[180], x[179], x[178], x[73], x[72], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[347], x[336], x[15], x[63], x[62], x[61]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[83], x[82], x[81], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[92], x[93], x[180], x[179], x[178], x[73], x[72], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[347], x[336], x[15], x[63], x[62], x[61]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[83], x[82], x[81], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[94], x[95], x[180], x[179], x[178], x[75], x[74], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[348], x[336], x[15], x[66], x[65], x[64]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[83], x[82], x[81], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[94], x[95], x[180], x[179], x[178], x[75], x[74], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[348], x[336], x[15], x[66], x[65], x[64]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[29], x[28], x[27], x[49], x[48], x[47], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[269], x[268], x[267], x[149], x[148], x[147], x[109], x[108], x[107], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[69], x[68], x[67], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[146], x[145], x[144], x[143], x[142], x[141], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[160], x[159], x[158], x[280], x[279], x[278], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[260], x[259], x[258], x[140], x[139], x[138], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[60], x[59], x[58], x[200], x[199], x[198], x[77], x[76], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[349], x[336], x[15], x[89], x[88], x[87]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[29], x[28], x[27], x[49], x[48], x[47], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[269], x[268], x[267], x[149], x[148], x[147], x[109], x[108], x[107], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[69], x[68], x[67], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[146], x[145], x[144], x[143], x[142], x[141], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[160], x[159], x[158], x[280], x[279], x[278], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[260], x[259], x[258], x[140], x[139], x[138], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[60], x[59], x[58], x[200], x[199], x[198], x[77], x[76], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[349], x[336], x[15], x[89], x[88], x[87]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[46], x[45], x[44], x[26], x[25], x[24], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[146], x[145], x[144], x[266], x[265], x[264], x[106], x[105], x[104], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[66], x[65], x[64], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[91], x[90], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[350], x[336], x[15], x[80], x[79], x[78]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[46], x[45], x[44], x[26], x[25], x[24], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[146], x[145], x[144], x[266], x[265], x[264], x[106], x[105], x[104], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[66], x[65], x[64], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[91], x[90], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[350], x[336], x[15], x[80], x[79], x[78]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[263], x[262], x[261], x[143], x[142], x[141], x[103], x[102], x[101], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[269], x[268], x[267], x[266], x[265], x[264], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[72], x[73], x[60], x[59], x[58], x[112], x[113], x[200], x[199], x[198], x[93], x[92], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[351], x[336], x[15], x[83], x[82], x[81]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[263], x[262], x[261], x[143], x[142], x[141], x[103], x[102], x[101], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[269], x[268], x[267], x[266], x[265], x[264], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[72], x[73], x[60], x[59], x[58], x[112], x[113], x[200], x[199], x[198], x[93], x[92], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[351], x[336], x[15], x[83], x[82], x[81]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[263], x[262], x[261], x[143], x[142], x[141], x[103], x[102], x[101], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[269], x[268], x[267], x[266], x[265], x[264], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[74], x[75], x[60], x[59], x[58], x[114], x[115], x[200], x[199], x[198], x[95], x[94], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[352], x[336], x[15], x[86], x[85], x[84]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[43], x[42], x[41], x[23], x[22], x[21], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[263], x[262], x[261], x[143], x[142], x[141], x[103], x[102], x[101], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[269], x[268], x[267], x[266], x[265], x[264], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[74], x[75], x[60], x[59], x[58], x[114], x[115], x[200], x[199], x[198], x[95], x[94], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[352], x[336], x[15], x[86], x[85], x[84]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[169], x[168], x[167], x[229], x[228], x[227], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[129], x[128], x[127], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[189], x[188], x[187], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[260], x[259], x[258], x[140], x[139], x[138], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[240], x[239], x[238], x[40], x[39], x[38], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[80], x[79], x[78], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[97], x[96], x[353], x[336], x[15], x[109], x[108], x[107]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[169], x[168], x[167], x[229], x[228], x[227], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[129], x[128], x[127], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[189], x[188], x[187], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[260], x[259], x[258], x[140], x[139], x[138], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[240], x[239], x[238], x[40], x[39], x[38], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[80], x[79], x[78], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[97], x[96], x[353], x[336], x[15], x[109], x[108], x[107]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[166], x[165], x[164], x[226], x[225], x[224], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[126], x[125], x[124], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[186], x[185], x[184], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[111], x[110], x[354], x[336], x[15], x[100], x[99], x[98]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[166], x[165], x[164], x[226], x[225], x[224], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[126], x[125], x[124], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[186], x[185], x[184], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[111], x[110], x[354], x[336], x[15], x[100], x[99], x[98]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[163], x[162], x[161], x[223], x[222], x[221], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[132], x[133], x[80], x[79], x[78], x[192], x[193], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[113], x[112], x[355], x[336], x[15], x[103], x[102], x[101]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[163], x[162], x[161], x[223], x[222], x[221], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[132], x[133], x[80], x[79], x[78], x[192], x[193], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[113], x[112], x[355], x[336], x[15], x[103], x[102], x[101]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[163], x[162], x[161], x[223], x[222], x[221], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[134], x[135], x[80], x[79], x[78], x[194], x[195], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[115], x[114], x[356], x[336], x[15], x[106], x[105], x[104]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[163], x[162], x[161], x[223], x[222], x[221], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[134], x[135], x[80], x[79], x[78], x[194], x[195], x[300], x[299], x[298], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[115], x[114], x[356], x[336], x[15], x[106], x[105], x[104]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[169], x[168], x[167], x[289], x[288], x[287], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[109], x[108], x[107], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[257], x[256], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[329], x[328], x[327], x[260], x[259], x[258], x[140], x[139], x[138], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[20], x[19], x[18], x[220], x[219], x[218], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[200], x[199], x[198], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[117], x[116], x[357], x[336], x[15], x[129], x[128], x[127]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[169], x[168], x[167], x[289], x[288], x[287], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[109], x[108], x[107], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[257], x[256], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[329], x[328], x[327], x[260], x[259], x[258], x[140], x[139], x[138], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[20], x[19], x[18], x[220], x[219], x[218], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[200], x[199], x[198], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[117], x[116], x[357], x[336], x[15], x[129], x[128], x[127]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[166], x[165], x[164], x[286], x[285], x[284], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[106], x[105], x[104], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[26], x[25], x[24], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[326], x[325], x[324], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[131], x[130], x[358], x[336], x[15], x[120], x[119], x[118]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[166], x[165], x[164], x[286], x[285], x[284], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[106], x[105], x[104], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[26], x[25], x[24], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[326], x[325], x[324], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[131], x[130], x[358], x[336], x[15], x[120], x[119], x[118]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[163], x[162], x[161], x[283], x[282], x[281], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[23], x[22], x[21], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[112], x[113], x[200], x[199], x[198], x[333], x[332], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[133], x[132], x[359], x[336], x[15], x[123], x[122], x[121]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[163], x[162], x[161], x[283], x[282], x[281], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[23], x[22], x[21], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[112], x[113], x[200], x[199], x[198], x[333], x[332], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[133], x[132], x[359], x[336], x[15], x[123], x[122], x[121]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[163], x[162], x[161], x[283], x[282], x[281], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[23], x[22], x[21], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[114], x[115], x[200], x[199], x[198], x[335], x[334], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[135], x[134], x[360], x[336], x[15], x[126], x[125], x[124]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[163], x[162], x[161], x[283], x[282], x[281], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[23], x[22], x[21], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[114], x[115], x[200], x[199], x[198], x[335], x[334], x[320], x[319], x[318], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[135], x[134], x[360], x[336], x[15], x[126], x[125], x[124]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[109], x[108], x[107], x[129], x[128], x[127], x[169], x[168], x[167], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[166], x[165], x[164], x[163], x[162], x[161], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[269], x[268], x[267], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[200], x[199], x[198], x[80], x[79], x[78], x[266], x[265], x[264], x[263], x[262], x[261], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[137], x[136], x[361], x[336], x[15], x[149], x[148], x[147]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[109], x[108], x[107], x[129], x[128], x[127], x[169], x[168], x[167], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[166], x[165], x[164], x[163], x[162], x[161], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[269], x[268], x[267], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[200], x[199], x[198], x[80], x[79], x[78], x[266], x[265], x[264], x[263], x[262], x[261], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[137], x[136], x[361], x[336], x[15], x[149], x[148], x[147]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[126], x[125], x[124], x[106], x[105], x[104], x[166], x[165], x[164], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[266], x[265], x[264], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[269], x[268], x[267], x[263], x[262], x[261], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[151], x[150], x[362], x[336], x[15], x[140], x[139], x[138]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[126], x[125], x[124], x[106], x[105], x[104], x[166], x[165], x[164], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[266], x[265], x[264], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[269], x[268], x[267], x[263], x[262], x[261], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[151], x[150], x[362], x[336], x[15], x[140], x[139], x[138]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[163], x[162], x[161], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[169], x[168], x[167], x[166], x[165], x[164], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[263], x[262], x[261], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[269], x[268], x[267], x[266], x[265], x[264], x[172], x[173], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[153], x[152], x[363], x[336], x[15], x[143], x[142], x[141]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[163], x[162], x[161], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[169], x[168], x[167], x[166], x[165], x[164], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[263], x[262], x[261], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[269], x[268], x[267], x[266], x[265], x[264], x[172], x[173], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[8], x[7], x[6], x[5], x[4], x[3], x[11], x[10], x[9], x[153], x[152], x[363], x[336], x[15], x[143], x[142], x[141]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[163], x[162], x[161], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[263], x[262], x[261], x[160], x[159], x[158], x[149], x[148], x[147], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[269], x[268], x[267], x[266], x[265], x[264], x[174], x[175], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[155], x[154], x[364], x[336], x[15], x[146], x[145], x[144]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[163], x[162], x[161], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[263], x[262], x[261], x[160], x[159], x[158], x[149], x[148], x[147], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[269], x[268], x[267], x[266], x[265], x[264], x[174], x[175], x[140], x[139], x[138], x[260], x[259], x[258], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[155], x[154], x[364], x[336], x[15], x[146], x[145], x[144]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[109], x[108], x[107], x[129], x[128], x[127], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[149], x[148], x[147], x[69], x[68], x[67], x[189], x[188], x[187], x[49], x[48], x[47], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[146], x[145], x[144], x[143], x[142], x[141], x[269], x[268], x[267], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[186], x[185], x[184], x[183], x[182], x[181], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[200], x[199], x[198], x[80], x[79], x[78], x[136], x[137], x[140], x[139], x[138], x[266], x[265], x[264], x[263], x[262], x[261], x[60], x[59], x[58], x[180], x[179], x[178], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[260], x[259], x[258], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[157], x[156], x[365], x[336], x[15], x[169], x[168], x[167]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[109], x[108], x[107], x[129], x[128], x[127], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[149], x[148], x[147], x[69], x[68], x[67], x[189], x[188], x[187], x[49], x[48], x[47], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[146], x[145], x[144], x[143], x[142], x[141], x[269], x[268], x[267], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[186], x[185], x[184], x[183], x[182], x[181], x[46], x[45], x[44], x[43], x[42], x[41], x[289], x[288], x[287], x[200], x[199], x[198], x[80], x[79], x[78], x[136], x[137], x[140], x[139], x[138], x[266], x[265], x[264], x[263], x[262], x[261], x[60], x[59], x[58], x[180], x[179], x[178], x[36], x[37], x[40], x[39], x[38], x[286], x[285], x[284], x[283], x[282], x[281], x[260], x[259], x[258], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[157], x[156], x[365], x[336], x[15], x[169], x[168], x[167]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[126], x[125], x[124], x[106], x[105], x[104], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[146], x[145], x[144], x[186], x[185], x[184], x[66], x[65], x[64], x[46], x[45], x[44], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[149], x[148], x[147], x[143], x[142], x[141], x[266], x[265], x[264], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[171], x[170], x[366], x[336], x[15], x[160], x[159], x[158]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[126], x[125], x[124], x[106], x[105], x[104], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[146], x[145], x[144], x[186], x[185], x[184], x[66], x[65], x[64], x[46], x[45], x[44], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[149], x[148], x[147], x[143], x[142], x[141], x[266], x[265], x[264], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[49], x[48], x[47], x[43], x[42], x[41], x[286], x[285], x[284], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[171], x[170], x[366], x[336], x[15], x[160], x[159], x[158]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[143], x[142], x[141], x[63], x[62], x[61], x[183], x[182], x[181], x[43], x[42], x[41], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[149], x[148], x[147], x[146], x[145], x[144], x[263], x[262], x[261], x[69], x[68], x[67], x[66], x[65], x[64], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[140], x[139], x[138], x[269], x[268], x[267], x[266], x[265], x[264], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[152], x[153], x[260], x[259], x[258], x[52], x[53], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[173], x[172], x[367], x[336], x[15], x[163], x[162], x[161]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[143], x[142], x[141], x[63], x[62], x[61], x[183], x[182], x[181], x[43], x[42], x[41], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[149], x[148], x[147], x[146], x[145], x[144], x[263], x[262], x[261], x[69], x[68], x[67], x[66], x[65], x[64], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[140], x[139], x[138], x[269], x[268], x[267], x[266], x[265], x[264], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[152], x[153], x[260], x[259], x[258], x[52], x[53], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[173], x[172], x[367], x[336], x[15], x[163], x[162], x[161]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[143], x[142], x[141], x[63], x[62], x[61], x[183], x[182], x[181], x[43], x[42], x[41], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[149], x[148], x[147], x[146], x[145], x[144], x[263], x[262], x[261], x[69], x[68], x[67], x[66], x[65], x[64], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[140], x[139], x[138], x[269], x[268], x[267], x[266], x[265], x[264], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[154], x[155], x[260], x[259], x[258], x[55], x[54], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[175], x[174], x[368], x[336], x[15], x[166], x[165], x[164]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[123], x[122], x[121], x[103], x[102], x[101], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[143], x[142], x[141], x[63], x[62], x[61], x[183], x[182], x[181], x[43], x[42], x[41], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[149], x[148], x[147], x[146], x[145], x[144], x[263], x[262], x[261], x[69], x[68], x[67], x[66], x[65], x[64], x[189], x[188], x[187], x[186], x[185], x[184], x[49], x[48], x[47], x[46], x[45], x[44], x[283], x[282], x[281], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[140], x[139], x[138], x[269], x[268], x[267], x[266], x[265], x[264], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[40], x[39], x[38], x[289], x[288], x[287], x[286], x[285], x[284], x[154], x[155], x[260], x[259], x[258], x[55], x[54], x[280], x[279], x[278], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[175], x[174], x[368], x[336], x[15], x[166], x[165], x[164]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[229], x[228], x[227], x[29], x[28], x[27], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[209], x[208], x[207], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[289], x[288], x[287], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[286], x[285], x[284], x[283], x[282], x[281], x[69], x[68], x[67], x[240], x[239], x[238], x[40], x[39], x[38], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[160], x[159], x[158], x[280], x[279], x[278], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[100], x[99], x[98], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[177], x[176], x[369], x[336], x[15], x[189], x[188], x[187]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[229], x[228], x[227], x[29], x[28], x[27], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[209], x[208], x[207], x[26], x[25], x[24], x[23], x[22], x[21], x[169], x[168], x[167], x[289], x[288], x[287], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[16], x[17], x[20], x[19], x[18], x[166], x[165], x[164], x[163], x[162], x[161], x[36], x[37], x[286], x[285], x[284], x[283], x[282], x[281], x[69], x[68], x[67], x[240], x[239], x[238], x[40], x[39], x[38], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[160], x[159], x[158], x[280], x[279], x[278], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[100], x[99], x[98], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[177], x[176], x[369], x[336], x[15], x[189], x[188], x[187]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[226], x[225], x[224], x[26], x[25], x[24], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[206], x[205], x[204], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[66], x[65], x[64], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[191], x[190], x[370], x[336], x[15], x[180], x[179], x[178]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[226], x[225], x[224], x[26], x[25], x[24], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[206], x[205], x[204], x[286], x[285], x[284], x[29], x[28], x[27], x[23], x[22], x[21], x[166], x[165], x[164], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[50], x[51], x[289], x[288], x[287], x[283], x[282], x[281], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[66], x[65], x[64], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[191], x[190], x[370], x[336], x[15], x[180], x[179], x[178]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[223], x[222], x[221], x[23], x[22], x[21], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[213], x[212], x[100], x[99], x[98], x[72], x[73], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[193], x[192], x[371], x[336], x[15], x[183], x[182], x[181]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[223], x[222], x[221], x[23], x[22], x[21], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[52], x[53], x[280], x[279], x[278], x[32], x[33], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[213], x[212], x[100], x[99], x[98], x[72], x[73], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[193], x[192], x[371], x[336], x[15], x[183], x[182], x[181]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[223], x[222], x[221], x[23], x[22], x[21], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[215], x[214], x[100], x[99], x[98], x[74], x[75], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[195], x[194], x[372], x[336], x[15], x[186], x[185], x[184]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[223], x[222], x[221], x[23], x[22], x[21], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[283], x[282], x[281], x[29], x[28], x[27], x[26], x[25], x[24], x[163], x[162], x[161], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[289], x[288], x[287], x[286], x[285], x[284], x[20], x[19], x[18], x[169], x[168], x[167], x[166], x[165], x[164], x[63], x[62], x[61], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[55], x[54], x[280], x[279], x[278], x[34], x[35], x[160], x[159], x[158], x[69], x[68], x[67], x[66], x[65], x[64], x[215], x[214], x[100], x[99], x[98], x[74], x[75], x[60], x[59], x[58], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[195], x[194], x[372], x[336], x[15], x[186], x[185], x[184]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[229], x[228], x[227], x[169], x[168], x[167], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[189], x[188], x[187], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[129], x[128], x[127], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[240], x[239], x[238], x[40], x[39], x[38], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[260], x[259], x[258], x[140], x[139], x[138], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[300], x[299], x[298], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[197], x[196], x[373], x[336], x[15], x[209], x[208], x[207]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[229], x[228], x[227], x[169], x[168], x[167], x[226], x[225], x[224], x[223], x[222], x[221], x[249], x[248], x[247], x[49], x[48], x[47], x[189], x[188], x[187], x[269], x[268], x[267], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[129], x[128], x[127], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[136], x[137], x[266], x[265], x[264], x[263], x[262], x[261], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[126], x[125], x[124], x[123], x[122], x[121], x[89], x[88], x[87], x[240], x[239], x[238], x[40], x[39], x[38], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[260], x[259], x[258], x[140], x[139], x[138], x[116], x[117], x[120], x[119], x[118], x[86], x[85], x[84], x[83], x[82], x[81], x[300], x[299], x[298], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[197], x[196], x[373], x[336], x[15], x[209], x[208], x[207]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[226], x[225], x[224], x[166], x[165], x[164], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[186], x[185], x[184], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[126], x[125], x[124], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[211], x[210], x[374], x[336], x[15], x[200], x[199], x[198]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[226], x[225], x[224], x[166], x[165], x[164], x[46], x[45], x[44], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[186], x[185], x[184], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[266], x[265], x[264], x[126], x[125], x[124], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[150], x[151], x[269], x[268], x[267], x[263], x[262], x[261], x[129], x[128], x[127], x[123], x[122], x[121], x[86], x[85], x[84], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[211], x[210], x[374], x[336], x[15], x[200], x[199], x[198]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[223], x[222], x[221], x[163], x[162], x[161], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[192], x[193], x[300], x[299], x[298], x[132], x[133], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[213], x[212], x[375], x[336], x[15], x[203], x[202], x[201]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[223], x[222], x[221], x[163], x[162], x[161], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[152], x[153], x[260], x[259], x[258], x[172], x[173], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[192], x[193], x[300], x[299], x[298], x[132], x[133], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[213], x[212], x[375], x[336], x[15], x[203], x[202], x[201]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[223], x[222], x[221], x[163], x[162], x[161], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[194], x[195], x[300], x[299], x[298], x[134], x[135], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[215], x[214], x[376], x[336], x[15], x[206], x[205], x[204]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[223], x[222], x[221], x[163], x[162], x[161], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[43], x[42], x[41], x[183], x[182], x[181], x[263], x[262], x[261], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[123], x[122], x[121], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[269], x[268], x[267], x[266], x[265], x[264], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[129], x[128], x[127], x[126], x[125], x[124], x[83], x[82], x[81], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[154], x[155], x[260], x[259], x[258], x[174], x[175], x[140], x[139], x[138], x[120], x[119], x[118], x[89], x[88], x[87], x[86], x[85], x[84], x[194], x[195], x[300], x[299], x[298], x[134], x[135], x[80], x[79], x[78], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[215], x[214], x[376], x[336], x[15], x[206], x[205], x[204]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[189], x[188], x[187], x[209], x[208], x[207], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[249], x[248], x[247], x[129], x[128], x[127], x[329], x[328], x[327], x[269], x[268], x[267], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[246], x[245], x[244], x[243], x[242], x[241], x[49], x[48], x[47], x[297], x[296], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[300], x[299], x[298], x[100], x[99], x[98], x[237], x[236], x[240], x[239], x[238], x[46], x[45], x[44], x[43], x[42], x[41], x[120], x[119], x[118], x[320], x[319], x[318], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[40], x[39], x[38], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[217], x[216], x[377], x[336], x[15], x[229], x[228], x[227]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[189], x[188], x[187], x[209], x[208], x[207], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[249], x[248], x[247], x[129], x[128], x[127], x[329], x[328], x[327], x[269], x[268], x[267], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[246], x[245], x[244], x[243], x[242], x[241], x[49], x[48], x[47], x[297], x[296], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[300], x[299], x[298], x[100], x[99], x[98], x[237], x[236], x[240], x[239], x[238], x[46], x[45], x[44], x[43], x[42], x[41], x[120], x[119], x[118], x[320], x[319], x[318], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[40], x[39], x[38], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[217], x[216], x[377], x[336], x[15], x[229], x[228], x[227]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[206], x[205], x[204], x[186], x[185], x[184], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[246], x[245], x[244], x[326], x[325], x[324], x[126], x[125], x[124], x[266], x[265], x[264], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[249], x[248], x[247], x[243], x[242], x[241], x[46], x[45], x[44], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[231], x[230], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[378], x[336], x[15], x[220], x[219], x[218]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[206], x[205], x[204], x[186], x[185], x[184], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[246], x[245], x[244], x[326], x[325], x[324], x[126], x[125], x[124], x[266], x[265], x[264], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[249], x[248], x[247], x[243], x[242], x[241], x[46], x[45], x[44], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[231], x[230], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[378], x[336], x[15], x[220], x[219], x[218]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[243], x[242], x[241], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[249], x[248], x[247], x[246], x[245], x[244], x[43], x[42], x[41], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[240], x[239], x[238], x[49], x[48], x[47], x[46], x[45], x[44], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[253], x[252], x[40], x[39], x[38], x[273], x[272], x[20], x[19], x[18], x[233], x[232], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[379], x[336], x[15], x[223], x[222], x[221]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[243], x[242], x[241], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[249], x[248], x[247], x[246], x[245], x[244], x[43], x[42], x[41], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[240], x[239], x[238], x[49], x[48], x[47], x[46], x[45], x[44], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[253], x[252], x[40], x[39], x[38], x[273], x[272], x[20], x[19], x[18], x[233], x[232], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[379], x[336], x[15], x[223], x[222], x[221]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[243], x[242], x[241], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[249], x[248], x[247], x[246], x[245], x[244], x[43], x[42], x[41], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[240], x[239], x[238], x[49], x[48], x[47], x[46], x[45], x[44], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[255], x[254], x[40], x[39], x[38], x[275], x[274], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[235], x[234], x[380], x[336], x[15], x[226], x[225], x[224]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[243], x[242], x[241], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[249], x[248], x[247], x[246], x[245], x[244], x[43], x[42], x[41], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[240], x[239], x[238], x[49], x[48], x[47], x[46], x[45], x[44], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[255], x[254], x[40], x[39], x[38], x[275], x[274], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[235], x[234], x[380], x[336], x[15], x[226], x[225], x[224]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[189], x[188], x[187], x[209], x[208], x[207], x[229], x[228], x[227], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[226], x[225], x[224], x[223], x[222], x[221], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[49], x[48], x[47], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[300], x[299], x[298], x[100], x[99], x[98], x[46], x[45], x[44], x[43], x[42], x[41], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[237], x[236], x[381], x[336], x[15], x[249], x[248], x[247]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[189], x[188], x[187], x[209], x[208], x[207], x[229], x[228], x[227], x[186], x[185], x[184], x[183], x[182], x[181], x[309], x[308], x[307], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[226], x[225], x[224], x[223], x[222], x[221], x[176], x[177], x[180], x[179], x[178], x[306], x[305], x[304], x[303], x[302], x[301], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[49], x[48], x[47], x[217], x[216], x[220], x[219], x[218], x[246], x[245], x[244], x[243], x[242], x[241], x[300], x[299], x[298], x[100], x[99], x[98], x[46], x[45], x[44], x[43], x[42], x[41], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[237], x[236], x[381], x[336], x[15], x[249], x[248], x[247]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[206], x[205], x[204], x[186], x[185], x[184], x[226], x[225], x[224], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[46], x[45], x[44], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[49], x[48], x[47], x[43], x[42], x[41], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[251], x[250], x[382], x[336], x[15], x[240], x[239], x[238]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[206], x[205], x[204], x[186], x[185], x[184], x[226], x[225], x[224], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[189], x[188], x[187], x[183], x[182], x[181], x[306], x[305], x[304], x[229], x[228], x[227], x[223], x[222], x[221], x[246], x[245], x[244], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[190], x[191], x[309], x[308], x[307], x[303], x[302], x[301], x[46], x[45], x[44], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[49], x[48], x[47], x[43], x[42], x[41], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[251], x[250], x[382], x[336], x[15], x[240], x[239], x[238]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[223], x[222], x[221], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[229], x[228], x[227], x[226], x[225], x[224], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[43], x[42], x[41], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[49], x[48], x[47], x[46], x[45], x[44], x[233], x[232], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[253], x[252], x[383], x[336], x[15], x[243], x[242], x[241]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[223], x[222], x[221], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[229], x[228], x[227], x[226], x[225], x[224], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[43], x[42], x[41], x[220], x[219], x[218], x[249], x[248], x[247], x[246], x[245], x[244], x[213], x[212], x[100], x[99], x[98], x[192], x[193], x[300], x[299], x[298], x[49], x[48], x[47], x[46], x[45], x[44], x[233], x[232], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[253], x[252], x[383], x[336], x[15], x[243], x[242], x[241]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[223], x[222], x[221], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[43], x[42], x[41], x[220], x[219], x[218], x[249], x[248], x[247], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[49], x[48], x[47], x[46], x[45], x[44], x[235], x[234], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[255], x[254], x[384], x[336], x[15], x[246], x[245], x[244]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[203], x[202], x[201], x[183], x[182], x[181], x[223], x[222], x[221], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[189], x[188], x[187], x[186], x[185], x[184], x[303], x[302], x[301], x[229], x[228], x[227], x[226], x[225], x[224], x[243], x[242], x[241], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[180], x[179], x[178], x[309], x[308], x[307], x[306], x[305], x[304], x[43], x[42], x[41], x[220], x[219], x[218], x[249], x[248], x[247], x[215], x[214], x[100], x[99], x[98], x[194], x[195], x[300], x[299], x[298], x[49], x[48], x[47], x[46], x[45], x[44], x[235], x[234], x[240], x[239], x[238], x[40], x[39], x[38], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[255], x[254], x[384], x[336], x[15], x[246], x[245], x[244]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[309], x[308], x[307], x[109], x[108], x[107], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[289], x[288], x[287], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[89], x[88], x[87], x[169], x[168], x[167], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[86], x[85], x[84], x[83], x[82], x[81], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[120], x[119], x[118], x[320], x[319], x[318], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[200], x[199], x[198], x[80], x[79], x[78], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[220], x[219], x[218], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[257], x[256], x[385], x[336], x[15], x[269], x[268], x[267]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[309], x[308], x[307], x[109], x[108], x[107], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[289], x[288], x[287], x[106], x[105], x[104], x[103], x[102], x[101], x[209], x[208], x[207], x[89], x[88], x[87], x[169], x[168], x[167], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[96], x[97], x[100], x[99], x[98], x[206], x[205], x[204], x[203], x[202], x[201], x[116], x[117], x[86], x[85], x[84], x[83], x[82], x[81], x[166], x[165], x[164], x[163], x[162], x[161], x[149], x[148], x[147], x[120], x[119], x[118], x[320], x[319], x[318], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[200], x[199], x[198], x[80], x[79], x[78], x[156], x[157], x[160], x[159], x[158], x[146], x[145], x[144], x[143], x[142], x[141], x[220], x[219], x[218], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[257], x[256], x[385], x[336], x[15], x[269], x[268], x[267]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[306], x[305], x[304], x[106], x[105], x[104], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[286], x[285], x[284], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[166], x[165], x[164], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[271], x[270], x[386], x[336], x[15], x[260], x[259], x[258]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[306], x[305], x[304], x[106], x[105], x[104], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[286], x[285], x[284], x[86], x[85], x[84], x[109], x[108], x[107], x[103], x[102], x[101], x[206], x[205], x[204], x[166], x[165], x[164], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[130], x[131], x[89], x[88], x[87], x[83], x[82], x[81], x[110], x[111], x[209], x[208], x[207], x[203], x[202], x[201], x[169], x[168], x[167], x[163], x[162], x[161], x[146], x[145], x[144], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[170], x[171], x[149], x[148], x[147], x[143], x[142], x[141], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[271], x[270], x[386], x[336], x[15], x[260], x[259], x[258]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[303], x[302], x[301], x[103], x[102], x[101], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[283], x[282], x[281], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[163], x[162], x[161], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[293], x[292], x[220], x[219], x[218], x[172], x[173], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[273], x[272], x[387], x[336], x[15], x[263], x[262], x[261]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[303], x[302], x[301], x[103], x[102], x[101], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[283], x[282], x[281], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[163], x[162], x[161], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[132], x[133], x[80], x[79], x[78], x[112], x[113], x[200], x[199], x[198], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[293], x[292], x[220], x[219], x[218], x[172], x[173], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[273], x[272], x[387], x[336], x[15], x[263], x[262], x[261]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[303], x[302], x[301], x[103], x[102], x[101], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[283], x[282], x[281], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[163], x[162], x[161], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[295], x[294], x[220], x[219], x[218], x[174], x[175], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[275], x[274], x[388], x[336], x[15], x[266], x[265], x[264]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[303], x[302], x[301], x[103], x[102], x[101], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[283], x[282], x[281], x[83], x[82], x[81], x[109], x[108], x[107], x[106], x[105], x[104], x[203], x[202], x[201], x[163], x[162], x[161], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[89], x[88], x[87], x[86], x[85], x[84], x[100], x[99], x[98], x[209], x[208], x[207], x[206], x[205], x[204], x[169], x[168], x[167], x[166], x[165], x[164], x[143], x[142], x[141], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[134], x[135], x[80], x[79], x[78], x[114], x[115], x[200], x[199], x[198], x[160], x[159], x[158], x[149], x[148], x[147], x[146], x[145], x[144], x[295], x[294], x[220], x[219], x[218], x[174], x[175], x[140], x[139], x[138], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[275], x[274], x[388], x[336], x[15], x[266], x[265], x[264]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[309], x[308], x[307], x[89], x[88], x[87], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[269], x[268], x[267], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[169], x[168], x[167], x[120], x[119], x[118], x[320], x[319], x[318], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[60], x[59], x[58], x[180], x[179], x[178], x[16], x[17], x[166], x[165], x[164], x[163], x[162], x[161], x[20], x[19], x[18], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[277], x[276], x[389], x[336], x[15], x[289], x[288], x[287]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[309], x[308], x[307], x[89], x[88], x[87], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[329], x[328], x[327], x[269], x[268], x[267], x[69], x[68], x[67], x[86], x[85], x[84], x[83], x[82], x[81], x[189], x[188], x[187], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[57], x[56], x[66], x[65], x[64], x[63], x[62], x[61], x[76], x[77], x[80], x[79], x[78], x[186], x[185], x[184], x[183], x[182], x[181], x[169], x[168], x[167], x[120], x[119], x[118], x[320], x[319], x[318], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[60], x[59], x[58], x[180], x[179], x[178], x[16], x[17], x[166], x[165], x[164], x[163], x[162], x[161], x[20], x[19], x[18], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[277], x[276], x[389], x[336], x[15], x[289], x[288], x[287]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[306], x[305], x[304], x[86], x[85], x[84], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[266], x[265], x[264], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[166], x[165], x[164], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[291], x[290], x[390], x[336], x[15], x[280], x[279], x[278]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[306], x[305], x[304], x[86], x[85], x[84], x[326], x[325], x[324], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[266], x[265], x[264], x[89], x[88], x[87], x[83], x[82], x[81], x[186], x[185], x[184], x[66], x[65], x[64], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[90], x[91], x[189], x[188], x[187], x[183], x[182], x[181], x[71], x[70], x[69], x[68], x[67], x[63], x[62], x[61], x[166], x[165], x[164], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[30], x[31], x[169], x[168], x[167], x[163], x[162], x[161], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[291], x[290], x[390], x[336], x[15], x[280], x[279], x[278]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[303], x[302], x[301], x[83], x[82], x[81], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[163], x[162], x[161], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[169], x[168], x[167], x[166], x[165], x[164], x[273], x[272], x[20], x[19], x[18], x[32], x[33], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[293], x[292], x[391], x[336], x[15], x[283], x[282], x[281]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[303], x[302], x[301], x[83], x[82], x[81], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[163], x[162], x[161], x[313], x[312], x[120], x[119], x[118], x[333], x[332], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[72], x[73], x[60], x[59], x[58], x[92], x[93], x[180], x[179], x[178], x[169], x[168], x[167], x[166], x[165], x[164], x[273], x[272], x[20], x[19], x[18], x[32], x[33], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[293], x[292], x[391], x[336], x[15], x[283], x[282], x[281]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[303], x[302], x[301], x[83], x[82], x[81], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[163], x[162], x[161], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[169], x[168], x[167], x[166], x[165], x[164], x[275], x[274], x[20], x[19], x[18], x[34], x[35], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[295], x[294], x[392], x[336], x[15], x[286], x[285], x[284]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[303], x[302], x[301], x[83], x[82], x[81], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[323], x[322], x[321], x[263], x[262], x[261], x[63], x[62], x[61], x[89], x[88], x[87], x[86], x[85], x[84], x[183], x[182], x[181], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[329], x[328], x[327], x[326], x[325], x[324], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[69], x[68], x[67], x[66], x[65], x[64], x[80], x[79], x[78], x[189], x[188], x[187], x[186], x[185], x[184], x[163], x[162], x[161], x[315], x[314], x[120], x[119], x[118], x[335], x[334], x[320], x[319], x[318], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[74], x[75], x[60], x[59], x[58], x[94], x[95], x[180], x[179], x[178], x[169], x[168], x[167], x[166], x[165], x[164], x[275], x[274], x[20], x[19], x[18], x[34], x[35], x[160], x[159], x[158], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[295], x[294], x[392], x[336], x[15], x[286], x[285], x[284]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[269], x[268], x[267], x[289], x[288], x[287], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[249], x[248], x[247], x[49], x[48], x[47], x[209], x[208], x[207], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[329], x[328], x[327], x[217], x[216], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[20], x[19], x[18], x[220], x[219], x[218], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[240], x[239], x[238], x[40], x[39], x[38], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[320], x[319], x[318], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[297], x[296], x[393], x[336], x[15], x[309], x[308], x[307]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[269], x[268], x[267], x[289], x[288], x[287], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[249], x[248], x[247], x[49], x[48], x[47], x[209], x[208], x[207], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[329], x[328], x[327], x[217], x[216], x[246], x[245], x[244], x[243], x[242], x[241], x[237], x[236], x[46], x[45], x[44], x[43], x[42], x[41], x[206], x[205], x[204], x[203], x[202], x[201], x[109], x[108], x[107], x[20], x[19], x[18], x[220], x[219], x[218], x[317], x[316], x[326], x[325], x[324], x[323], x[322], x[321], x[240], x[239], x[238], x[40], x[39], x[38], x[197], x[196], x[200], x[199], x[198], x[106], x[105], x[104], x[103], x[102], x[101], x[320], x[319], x[318], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[297], x[296], x[393], x[336], x[15], x[309], x[308], x[307]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[286], x[285], x[284], x[266], x[265], x[264], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[46], x[45], x[44], x[246], x[245], x[244], x[206], x[205], x[204], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[326], x[325], x[324], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[311], x[310], x[394], x[336], x[15], x[300], x[299], x[298]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[286], x[285], x[284], x[266], x[265], x[264], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[46], x[45], x[44], x[246], x[245], x[244], x[206], x[205], x[204], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[326], x[325], x[324], x[251], x[250], x[49], x[48], x[47], x[43], x[42], x[41], x[231], x[230], x[249], x[248], x[247], x[243], x[242], x[241], x[209], x[208], x[207], x[203], x[202], x[201], x[106], x[105], x[104], x[331], x[330], x[329], x[328], x[327], x[323], x[322], x[321], x[211], x[210], x[109], x[108], x[107], x[103], x[102], x[101], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[311], x[310], x[394], x[336], x[15], x[300], x[299], x[298]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[333], x[332], x[320], x[319], x[318], x[213], x[212], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[313], x[312], x[395], x[336], x[15], x[303], x[302], x[301]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[233], x[232], x[240], x[239], x[238], x[253], x[252], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[333], x[332], x[320], x[319], x[318], x[213], x[212], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[313], x[312], x[395], x[336], x[15], x[303], x[302], x[301]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[335], x[334], x[320], x[319], x[318], x[215], x[214], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[315], x[314], x[396], x[336], x[15], x[306], x[305], x[304]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[243], x[242], x[241], x[43], x[42], x[41], x[203], x[202], x[201], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[323], x[322], x[321], x[249], x[248], x[247], x[246], x[245], x[244], x[49], x[48], x[47], x[46], x[45], x[44], x[209], x[208], x[207], x[206], x[205], x[204], x[103], x[102], x[101], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[329], x[328], x[327], x[326], x[325], x[324], x[235], x[234], x[240], x[239], x[238], x[255], x[254], x[40], x[39], x[38], x[200], x[199], x[198], x[109], x[108], x[107], x[106], x[105], x[104], x[335], x[334], x[320], x[319], x[318], x[215], x[214], x[100], x[99], x[98], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[315], x[314], x[396], x[336], x[15], x[306], x[305], x[304]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[269], x[268], x[267], x[289], x[288], x[287], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[309], x[308], x[307], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[20], x[19], x[18], x[220], x[219], x[218], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[317], x[316], x[397], x[336], x[15], x[329], x[328], x[327]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[269], x[268], x[267], x[289], x[288], x[287], x[266], x[265], x[264], x[263], x[262], x[261], x[29], x[28], x[27], x[286], x[285], x[284], x[283], x[282], x[281], x[229], x[228], x[227], x[309], x[308], x[307], x[257], x[256], x[260], x[259], x[258], x[26], x[25], x[24], x[23], x[22], x[21], x[277], x[276], x[280], x[279], x[278], x[226], x[225], x[224], x[223], x[222], x[221], x[306], x[305], x[304], x[303], x[302], x[301], x[129], x[128], x[127], x[20], x[19], x[18], x[220], x[219], x[218], x[297], x[296], x[300], x[299], x[298], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[317], x[316], x[397], x[336], x[15], x[329], x[328], x[327]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[286], x[285], x[284], x[266], x[265], x[264], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[306], x[305], x[304], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[331], x[330], x[398], x[336], x[15], x[320], x[319], x[318]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[286], x[285], x[284], x[266], x[265], x[264], x[289], x[288], x[287], x[283], x[282], x[281], x[226], x[225], x[224], x[269], x[268], x[267], x[263], x[262], x[261], x[26], x[25], x[24], x[306], x[305], x[304], x[291], x[290], x[229], x[228], x[227], x[223], x[222], x[221], x[271], x[270], x[29], x[28], x[27], x[23], x[22], x[21], x[309], x[308], x[307], x[303], x[302], x[301], x[126], x[125], x[124], x[311], x[310], x[129], x[128], x[127], x[123], x[122], x[121], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[331], x[330], x[398], x[336], x[15], x[320], x[319], x[318]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[303], x[302], x[301], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[313], x[312], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[333], x[332], x[399], x[336], x[15], x[323], x[322], x[321]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[303], x[302], x[301], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[293], x[292], x[220], x[219], x[218], x[273], x[272], x[20], x[19], x[18], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[313], x[312], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[333], x[332], x[399], x[336], x[15], x[323], x[322], x[321]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[303], x[302], x[301], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[315], x[314], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[335], x[334], x[400], x[336], x[15], x[326], x[325], x[324]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[283], x[282], x[281], x[263], x[262], x[261], x[289], x[288], x[287], x[286], x[285], x[284], x[223], x[222], x[221], x[269], x[268], x[267], x[266], x[265], x[264], x[23], x[22], x[21], x[303], x[302], x[301], x[280], x[279], x[278], x[229], x[228], x[227], x[226], x[225], x[224], x[260], x[259], x[258], x[29], x[28], x[27], x[26], x[25], x[24], x[309], x[308], x[307], x[306], x[305], x[304], x[123], x[122], x[121], x[295], x[294], x[220], x[219], x[218], x[275], x[274], x[20], x[19], x[18], x[300], x[299], x[298], x[129], x[128], x[127], x[126], x[125], x[124], x[315], x[314], x[120], x[119], x[118], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[335], x[334], x[400], x[336], x[15], x[326], x[325], x[324]}), .y(y[267]));
endmodule

