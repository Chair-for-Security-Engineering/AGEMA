/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module Midori64_HPC2_BDDcudd_Pipeline_d1 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, DataIn_s1, Fresh, DataOut_s0, done, DataOut_s1);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [63:0] DataIn_s1 ;
    input [230:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    wire signal_201 ;
    wire signal_203 ;
    wire signal_205 ;
    wire signal_207 ;
    wire signal_209 ;
    wire signal_211 ;
    wire signal_213 ;
    wire signal_215 ;
    wire signal_217 ;
    wire signal_219 ;
    wire signal_221 ;
    wire signal_223 ;
    wire signal_225 ;
    wire signal_227 ;
    wire signal_229 ;
    wire signal_231 ;
    wire signal_233 ;
    wire signal_235 ;
    wire signal_237 ;
    wire signal_239 ;
    wire signal_241 ;
    wire signal_243 ;
    wire signal_245 ;
    wire signal_247 ;
    wire signal_249 ;
    wire signal_251 ;
    wire signal_253 ;
    wire signal_255 ;
    wire signal_257 ;
    wire signal_259 ;
    wire signal_261 ;
    wire signal_263 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1625 ;
    wire signal_1628 ;
    wire signal_1631 ;
    wire signal_1634 ;
    wire signal_1637 ;
    wire signal_1640 ;
    wire signal_1643 ;
    wire signal_1646 ;
    wire signal_1649 ;
    wire signal_1652 ;
    wire signal_1655 ;
    wire signal_1658 ;
    wire signal_1661 ;
    wire signal_1664 ;
    wire signal_1667 ;
    wire signal_1670 ;
    wire signal_1673 ;
    wire signal_1676 ;
    wire signal_1679 ;
    wire signal_1682 ;
    wire signal_1685 ;
    wire signal_1688 ;
    wire signal_1691 ;
    wire signal_1694 ;
    wire signal_1697 ;
    wire signal_1700 ;
    wire signal_1703 ;
    wire signal_1706 ;
    wire signal_1709 ;
    wire signal_1712 ;
    wire signal_1715 ;
    wire signal_1718 ;
    wire signal_1721 ;
    wire signal_1724 ;
    wire signal_1727 ;
    wire signal_1730 ;
    wire signal_1733 ;
    wire signal_1736 ;
    wire signal_1739 ;
    wire signal_1742 ;
    wire signal_1745 ;
    wire signal_1748 ;
    wire signal_1751 ;
    wire signal_1754 ;
    wire signal_1757 ;
    wire signal_1760 ;
    wire signal_1763 ;
    wire signal_1766 ;
    wire signal_1769 ;
    wire signal_1772 ;
    wire signal_1775 ;
    wire signal_1778 ;
    wire signal_1781 ;
    wire signal_1784 ;
    wire signal_1787 ;
    wire signal_1790 ;
    wire signal_1793 ;
    wire signal_1796 ;
    wire signal_1799 ;
    wire signal_1802 ;
    wire signal_1805 ;
    wire signal_1808 ;
    wire signal_1811 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1891 ;
    wire signal_1893 ;
    wire signal_1895 ;
    wire signal_1897 ;
    wire signal_1899 ;
    wire signal_1901 ;
    wire signal_1903 ;
    wire signal_1905 ;
    wire signal_1907 ;
    wire signal_1909 ;
    wire signal_1911 ;
    wire signal_1913 ;
    wire signal_1915 ;
    wire signal_1917 ;
    wire signal_1919 ;
    wire signal_1921 ;
    wire signal_1923 ;
    wire signal_1925 ;
    wire signal_1927 ;
    wire signal_1929 ;
    wire signal_1931 ;
    wire signal_1933 ;
    wire signal_1935 ;
    wire signal_1937 ;
    wire signal_1939 ;
    wire signal_1941 ;
    wire signal_1943 ;
    wire signal_1945 ;
    wire signal_1947 ;
    wire signal_1949 ;
    wire signal_1951 ;
    wire signal_1953 ;
    wire signal_1955 ;
    wire signal_1957 ;
    wire signal_1959 ;
    wire signal_1961 ;
    wire signal_1963 ;
    wire signal_1965 ;
    wire signal_1967 ;
    wire signal_1969 ;
    wire signal_1971 ;
    wire signal_1973 ;
    wire signal_1975 ;
    wire signal_1977 ;
    wire signal_1979 ;
    wire signal_1981 ;
    wire signal_1983 ;
    wire signal_1985 ;
    wire signal_1987 ;
    wire signal_1989 ;
    wire signal_1991 ;
    wire signal_1993 ;
    wire signal_1995 ;
    wire signal_1997 ;
    wire signal_1999 ;
    wire signal_2001 ;
    wire signal_2003 ;
    wire signal_2005 ;
    wire signal_2007 ;
    wire signal_2009 ;
    wire signal_2011 ;
    wire signal_2013 ;
    wire signal_2015 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3111 ;
    wire signal_3113 ;
    wire signal_3115 ;
    wire signal_3117 ;
    wire signal_3119 ;
    wire signal_3121 ;
    wire signal_3123 ;
    wire signal_3125 ;
    wire signal_3127 ;
    wire signal_3129 ;
    wire signal_3131 ;
    wire signal_3133 ;
    wire signal_3135 ;
    wire signal_3137 ;
    wire signal_3139 ;
    wire signal_3141 ;
    wire signal_3143 ;
    wire signal_3145 ;
    wire signal_3147 ;
    wire signal_3149 ;
    wire signal_3151 ;
    wire signal_3153 ;
    wire signal_3155 ;
    wire signal_3157 ;
    wire signal_3159 ;
    wire signal_3161 ;
    wire signal_3163 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_0 ( .a ({key_s1[73], key_s0[73]}), .b ({key_s1[9], key_s0[9]}), .c ({signal_1625, signal_914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1 ( .a ({key_s1[72], key_s0[72]}), .b ({key_s1[8], key_s0[8]}), .c ({signal_1628, signal_915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_2 ( .a ({key_s1[71], key_s0[71]}), .b ({key_s1[7], key_s0[7]}), .c ({signal_1631, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3 ( .a ({key_s1[6], key_s0[6]}), .b ({key_s1[70], key_s0[70]}), .c ({signal_1634, signal_917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4 ( .a ({key_s1[127], key_s0[127]}), .b ({key_s1[63], key_s0[63]}), .c ({signal_1637, signal_860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5 ( .a ({key_s1[126], key_s0[126]}), .b ({key_s1[62], key_s0[62]}), .c ({signal_1640, signal_861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6 ( .a ({key_s1[125], key_s0[125]}), .b ({key_s1[61], key_s0[61]}), .c ({signal_1643, signal_862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7 ( .a ({key_s1[124], key_s0[124]}), .b ({key_s1[60], key_s0[60]}), .c ({signal_1646, signal_863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_8 ( .a ({key_s1[5], key_s0[5]}), .b ({key_s1[69], key_s0[69]}), .c ({signal_1649, signal_918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_9 ( .a ({key_s1[123], key_s0[123]}), .b ({key_s1[59], key_s0[59]}), .c ({signal_1652, signal_864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_10 ( .a ({key_s1[122], key_s0[122]}), .b ({key_s1[58], key_s0[58]}), .c ({signal_1655, signal_865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_11 ( .a ({key_s1[121], key_s0[121]}), .b ({key_s1[57], key_s0[57]}), .c ({signal_1658, signal_866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_12 ( .a ({key_s1[120], key_s0[120]}), .b ({key_s1[56], key_s0[56]}), .c ({signal_1661, signal_867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_13 ( .a ({key_s1[119], key_s0[119]}), .b ({key_s1[55], key_s0[55]}), .c ({signal_1664, signal_868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_14 ( .a ({key_s1[118], key_s0[118]}), .b ({key_s1[54], key_s0[54]}), .c ({signal_1667, signal_869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_15 ( .a ({key_s1[117], key_s0[117]}), .b ({key_s1[53], key_s0[53]}), .c ({signal_1670, signal_870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_16 ( .a ({key_s1[116], key_s0[116]}), .b ({key_s1[52], key_s0[52]}), .c ({signal_1673, signal_871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_17 ( .a ({key_s1[115], key_s0[115]}), .b ({key_s1[51], key_s0[51]}), .c ({signal_1676, signal_872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_18 ( .a ({key_s1[114], key_s0[114]}), .b ({key_s1[50], key_s0[50]}), .c ({signal_1679, signal_873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_19 ( .a ({key_s1[4], key_s0[4]}), .b ({key_s1[68], key_s0[68]}), .c ({signal_1682, signal_919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_20 ( .a ({key_s1[113], key_s0[113]}), .b ({key_s1[49], key_s0[49]}), .c ({signal_1685, signal_874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_21 ( .a ({key_s1[112], key_s0[112]}), .b ({key_s1[48], key_s0[48]}), .c ({signal_1688, signal_875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_22 ( .a ({key_s1[111], key_s0[111]}), .b ({key_s1[47], key_s0[47]}), .c ({signal_1691, signal_876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_23 ( .a ({key_s1[110], key_s0[110]}), .b ({key_s1[46], key_s0[46]}), .c ({signal_1694, signal_877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_24 ( .a ({key_s1[109], key_s0[109]}), .b ({key_s1[45], key_s0[45]}), .c ({signal_1697, signal_878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_25 ( .a ({key_s1[108], key_s0[108]}), .b ({key_s1[44], key_s0[44]}), .c ({signal_1700, signal_879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_26 ( .a ({key_s1[107], key_s0[107]}), .b ({key_s1[43], key_s0[43]}), .c ({signal_1703, signal_880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_27 ( .a ({key_s1[106], key_s0[106]}), .b ({key_s1[42], key_s0[42]}), .c ({signal_1706, signal_881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_28 ( .a ({key_s1[105], key_s0[105]}), .b ({key_s1[41], key_s0[41]}), .c ({signal_1709, signal_882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_29 ( .a ({key_s1[104], key_s0[104]}), .b ({key_s1[40], key_s0[40]}), .c ({signal_1712, signal_883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_30 ( .a ({key_s1[3], key_s0[3]}), .b ({key_s1[67], key_s0[67]}), .c ({signal_1715, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_31 ( .a ({key_s1[103], key_s0[103]}), .b ({key_s1[39], key_s0[39]}), .c ({signal_1718, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_32 ( .a ({key_s1[102], key_s0[102]}), .b ({key_s1[38], key_s0[38]}), .c ({signal_1721, signal_885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_33 ( .a ({key_s1[101], key_s0[101]}), .b ({key_s1[37], key_s0[37]}), .c ({signal_1724, signal_886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_34 ( .a ({key_s1[100], key_s0[100]}), .b ({key_s1[36], key_s0[36]}), .c ({signal_1727, signal_887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_35 ( .a ({key_s1[35], key_s0[35]}), .b ({key_s1[99], key_s0[99]}), .c ({signal_1730, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_36 ( .a ({key_s1[34], key_s0[34]}), .b ({key_s1[98], key_s0[98]}), .c ({signal_1733, signal_889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_37 ( .a ({key_s1[33], key_s0[33]}), .b ({key_s1[97], key_s0[97]}), .c ({signal_1736, signal_890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_38 ( .a ({key_s1[32], key_s0[32]}), .b ({key_s1[96], key_s0[96]}), .c ({signal_1739, signal_891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_39 ( .a ({key_s1[31], key_s0[31]}), .b ({key_s1[95], key_s0[95]}), .c ({signal_1742, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_40 ( .a ({key_s1[30], key_s0[30]}), .b ({key_s1[94], key_s0[94]}), .c ({signal_1745, signal_893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_41 ( .a ({key_s1[2], key_s0[2]}), .b ({key_s1[66], key_s0[66]}), .c ({signal_1748, signal_921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_42 ( .a ({key_s1[29], key_s0[29]}), .b ({key_s1[93], key_s0[93]}), .c ({signal_1751, signal_894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_43 ( .a ({key_s1[28], key_s0[28]}), .b ({key_s1[92], key_s0[92]}), .c ({signal_1754, signal_895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_44 ( .a ({key_s1[27], key_s0[27]}), .b ({key_s1[91], key_s0[91]}), .c ({signal_1757, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_45 ( .a ({key_s1[26], key_s0[26]}), .b ({key_s1[90], key_s0[90]}), .c ({signal_1760, signal_897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_46 ( .a ({key_s1[25], key_s0[25]}), .b ({key_s1[89], key_s0[89]}), .c ({signal_1763, signal_898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_47 ( .a ({key_s1[24], key_s0[24]}), .b ({key_s1[88], key_s0[88]}), .c ({signal_1766, signal_899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_48 ( .a ({key_s1[23], key_s0[23]}), .b ({key_s1[87], key_s0[87]}), .c ({signal_1769, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_49 ( .a ({key_s1[22], key_s0[22]}), .b ({key_s1[86], key_s0[86]}), .c ({signal_1772, signal_901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_50 ( .a ({key_s1[21], key_s0[21]}), .b ({key_s1[85], key_s0[85]}), .c ({signal_1775, signal_902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_51 ( .a ({key_s1[20], key_s0[20]}), .b ({key_s1[84], key_s0[84]}), .c ({signal_1778, signal_903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_52 ( .a ({key_s1[1], key_s0[1]}), .b ({key_s1[65], key_s0[65]}), .c ({signal_1781, signal_922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_53 ( .a ({key_s1[19], key_s0[19]}), .b ({key_s1[83], key_s0[83]}), .c ({signal_1784, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_54 ( .a ({key_s1[18], key_s0[18]}), .b ({key_s1[82], key_s0[82]}), .c ({signal_1787, signal_905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_55 ( .a ({key_s1[17], key_s0[17]}), .b ({key_s1[81], key_s0[81]}), .c ({signal_1790, signal_906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_56 ( .a ({key_s1[16], key_s0[16]}), .b ({key_s1[80], key_s0[80]}), .c ({signal_1793, signal_907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_57 ( .a ({key_s1[15], key_s0[15]}), .b ({key_s1[79], key_s0[79]}), .c ({signal_1796, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_58 ( .a ({key_s1[14], key_s0[14]}), .b ({key_s1[78], key_s0[78]}), .c ({signal_1799, signal_909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_59 ( .a ({key_s1[13], key_s0[13]}), .b ({key_s1[77], key_s0[77]}), .c ({signal_1802, signal_910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_60 ( .a ({key_s1[12], key_s0[12]}), .b ({key_s1[76], key_s0[76]}), .c ({signal_1805, signal_911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_61 ( .a ({key_s1[11], key_s0[11]}), .b ({key_s1[75], key_s0[75]}), .c ({signal_1808, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_62 ( .a ({key_s1[10], key_s0[10]}), .b ({key_s1[74], key_s0[74]}), .c ({signal_1811, signal_913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_63 ( .a ({key_s1[0], key_s0[0]}), .b ({key_s1[64], key_s0[64]}), .c ({signal_1814, signal_923}) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_266), .A2 (signal_267), .ZN (signal_265) ) ;
    NAND2_X1 cell_65 ( .A1 (signal_927), .A2 (signal_926), .ZN (signal_267) ) ;
    NAND2_X1 cell_66 ( .A1 (signal_925), .A2 (signal_924), .ZN (signal_266) ) ;
    INV_X1 cell_67 ( .A (signal_268), .ZN (signal_278) ) ;
    MUX2_X1 cell_68 ( .S (signal_281), .A (signal_269), .B (signal_270), .Z (signal_268) ) ;
    NOR2_X1 cell_69 ( .A1 (reset), .A2 (signal_271), .ZN (signal_282) ) ;
    XNOR2_X1 cell_70 ( .A (signal_927), .B (signal_926), .ZN (signal_271) ) ;
    MUX2_X1 cell_71 ( .S (signal_924), .A (signal_272), .B (signal_273), .Z (signal_280) ) ;
    NAND2_X1 cell_72 ( .A1 (signal_269), .A2 (signal_274), .ZN (signal_273) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_281), .A2 (signal_277), .ZN (signal_274) ) ;
    NOR2_X1 cell_74 ( .A1 (signal_275), .A2 (signal_283), .ZN (signal_269) ) ;
    NOR2_X1 cell_75 ( .A1 (signal_926), .A2 (reset), .ZN (signal_275) ) ;
    NOR2_X1 cell_76 ( .A1 (signal_281), .A2 (signal_270), .ZN (signal_272) ) ;
    NAND2_X1 cell_77 ( .A1 (signal_926), .A2 (signal_276), .ZN (signal_270) ) ;
    NOR2_X1 cell_78 ( .A1 (reset), .A2 (signal_279), .ZN (signal_276) ) ;
    NOR2_X1 cell_79 ( .A1 (reset), .A2 (signal_927), .ZN (signal_283) ) ;
    INV_X1 cell_80 ( .A (reset), .ZN (signal_277) ) ;
    INV_X1 cell_81 ( .A (signal_927), .ZN (signal_279) ) ;
    INV_X1 cell_85 ( .A (signal_925), .ZN (signal_281) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_153 ( .a ({signal_1625, signal_914}), .b ({DataIn_s1[9], DataIn_s0[9]}), .c ({signal_1891, signal_982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_154 ( .a ({signal_1628, signal_915}), .b ({DataIn_s1[8], DataIn_s0[8]}), .c ({signal_1893, signal_983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_155 ( .a ({signal_1631, signal_916}), .b ({DataIn_s1[7], DataIn_s0[7]}), .c ({signal_1895, signal_984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_156 ( .a ({signal_1634, signal_917}), .b ({DataIn_s1[6], DataIn_s0[6]}), .c ({signal_1897, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_157 ( .a ({signal_1637, signal_860}), .b ({DataIn_s1[63], DataIn_s0[63]}), .c ({signal_1899, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_158 ( .a ({signal_1640, signal_861}), .b ({DataIn_s1[62], DataIn_s0[62]}), .c ({signal_1901, signal_929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_159 ( .a ({signal_1643, signal_862}), .b ({DataIn_s1[61], DataIn_s0[61]}), .c ({signal_1903, signal_930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_160 ( .a ({signal_1646, signal_863}), .b ({DataIn_s1[60], DataIn_s0[60]}), .c ({signal_1905, signal_931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_161 ( .a ({signal_1649, signal_918}), .b ({DataIn_s1[5], DataIn_s0[5]}), .c ({signal_1907, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_162 ( .a ({signal_1652, signal_864}), .b ({DataIn_s1[59], DataIn_s0[59]}), .c ({signal_1909, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_163 ( .a ({signal_1655, signal_865}), .b ({DataIn_s1[58], DataIn_s0[58]}), .c ({signal_1911, signal_933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_164 ( .a ({signal_1658, signal_866}), .b ({DataIn_s1[57], DataIn_s0[57]}), .c ({signal_1913, signal_934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_165 ( .a ({signal_1661, signal_867}), .b ({DataIn_s1[56], DataIn_s0[56]}), .c ({signal_1915, signal_935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_166 ( .a ({signal_1664, signal_868}), .b ({DataIn_s1[55], DataIn_s0[55]}), .c ({signal_1917, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_167 ( .a ({signal_1667, signal_869}), .b ({DataIn_s1[54], DataIn_s0[54]}), .c ({signal_1919, signal_937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_168 ( .a ({signal_1670, signal_870}), .b ({DataIn_s1[53], DataIn_s0[53]}), .c ({signal_1921, signal_938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_169 ( .a ({signal_1673, signal_871}), .b ({DataIn_s1[52], DataIn_s0[52]}), .c ({signal_1923, signal_939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_170 ( .a ({signal_1676, signal_872}), .b ({DataIn_s1[51], DataIn_s0[51]}), .c ({signal_1925, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_171 ( .a ({signal_1679, signal_873}), .b ({DataIn_s1[50], DataIn_s0[50]}), .c ({signal_1927, signal_941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_172 ( .a ({signal_1682, signal_919}), .b ({DataIn_s1[4], DataIn_s0[4]}), .c ({signal_1929, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_173 ( .a ({signal_1685, signal_874}), .b ({DataIn_s1[49], DataIn_s0[49]}), .c ({signal_1931, signal_942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_174 ( .a ({signal_1688, signal_875}), .b ({DataIn_s1[48], DataIn_s0[48]}), .c ({signal_1933, signal_943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_175 ( .a ({signal_1691, signal_876}), .b ({DataIn_s1[47], DataIn_s0[47]}), .c ({signal_1935, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_176 ( .a ({signal_1694, signal_877}), .b ({DataIn_s1[46], DataIn_s0[46]}), .c ({signal_1937, signal_945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_177 ( .a ({signal_1697, signal_878}), .b ({DataIn_s1[45], DataIn_s0[45]}), .c ({signal_1939, signal_946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .a ({signal_1700, signal_879}), .b ({DataIn_s1[44], DataIn_s0[44]}), .c ({signal_1941, signal_947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .a ({signal_1703, signal_880}), .b ({DataIn_s1[43], DataIn_s0[43]}), .c ({signal_1943, signal_948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .a ({signal_1706, signal_881}), .b ({DataIn_s1[42], DataIn_s0[42]}), .c ({signal_1945, signal_949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .a ({signal_1709, signal_882}), .b ({DataIn_s1[41], DataIn_s0[41]}), .c ({signal_1947, signal_950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .a ({signal_1712, signal_883}), .b ({DataIn_s1[40], DataIn_s0[40]}), .c ({signal_1949, signal_951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .a ({signal_1715, signal_920}), .b ({DataIn_s1[3], DataIn_s0[3]}), .c ({signal_1951, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .a ({signal_1718, signal_884}), .b ({DataIn_s1[39], DataIn_s0[39]}), .c ({signal_1953, signal_952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .a ({signal_1721, signal_885}), .b ({DataIn_s1[38], DataIn_s0[38]}), .c ({signal_1955, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .a ({signal_1724, signal_886}), .b ({DataIn_s1[37], DataIn_s0[37]}), .c ({signal_1957, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .a ({signal_1727, signal_887}), .b ({DataIn_s1[36], DataIn_s0[36]}), .c ({signal_1959, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .a ({signal_1730, signal_888}), .b ({DataIn_s1[35], DataIn_s0[35]}), .c ({signal_1961, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .a ({signal_1733, signal_889}), .b ({DataIn_s1[34], DataIn_s0[34]}), .c ({signal_1963, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .a ({signal_1736, signal_890}), .b ({DataIn_s1[33], DataIn_s0[33]}), .c ({signal_1965, signal_958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .a ({signal_1739, signal_891}), .b ({DataIn_s1[32], DataIn_s0[32]}), .c ({signal_1967, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .a ({signal_1742, signal_892}), .b ({DataIn_s1[31], DataIn_s0[31]}), .c ({signal_1969, signal_960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_193 ( .a ({signal_1745, signal_893}), .b ({DataIn_s1[30], DataIn_s0[30]}), .c ({signal_1971, signal_961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_194 ( .a ({signal_1748, signal_921}), .b ({DataIn_s1[2], DataIn_s0[2]}), .c ({signal_1973, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_195 ( .a ({signal_1751, signal_894}), .b ({DataIn_s1[29], DataIn_s0[29]}), .c ({signal_1975, signal_962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_196 ( .a ({signal_1754, signal_895}), .b ({DataIn_s1[28], DataIn_s0[28]}), .c ({signal_1977, signal_963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .a ({signal_1757, signal_896}), .b ({DataIn_s1[27], DataIn_s0[27]}), .c ({signal_1979, signal_964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .a ({signal_1760, signal_897}), .b ({DataIn_s1[26], DataIn_s0[26]}), .c ({signal_1981, signal_965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .a ({signal_1763, signal_898}), .b ({DataIn_s1[25], DataIn_s0[25]}), .c ({signal_1983, signal_966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .a ({signal_1766, signal_899}), .b ({DataIn_s1[24], DataIn_s0[24]}), .c ({signal_1985, signal_967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .a ({signal_1769, signal_900}), .b ({DataIn_s1[23], DataIn_s0[23]}), .c ({signal_1987, signal_968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .a ({signal_1772, signal_901}), .b ({DataIn_s1[22], DataIn_s0[22]}), .c ({signal_1989, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .a ({signal_1775, signal_902}), .b ({DataIn_s1[21], DataIn_s0[21]}), .c ({signal_1991, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .a ({signal_1778, signal_903}), .b ({DataIn_s1[20], DataIn_s0[20]}), .c ({signal_1993, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .a ({signal_1781, signal_922}), .b ({DataIn_s1[1], DataIn_s0[1]}), .c ({signal_1995, signal_990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .a ({signal_1784, signal_904}), .b ({DataIn_s1[19], DataIn_s0[19]}), .c ({signal_1997, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_207 ( .a ({signal_1787, signal_905}), .b ({DataIn_s1[18], DataIn_s0[18]}), .c ({signal_1999, signal_973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_208 ( .a ({signal_1790, signal_906}), .b ({DataIn_s1[17], DataIn_s0[17]}), .c ({signal_2001, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_209 ( .a ({signal_1793, signal_907}), .b ({DataIn_s1[16], DataIn_s0[16]}), .c ({signal_2003, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_210 ( .a ({signal_1796, signal_908}), .b ({DataIn_s1[15], DataIn_s0[15]}), .c ({signal_2005, signal_976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_211 ( .a ({signal_1799, signal_909}), .b ({DataIn_s1[14], DataIn_s0[14]}), .c ({signal_2007, signal_977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_212 ( .a ({signal_1802, signal_910}), .b ({DataIn_s1[13], DataIn_s0[13]}), .c ({signal_2009, signal_978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_213 ( .a ({signal_1805, signal_911}), .b ({DataIn_s1[12], DataIn_s0[12]}), .c ({signal_2011, signal_979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_214 ( .a ({signal_1808, signal_912}), .b ({DataIn_s1[11], DataIn_s0[11]}), .c ({signal_2013, signal_980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .a ({signal_1811, signal_913}), .b ({DataIn_s1[10], DataIn_s0[10]}), .c ({signal_2015, signal_981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .a ({signal_1814, signal_923}), .b ({DataIn_s1[0], DataIn_s0[0]}), .c ({signal_2017, signal_991}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .a ({signal_1820, signal_310}), .b ({1'b0, signal_1453}), .c ({signal_2566, signal_286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_290 ( .a ({signal_2186, signal_362}), .b ({1'b0, signal_1440}), .c ({signal_2622, signal_287}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_296 ( .a ({signal_2182, signal_358}), .b ({1'b0, signal_1441}), .c ({signal_2623, signal_288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_301 ( .a ({signal_2178, signal_354}), .b ({1'b0, signal_1442}), .c ({signal_2624, signal_289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_305 ( .a ({signal_1819, signal_306}), .b ({1'b0, signal_1454}), .c ({signal_2625, signal_290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_308 ( .a ({signal_2174, signal_350}), .b ({1'b0, signal_1443}), .c ({signal_2712, signal_291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_313 ( .a ({signal_2170, signal_346}), .b ({1'b0, signal_1444}), .c ({signal_2573, signal_292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_318 ( .a ({signal_2166, signal_342}), .b ({1'b0, signal_1445}), .c ({signal_2626, signal_293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_324 ( .a ({signal_2162, signal_338}), .b ({1'b0, signal_1446}), .c ({signal_2576, signal_294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_329 ( .a ({signal_2158, signal_334}), .b ({1'b0, signal_1447}), .c ({signal_2627, signal_295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_335 ( .a ({signal_2154, signal_330}), .b ({1'b0, signal_1448}), .c ({signal_2690, signal_296}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_340 ( .a ({signal_2151, signal_326}), .b ({1'b0, signal_1449}), .c ({signal_2628, signal_297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_345 ( .a ({signal_2147, signal_322}), .b ({1'b0, signal_1450}), .c ({signal_2582, signal_298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_351 ( .a ({signal_2143, signal_318}), .b ({1'b0, signal_1451}), .c ({signal_2629, signal_299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_356 ( .a ({signal_2142, signal_314}), .b ({1'b0, signal_1452}), .c ({signal_2630, signal_300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_360 ( .a ({signal_1815, signal_302}), .b ({1'b0, signal_1455}), .c ({signal_2631, signal_301}) ) ;
    NAND2_X1 cell_361 ( .A1 (signal_366), .A2 (signal_367), .ZN (signal_1446) ) ;
    NOR2_X1 cell_362 ( .A1 (signal_368), .A2 (signal_369), .ZN (signal_366) ) ;
    OR2_X1 cell_363 ( .A1 (signal_370), .A2 (signal_371), .ZN (signal_369) ) ;
    NAND2_X1 cell_364 ( .A1 (signal_372), .A2 (signal_373), .ZN (signal_1447) ) ;
    NAND2_X1 cell_365 ( .A1 (signal_374), .A2 (signal_375), .ZN (signal_1448) ) ;
    NOR2_X1 cell_366 ( .A1 (signal_1444), .A2 (signal_376), .ZN (signal_375) ) ;
    NAND2_X1 cell_367 ( .A1 (signal_377), .A2 (signal_378), .ZN (signal_376) ) ;
    NOR2_X1 cell_368 ( .A1 (signal_379), .A2 (signal_380), .ZN (signal_377) ) ;
    NAND2_X1 cell_369 ( .A1 (signal_381), .A2 (signal_382), .ZN (signal_1449) ) ;
    NOR2_X1 cell_370 ( .A1 (signal_383), .A2 (signal_384), .ZN (signal_382) ) ;
    NAND2_X1 cell_371 ( .A1 (signal_385), .A2 (signal_386), .ZN (signal_1450) ) ;
    NOR2_X1 cell_372 ( .A1 (signal_371), .A2 (signal_387), .ZN (signal_386) ) ;
    NAND2_X1 cell_373 ( .A1 (signal_388), .A2 (signal_378), .ZN (signal_387) ) ;
    NAND2_X1 cell_374 ( .A1 (signal_389), .A2 (signal_388), .ZN (signal_1451) ) ;
    NOR2_X1 cell_375 ( .A1 (signal_390), .A2 (signal_391), .ZN (signal_388) ) ;
    NAND2_X1 cell_376 ( .A1 (signal_392), .A2 (signal_393), .ZN (signal_1452) ) ;
    NOR2_X1 cell_377 ( .A1 (signal_368), .A2 (signal_394), .ZN (signal_392) ) ;
    NAND2_X1 cell_378 ( .A1 (signal_395), .A2 (signal_378), .ZN (signal_394) ) ;
    INV_X1 cell_379 ( .A (signal_396), .ZN (signal_395) ) ;
    OR2_X1 cell_380 ( .A1 (signal_368), .A2 (signal_397), .ZN (signal_1453) ) ;
    NAND2_X1 cell_381 ( .A1 (signal_381), .A2 (signal_398), .ZN (signal_397) ) ;
    NOR2_X1 cell_382 ( .A1 (signal_399), .A2 (signal_371), .ZN (signal_381) ) ;
    NAND2_X1 cell_383 ( .A1 (signal_400), .A2 (signal_373), .ZN (signal_368) ) ;
    NAND2_X1 cell_384 ( .A1 (signal_401), .A2 (signal_402), .ZN (signal_1454) ) ;
    NOR2_X1 cell_385 ( .A1 (signal_396), .A2 (signal_403), .ZN (signal_402) ) ;
    OR2_X1 cell_386 ( .A1 (signal_371), .A2 (signal_379), .ZN (signal_403) ) ;
    INV_X1 cell_387 ( .A (signal_400), .ZN (signal_379) ) ;
    NAND2_X1 cell_388 ( .A1 (signal_404), .A2 (signal_405), .ZN (signal_400) ) ;
    NAND2_X1 cell_389 ( .A1 (signal_406), .A2 (signal_407), .ZN (signal_405) ) ;
    NOR2_X1 cell_390 ( .A1 (signal_455), .A2 (signal_408), .ZN (signal_371) ) ;
    MUX2_X1 cell_391 ( .S (signal_925), .A (signal_409), .B (signal_410), .Z (signal_408) ) ;
    NAND2_X1 cell_392 ( .A1 (signal_411), .A2 (signal_412), .ZN (signal_1440) ) ;
    NOR2_X1 cell_393 ( .A1 (signal_383), .A2 (signal_396), .ZN (signal_411) ) ;
    NAND2_X1 cell_394 ( .A1 (signal_413), .A2 (signal_389), .ZN (signal_1441) ) ;
    NOR2_X1 cell_395 ( .A1 (signal_414), .A2 (signal_415), .ZN (signal_389) ) ;
    NAND2_X1 cell_396 ( .A1 (signal_367), .A2 (signal_378), .ZN (signal_415) ) ;
    OR2_X1 cell_397 ( .A1 (signal_454), .A2 (signal_416), .ZN (signal_378) ) ;
    MUX2_X1 cell_398 ( .S (signal_925), .A (signal_417), .B (signal_418), .Z (signal_416) ) ;
    NAND2_X1 cell_399 ( .A1 (signal_398), .A2 (signal_419), .ZN (signal_1442) ) ;
    NOR2_X1 cell_400 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_419) ) ;
    INV_X1 cell_401 ( .A (signal_413), .ZN (signal_421) ) ;
    NOR2_X1 cell_402 ( .A1 (signal_422), .A2 (signal_391), .ZN (signal_398) ) ;
    NAND2_X1 cell_403 ( .A1 (signal_423), .A2 (signal_393), .ZN (signal_1443) ) ;
    INV_X1 cell_404 ( .A (signal_399), .ZN (signal_393) ) ;
    NOR2_X1 cell_405 ( .A1 (signal_380), .A2 (signal_424), .ZN (signal_423) ) ;
    NAND2_X1 cell_406 ( .A1 (signal_372), .A2 (signal_413), .ZN (signal_424) ) ;
    NOR2_X1 cell_407 ( .A1 (signal_390), .A2 (signal_414), .ZN (signal_372) ) ;
    NAND2_X1 cell_408 ( .A1 (signal_385), .A2 (signal_425), .ZN (signal_414) ) ;
    NAND2_X1 cell_409 ( .A1 (signal_454), .A2 (signal_426), .ZN (signal_425) ) ;
    NAND2_X1 cell_410 ( .A1 (signal_418), .A2 (signal_406), .ZN (signal_426) ) ;
    NOR2_X1 cell_411 ( .A1 (signal_383), .A2 (signal_427), .ZN (signal_385) ) ;
    NOR2_X1 cell_412 ( .A1 (signal_455), .A2 (signal_428), .ZN (signal_427) ) ;
    MUX2_X1 cell_413 ( .S (signal_925), .A (signal_407), .B (signal_417), .Z (signal_428) ) ;
    NOR2_X1 cell_414 ( .A1 (signal_454), .A2 (signal_429), .ZN (signal_383) ) ;
    MUX2_X1 cell_415 ( .S (signal_925), .A (signal_409), .B (signal_430), .Z (signal_429) ) ;
    OR2_X1 cell_416 ( .A1 (signal_384), .A2 (signal_370), .ZN (signal_1444) ) ;
    NAND2_X1 cell_417 ( .A1 (signal_413), .A2 (signal_373), .ZN (signal_384) ) ;
    NAND2_X1 cell_418 ( .A1 (signal_431), .A2 (signal_432), .ZN (signal_373) ) ;
    AND2_X1 cell_419 ( .A1 (signal_455), .A2 (signal_925), .ZN (signal_432) ) ;
    NOR2_X1 cell_420 ( .A1 (signal_433), .A2 (signal_396), .ZN (signal_413) ) ;
    NOR2_X1 cell_421 ( .A1 (signal_454), .A2 (signal_434), .ZN (signal_396) ) ;
    MUX2_X1 cell_422 ( .S (signal_925), .A (signal_418), .B (signal_417), .Z (signal_434) ) ;
    NOR2_X1 cell_423 ( .A1 (signal_454), .A2 (signal_435), .ZN (signal_433) ) ;
    MUX2_X1 cell_424 ( .S (signal_925), .A (signal_430), .B (signal_409), .Z (signal_435) ) ;
    NAND2_X1 cell_425 ( .A1 (signal_436), .A2 (signal_412), .ZN (signal_1445) ) ;
    NOR2_X1 cell_426 ( .A1 (signal_437), .A2 (signal_370), .ZN (signal_412) ) ;
    NOR2_X1 cell_427 ( .A1 (signal_455), .A2 (signal_438), .ZN (signal_370) ) ;
    MUX2_X1 cell_428 ( .S (signal_925), .A (signal_418), .B (signal_406), .Z (signal_438) ) ;
    INV_X1 cell_429 ( .A (signal_439), .ZN (signal_437) ) ;
    INV_X1 cell_430 ( .A (signal_390), .ZN (signal_436) ) ;
    NAND2_X1 cell_431 ( .A1 (signal_401), .A2 (signal_439), .ZN (signal_1455) ) ;
    NOR2_X1 cell_432 ( .A1 (signal_380), .A2 (signal_391), .ZN (signal_439) ) ;
    NOR2_X1 cell_433 ( .A1 (signal_455), .A2 (signal_440), .ZN (signal_391) ) ;
    MUX2_X1 cell_434 ( .S (signal_925), .A (signal_410), .B (signal_409), .Z (signal_440) ) ;
    NAND2_X1 cell_435 ( .A1 (signal_441), .A2 (signal_442), .ZN (signal_409) ) ;
    NAND2_X1 cell_436 ( .A1 (signal_443), .A2 (signal_926), .ZN (signal_410) ) ;
    NOR2_X1 cell_437 ( .A1 (signal_455), .A2 (signal_444), .ZN (signal_380) ) ;
    MUX2_X1 cell_438 ( .S (signal_925), .A (signal_417), .B (signal_407), .Z (signal_444) ) ;
    NAND2_X1 cell_439 ( .A1 (enc_dec), .A2 (signal_431), .ZN (signal_407) ) ;
    NOR2_X1 cell_440 ( .A1 (signal_924), .A2 (signal_442), .ZN (signal_431) ) ;
    NAND2_X1 cell_441 ( .A1 (signal_445), .A2 (signal_442), .ZN (signal_417) ) ;
    NOR2_X1 cell_442 ( .A1 (signal_399), .A2 (signal_446), .ZN (signal_401) ) ;
    NAND2_X1 cell_443 ( .A1 (signal_374), .A2 (signal_367), .ZN (signal_446) ) ;
    NAND2_X1 cell_444 ( .A1 (signal_420), .A2 (signal_447), .ZN (signal_367) ) ;
    OR2_X1 cell_445 ( .A1 (signal_443), .A2 (signal_441), .ZN (signal_447) ) ;
    AND2_X1 cell_446 ( .A1 (signal_926), .A2 (signal_404), .ZN (signal_420) ) ;
    NOR2_X1 cell_447 ( .A1 (signal_454), .A2 (signal_925), .ZN (signal_404) ) ;
    NOR2_X1 cell_448 ( .A1 (signal_390), .A2 (signal_422), .ZN (signal_374) ) ;
    NOR2_X1 cell_449 ( .A1 (signal_455), .A2 (signal_448), .ZN (signal_422) ) ;
    MUX2_X1 cell_450 ( .S (signal_925), .A (signal_406), .B (signal_418), .Z (signal_448) ) ;
    NAND2_X1 cell_451 ( .A1 (enc_dec), .A2 (signal_449), .ZN (signal_418) ) ;
    NOR2_X1 cell_452 ( .A1 (signal_924), .A2 (signal_926), .ZN (signal_449) ) ;
    NAND2_X1 cell_453 ( .A1 (signal_926), .A2 (signal_445), .ZN (signal_406) ) ;
    NOR2_X1 cell_454 ( .A1 (enc_dec), .A2 (signal_450), .ZN (signal_445) ) ;
    INV_X1 cell_455 ( .A (signal_924), .ZN (signal_450) ) ;
    NOR2_X1 cell_456 ( .A1 (signal_455), .A2 (signal_451), .ZN (signal_390) ) ;
    MUX2_X1 cell_457 ( .S (signal_925), .A (signal_430), .B (signal_452), .Z (signal_451) ) ;
    NOR2_X1 cell_458 ( .A1 (signal_455), .A2 (signal_453), .ZN (signal_399) ) ;
    MUX2_X1 cell_459 ( .S (signal_925), .A (signal_452), .B (signal_430), .Z (signal_453) ) ;
    NAND2_X1 cell_460 ( .A1 (signal_443), .A2 (signal_442), .ZN (signal_430) ) ;
    INV_X1 cell_461 ( .A (signal_926), .ZN (signal_442) ) ;
    NOR2_X1 cell_462 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_443) ) ;
    NAND2_X1 cell_463 ( .A1 (signal_441), .A2 (signal_926), .ZN (signal_452) ) ;
    AND2_X1 cell_464 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_441) ) ;
    INV_X1 cell_465 ( .A (signal_454), .ZN (signal_455) ) ;
    INV_X1 cell_466 ( .A (signal_927), .ZN (signal_454) ) ;
    INV_X1 cell_467 ( .A (signal_927), .ZN (signal_456) ) ;
    INV_X1 cell_468 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_469 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_470 ( .A (signal_456), .ZN (signal_457) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_471 ( .s (signal_927), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1815, signal_302}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_472 ( .s (signal_927), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1816, signal_303}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_473 ( .s (signal_927), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1817, signal_304}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_474 ( .s (signal_927), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1818, signal_305}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_475 ( .s (signal_927), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1819, signal_306}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_476 ( .s (signal_459), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_2139, signal_307}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_477 ( .s (signal_457), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_2140, signal_308}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_478 ( .s (signal_458), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_2141, signal_309}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_479 ( .s (signal_927), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1820, signal_310}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_480 ( .s (signal_927), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1821, signal_311}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_481 ( .s (signal_927), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1822, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_482 ( .s (signal_927), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1823, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_483 ( .s (signal_458), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_2142, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_484 ( .s (signal_927), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1824, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_485 ( .s (signal_927), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1825, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_486 ( .s (signal_927), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1826, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_487 ( .s (signal_457), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_2143, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_488 ( .s (signal_459), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_2144, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_489 ( .s (signal_457), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_2145, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_490 ( .s (signal_457), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_2146, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_491 ( .s (signal_457), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_2147, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_492 ( .s (signal_457), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_2148, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_493 ( .s (signal_458), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_2149, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_494 ( .s (signal_459), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_2150, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_495 ( .s (signal_457), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_2151, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_496 ( .s (signal_458), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_2152, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_497 ( .s (signal_927), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1827, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_498 ( .s (signal_457), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_2153, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_499 ( .s (signal_457), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_2154, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_500 ( .s (signal_457), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_2155, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_501 ( .s (signal_457), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_2156, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_502 ( .s (signal_457), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_2157, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_503 ( .s (signal_457), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_2158, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_504 ( .s (signal_457), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_2159, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_505 ( .s (signal_457), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_2160, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_506 ( .s (signal_457), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_2161, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_507 ( .s (signal_457), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_2162, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_508 ( .s (signal_457), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_2163, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_509 ( .s (signal_457), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_2164, signal_340}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_510 ( .s (signal_457), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_2165, signal_341}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_511 ( .s (signal_458), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_2166, signal_342}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_512 ( .s (signal_458), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_2167, signal_343}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_513 ( .s (signal_458), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_2168, signal_344}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_514 ( .s (signal_458), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_2169, signal_345}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_515 ( .s (signal_458), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_2170, signal_346}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_516 ( .s (signal_458), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_2171, signal_347}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_517 ( .s (signal_458), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_2172, signal_348}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_518 ( .s (signal_458), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_2173, signal_349}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_519 ( .s (signal_458), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_2174, signal_350}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_520 ( .s (signal_458), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_2175, signal_351}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_521 ( .s (signal_458), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_2176, signal_352}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_522 ( .s (signal_458), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_2177, signal_353}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_523 ( .s (signal_459), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_2178, signal_354}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_524 ( .s (signal_459), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_2179, signal_355}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_525 ( .s (signal_459), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_2180, signal_356}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_526 ( .s (signal_459), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_2181, signal_357}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_527 ( .s (signal_459), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_2182, signal_358}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_528 ( .s (signal_459), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_2183, signal_359}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_529 ( .s (signal_459), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_2184, signal_360}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_530 ( .s (signal_459), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_2185, signal_361}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_531 ( .s (signal_459), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_2186, signal_362}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_532 ( .s (signal_459), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_2187, signal_363}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_533 ( .s (signal_459), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_2188, signal_364}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_534 ( .s (signal_459), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_2189, signal_365}) ) ;

    /* cells in depth 1 */
    buf_clk cell_1550 ( .C (clk), .D (signal_265), .Q (signal_3093) ) ;
    buf_clk cell_1622 ( .C (clk), .D (signal_1341), .Q (signal_3165) ) ;
    buf_clk cell_1624 ( .C (clk), .D (signal_2018), .Q (signal_3167) ) ;
    buf_clk cell_1626 ( .C (clk), .D (signal_1372), .Q (signal_3169) ) ;
    buf_clk cell_1628 ( .C (clk), .D (signal_1846), .Q (signal_3171) ) ;
    buf_clk cell_1630 ( .C (clk), .D (signal_1368), .Q (signal_3173) ) ;
    buf_clk cell_1632 ( .C (clk), .D (signal_1828), .Q (signal_3175) ) ;
    buf_clk cell_1634 ( .C (clk), .D (signal_1325), .Q (signal_3177) ) ;
    buf_clk cell_1636 ( .C (clk), .D (signal_2022), .Q (signal_3179) ) ;
    buf_clk cell_1638 ( .C (clk), .D (signal_1323), .Q (signal_3181) ) ;
    buf_clk cell_1640 ( .C (clk), .D (signal_2024), .Q (signal_3183) ) ;
    buf_clk cell_1642 ( .C (clk), .D (signal_1313), .Q (signal_3185) ) ;
    buf_clk cell_1644 ( .C (clk), .D (signal_2026), .Q (signal_3187) ) ;
    buf_clk cell_1646 ( .C (clk), .D (signal_1321), .Q (signal_3189) ) ;
    buf_clk cell_1648 ( .C (clk), .D (signal_2030), .Q (signal_3191) ) ;
    buf_clk cell_1650 ( .C (clk), .D (signal_1364), .Q (signal_3193) ) ;
    buf_clk cell_1652 ( .C (clk), .D (signal_1888), .Q (signal_3195) ) ;
    buf_clk cell_1654 ( .C (clk), .D (signal_1333), .Q (signal_3197) ) ;
    buf_clk cell_1656 ( .C (clk), .D (signal_2033), .Q (signal_3199) ) ;
    buf_clk cell_1658 ( .C (clk), .D (signal_1337), .Q (signal_3201) ) ;
    buf_clk cell_1660 ( .C (clk), .D (signal_2035), .Q (signal_3203) ) ;
    buf_clk cell_1662 ( .C (clk), .D (signal_1317), .Q (signal_3205) ) ;
    buf_clk cell_1664 ( .C (clk), .D (signal_2038), .Q (signal_3207) ) ;
    buf_clk cell_1666 ( .C (clk), .D (signal_1331), .Q (signal_3209) ) ;
    buf_clk cell_1668 ( .C (clk), .D (signal_2043), .Q (signal_3211) ) ;
    buf_clk cell_1670 ( .C (clk), .D (signal_1319), .Q (signal_3213) ) ;
    buf_clk cell_1672 ( .C (clk), .D (signal_2045), .Q (signal_3215) ) ;
    buf_clk cell_1674 ( .C (clk), .D (signal_1375), .Q (signal_3217) ) ;
    buf_clk cell_1676 ( .C (clk), .D (signal_2052), .Q (signal_3219) ) ;
    buf_clk cell_1678 ( .C (clk), .D (signal_1339), .Q (signal_3221) ) ;
    buf_clk cell_1680 ( .C (clk), .D (signal_2056), .Q (signal_3223) ) ;
    buf_clk cell_1682 ( .C (clk), .D (signal_1329), .Q (signal_3225) ) ;
    buf_clk cell_1684 ( .C (clk), .D (signal_2059), .Q (signal_3227) ) ;
    buf_clk cell_1686 ( .C (clk), .D (signal_1335), .Q (signal_3229) ) ;
    buf_clk cell_1688 ( .C (clk), .D (signal_2064), .Q (signal_3231) ) ;
    buf_clk cell_1690 ( .C (clk), .D (signal_1347), .Q (signal_3233) ) ;
    buf_clk cell_1692 ( .C (clk), .D (signal_2067), .Q (signal_3235) ) ;
    buf_clk cell_1694 ( .C (clk), .D (signal_1343), .Q (signal_3237) ) ;
    buf_clk cell_1696 ( .C (clk), .D (signal_2070), .Q (signal_3239) ) ;
    buf_clk cell_1698 ( .C (clk), .D (signal_1371), .Q (signal_3241) ) ;
    buf_clk cell_1700 ( .C (clk), .D (signal_2072), .Q (signal_3243) ) ;
    buf_clk cell_1702 ( .C (clk), .D (signal_1315), .Q (signal_3245) ) ;
    buf_clk cell_1704 ( .C (clk), .D (signal_2075), .Q (signal_3247) ) ;
    buf_clk cell_1706 ( .C (clk), .D (signal_1327), .Q (signal_3249) ) ;
    buf_clk cell_1708 ( .C (clk), .D (signal_2094), .Q (signal_3251) ) ;
    buf_clk cell_1710 ( .C (clk), .D (signal_1345), .Q (signal_3253) ) ;
    buf_clk cell_1712 ( .C (clk), .D (signal_2098), .Q (signal_3255) ) ;
    buf_clk cell_1714 ( .C (clk), .D (signal_1351), .Q (signal_3257) ) ;
    buf_clk cell_1716 ( .C (clk), .D (signal_2106), .Q (signal_3259) ) ;
    buf_clk cell_1718 ( .C (clk), .D (signal_1348), .Q (signal_3261) ) ;
    buf_clk cell_1720 ( .C (clk), .D (signal_1870), .Q (signal_3263) ) ;
    buf_clk cell_1722 ( .C (clk), .D (signal_1355), .Q (signal_3265) ) ;
    buf_clk cell_1724 ( .C (clk), .D (signal_2113), .Q (signal_3267) ) ;
    buf_clk cell_1726 ( .C (clk), .D (signal_1352), .Q (signal_3269) ) ;
    buf_clk cell_1728 ( .C (clk), .D (signal_1875), .Q (signal_3271) ) ;
    buf_clk cell_1730 ( .C (clk), .D (signal_1359), .Q (signal_3273) ) ;
    buf_clk cell_1732 ( .C (clk), .D (signal_2121), .Q (signal_3275) ) ;
    buf_clk cell_1734 ( .C (clk), .D (signal_1356), .Q (signal_3277) ) ;
    buf_clk cell_1736 ( .C (clk), .D (signal_1880), .Q (signal_3279) ) ;
    buf_clk cell_1738 ( .C (clk), .D (signal_1363), .Q (signal_3281) ) ;
    buf_clk cell_1740 ( .C (clk), .D (signal_2128), .Q (signal_3283) ) ;
    buf_clk cell_1742 ( .C (clk), .D (signal_1360), .Q (signal_3285) ) ;
    buf_clk cell_1744 ( .C (clk), .D (signal_1885), .Q (signal_3287) ) ;
    buf_clk cell_1746 ( .C (clk), .D (signal_1367), .Q (signal_3289) ) ;
    buf_clk cell_1748 ( .C (clk), .D (signal_2135), .Q (signal_3291) ) ;
    buf_clk cell_1750 ( .C (clk), .D (signal_914), .Q (signal_3293) ) ;
    buf_clk cell_1756 ( .C (clk), .D (signal_1625), .Q (signal_3299) ) ;
    buf_clk cell_1762 ( .C (clk), .D (signal_916), .Q (signal_3305) ) ;
    buf_clk cell_1768 ( .C (clk), .D (signal_1631), .Q (signal_3311) ) ;
    buf_clk cell_1774 ( .C (clk), .D (signal_860), .Q (signal_3317) ) ;
    buf_clk cell_1780 ( .C (clk), .D (signal_1637), .Q (signal_3323) ) ;
    buf_clk cell_1786 ( .C (clk), .D (signal_862), .Q (signal_3329) ) ;
    buf_clk cell_1792 ( .C (clk), .D (signal_1643), .Q (signal_3335) ) ;
    buf_clk cell_1798 ( .C (clk), .D (signal_918), .Q (signal_3341) ) ;
    buf_clk cell_1804 ( .C (clk), .D (signal_1649), .Q (signal_3347) ) ;
    buf_clk cell_1810 ( .C (clk), .D (signal_864), .Q (signal_3353) ) ;
    buf_clk cell_1816 ( .C (clk), .D (signal_1652), .Q (signal_3359) ) ;
    buf_clk cell_1822 ( .C (clk), .D (signal_866), .Q (signal_3365) ) ;
    buf_clk cell_1828 ( .C (clk), .D (signal_1658), .Q (signal_3371) ) ;
    buf_clk cell_1834 ( .C (clk), .D (signal_868), .Q (signal_3377) ) ;
    buf_clk cell_1840 ( .C (clk), .D (signal_1664), .Q (signal_3383) ) ;
    buf_clk cell_1846 ( .C (clk), .D (signal_870), .Q (signal_3389) ) ;
    buf_clk cell_1852 ( .C (clk), .D (signal_1670), .Q (signal_3395) ) ;
    buf_clk cell_1858 ( .C (clk), .D (signal_872), .Q (signal_3401) ) ;
    buf_clk cell_1864 ( .C (clk), .D (signal_1676), .Q (signal_3407) ) ;
    buf_clk cell_1870 ( .C (clk), .D (signal_874), .Q (signal_3413) ) ;
    buf_clk cell_1876 ( .C (clk), .D (signal_1685), .Q (signal_3419) ) ;
    buf_clk cell_1882 ( .C (clk), .D (signal_876), .Q (signal_3425) ) ;
    buf_clk cell_1888 ( .C (clk), .D (signal_1691), .Q (signal_3431) ) ;
    buf_clk cell_1894 ( .C (clk), .D (signal_878), .Q (signal_3437) ) ;
    buf_clk cell_1900 ( .C (clk), .D (signal_1697), .Q (signal_3443) ) ;
    buf_clk cell_1906 ( .C (clk), .D (signal_880), .Q (signal_3449) ) ;
    buf_clk cell_1912 ( .C (clk), .D (signal_1703), .Q (signal_3455) ) ;
    buf_clk cell_1918 ( .C (clk), .D (signal_882), .Q (signal_3461) ) ;
    buf_clk cell_1924 ( .C (clk), .D (signal_1709), .Q (signal_3467) ) ;
    buf_clk cell_1930 ( .C (clk), .D (signal_920), .Q (signal_3473) ) ;
    buf_clk cell_1936 ( .C (clk), .D (signal_1715), .Q (signal_3479) ) ;
    buf_clk cell_1942 ( .C (clk), .D (signal_884), .Q (signal_3485) ) ;
    buf_clk cell_1948 ( .C (clk), .D (signal_1718), .Q (signal_3491) ) ;
    buf_clk cell_1954 ( .C (clk), .D (signal_886), .Q (signal_3497) ) ;
    buf_clk cell_1960 ( .C (clk), .D (signal_1724), .Q (signal_3503) ) ;
    buf_clk cell_1966 ( .C (clk), .D (signal_888), .Q (signal_3509) ) ;
    buf_clk cell_1972 ( .C (clk), .D (signal_1730), .Q (signal_3515) ) ;
    buf_clk cell_1978 ( .C (clk), .D (signal_890), .Q (signal_3521) ) ;
    buf_clk cell_1984 ( .C (clk), .D (signal_1736), .Q (signal_3527) ) ;
    buf_clk cell_1990 ( .C (clk), .D (signal_892), .Q (signal_3533) ) ;
    buf_clk cell_1996 ( .C (clk), .D (signal_1742), .Q (signal_3539) ) ;
    buf_clk cell_2002 ( .C (clk), .D (signal_894), .Q (signal_3545) ) ;
    buf_clk cell_2008 ( .C (clk), .D (signal_1751), .Q (signal_3551) ) ;
    buf_clk cell_2014 ( .C (clk), .D (signal_896), .Q (signal_3557) ) ;
    buf_clk cell_2020 ( .C (clk), .D (signal_1757), .Q (signal_3563) ) ;
    buf_clk cell_2026 ( .C (clk), .D (signal_898), .Q (signal_3569) ) ;
    buf_clk cell_2032 ( .C (clk), .D (signal_1763), .Q (signal_3575) ) ;
    buf_clk cell_2038 ( .C (clk), .D (signal_900), .Q (signal_3581) ) ;
    buf_clk cell_2044 ( .C (clk), .D (signal_1769), .Q (signal_3587) ) ;
    buf_clk cell_2050 ( .C (clk), .D (signal_902), .Q (signal_3593) ) ;
    buf_clk cell_2056 ( .C (clk), .D (signal_1775), .Q (signal_3599) ) ;
    buf_clk cell_2062 ( .C (clk), .D (signal_922), .Q (signal_3605) ) ;
    buf_clk cell_2068 ( .C (clk), .D (signal_1781), .Q (signal_3611) ) ;
    buf_clk cell_2074 ( .C (clk), .D (signal_904), .Q (signal_3617) ) ;
    buf_clk cell_2080 ( .C (clk), .D (signal_1784), .Q (signal_3623) ) ;
    buf_clk cell_2086 ( .C (clk), .D (signal_906), .Q (signal_3629) ) ;
    buf_clk cell_2092 ( .C (clk), .D (signal_1790), .Q (signal_3635) ) ;
    buf_clk cell_2098 ( .C (clk), .D (signal_908), .Q (signal_3641) ) ;
    buf_clk cell_2104 ( .C (clk), .D (signal_1796), .Q (signal_3647) ) ;
    buf_clk cell_2110 ( .C (clk), .D (signal_910), .Q (signal_3653) ) ;
    buf_clk cell_2116 ( .C (clk), .D (signal_1802), .Q (signal_3659) ) ;
    buf_clk cell_2122 ( .C (clk), .D (signal_912), .Q (signal_3665) ) ;
    buf_clk cell_2128 ( .C (clk), .D (signal_1808), .Q (signal_3671) ) ;
    buf_clk cell_2134 ( .C (clk), .D (signal_311), .Q (signal_3677) ) ;
    buf_clk cell_2140 ( .C (clk), .D (signal_1821), .Q (signal_3683) ) ;
    buf_clk cell_2146 ( .C (clk), .D (signal_309), .Q (signal_3689) ) ;
    buf_clk cell_2152 ( .C (clk), .D (signal_2141), .Q (signal_3695) ) ;
    buf_clk cell_2158 ( .C (clk), .D (signal_365), .Q (signal_3701) ) ;
    buf_clk cell_2164 ( .C (clk), .D (signal_2189), .Q (signal_3707) ) ;
    buf_clk cell_2170 ( .C (clk), .D (signal_363), .Q (signal_3713) ) ;
    buf_clk cell_2176 ( .C (clk), .D (signal_2187), .Q (signal_3719) ) ;
    buf_clk cell_2182 ( .C (clk), .D (signal_307), .Q (signal_3725) ) ;
    buf_clk cell_2188 ( .C (clk), .D (signal_2139), .Q (signal_3731) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_361), .Q (signal_3737) ) ;
    buf_clk cell_2200 ( .C (clk), .D (signal_2185), .Q (signal_3743) ) ;
    buf_clk cell_2206 ( .C (clk), .D (signal_359), .Q (signal_3749) ) ;
    buf_clk cell_2212 ( .C (clk), .D (signal_2183), .Q (signal_3755) ) ;
    buf_clk cell_2218 ( .C (clk), .D (signal_357), .Q (signal_3761) ) ;
    buf_clk cell_2224 ( .C (clk), .D (signal_2181), .Q (signal_3767) ) ;
    buf_clk cell_2230 ( .C (clk), .D (signal_355), .Q (signal_3773) ) ;
    buf_clk cell_2236 ( .C (clk), .D (signal_2179), .Q (signal_3779) ) ;
    buf_clk cell_2242 ( .C (clk), .D (signal_353), .Q (signal_3785) ) ;
    buf_clk cell_2248 ( .C (clk), .D (signal_2177), .Q (signal_3791) ) ;
    buf_clk cell_2254 ( .C (clk), .D (signal_351), .Q (signal_3797) ) ;
    buf_clk cell_2260 ( .C (clk), .D (signal_2175), .Q (signal_3803) ) ;
    buf_clk cell_2266 ( .C (clk), .D (signal_349), .Q (signal_3809) ) ;
    buf_clk cell_2272 ( .C (clk), .D (signal_2173), .Q (signal_3815) ) ;
    buf_clk cell_2278 ( .C (clk), .D (signal_347), .Q (signal_3821) ) ;
    buf_clk cell_2284 ( .C (clk), .D (signal_2171), .Q (signal_3827) ) ;
    buf_clk cell_2290 ( .C (clk), .D (signal_345), .Q (signal_3833) ) ;
    buf_clk cell_2296 ( .C (clk), .D (signal_2169), .Q (signal_3839) ) ;
    buf_clk cell_2302 ( .C (clk), .D (signal_343), .Q (signal_3845) ) ;
    buf_clk cell_2308 ( .C (clk), .D (signal_2167), .Q (signal_3851) ) ;
    buf_clk cell_2314 ( .C (clk), .D (signal_305), .Q (signal_3857) ) ;
    buf_clk cell_2320 ( .C (clk), .D (signal_1818), .Q (signal_3863) ) ;
    buf_clk cell_2326 ( .C (clk), .D (signal_341), .Q (signal_3869) ) ;
    buf_clk cell_2332 ( .C (clk), .D (signal_2165), .Q (signal_3875) ) ;
    buf_clk cell_2338 ( .C (clk), .D (signal_339), .Q (signal_3881) ) ;
    buf_clk cell_2344 ( .C (clk), .D (signal_2163), .Q (signal_3887) ) ;
    buf_clk cell_2350 ( .C (clk), .D (signal_337), .Q (signal_3893) ) ;
    buf_clk cell_2356 ( .C (clk), .D (signal_2161), .Q (signal_3899) ) ;
    buf_clk cell_2362 ( .C (clk), .D (signal_335), .Q (signal_3905) ) ;
    buf_clk cell_2368 ( .C (clk), .D (signal_2159), .Q (signal_3911) ) ;
    buf_clk cell_2374 ( .C (clk), .D (signal_333), .Q (signal_3917) ) ;
    buf_clk cell_2380 ( .C (clk), .D (signal_2157), .Q (signal_3923) ) ;
    buf_clk cell_2386 ( .C (clk), .D (signal_331), .Q (signal_3929) ) ;
    buf_clk cell_2392 ( .C (clk), .D (signal_2155), .Q (signal_3935) ) ;
    buf_clk cell_2398 ( .C (clk), .D (signal_329), .Q (signal_3941) ) ;
    buf_clk cell_2404 ( .C (clk), .D (signal_2153), .Q (signal_3947) ) ;
    buf_clk cell_2410 ( .C (clk), .D (signal_327), .Q (signal_3953) ) ;
    buf_clk cell_2416 ( .C (clk), .D (signal_2152), .Q (signal_3959) ) ;
    buf_clk cell_2422 ( .C (clk), .D (signal_325), .Q (signal_3965) ) ;
    buf_clk cell_2428 ( .C (clk), .D (signal_2150), .Q (signal_3971) ) ;
    buf_clk cell_2434 ( .C (clk), .D (signal_323), .Q (signal_3977) ) ;
    buf_clk cell_2440 ( .C (clk), .D (signal_2148), .Q (signal_3983) ) ;
    buf_clk cell_2446 ( .C (clk), .D (signal_303), .Q (signal_3989) ) ;
    buf_clk cell_2452 ( .C (clk), .D (signal_1816), .Q (signal_3995) ) ;
    buf_clk cell_2458 ( .C (clk), .D (signal_321), .Q (signal_4001) ) ;
    buf_clk cell_2464 ( .C (clk), .D (signal_2146), .Q (signal_4007) ) ;
    buf_clk cell_2470 ( .C (clk), .D (signal_319), .Q (signal_4013) ) ;
    buf_clk cell_2476 ( .C (clk), .D (signal_2144), .Q (signal_4019) ) ;
    buf_clk cell_2482 ( .C (clk), .D (signal_317), .Q (signal_4025) ) ;
    buf_clk cell_2488 ( .C (clk), .D (signal_1826), .Q (signal_4031) ) ;
    buf_clk cell_2494 ( .C (clk), .D (signal_315), .Q (signal_4037) ) ;
    buf_clk cell_2500 ( .C (clk), .D (signal_1824), .Q (signal_4043) ) ;
    buf_clk cell_2506 ( .C (clk), .D (signal_313), .Q (signal_4049) ) ;
    buf_clk cell_2512 ( .C (clk), .D (signal_1823), .Q (signal_4055) ) ;
    buf_clk cell_2518 ( .C (clk), .D (reset), .Q (signal_4061) ) ;
    buf_clk cell_2524 ( .C (clk), .D (signal_990), .Q (signal_4067) ) ;
    buf_clk cell_2530 ( .C (clk), .D (signal_1995), .Q (signal_4073) ) ;
    buf_clk cell_2536 ( .C (clk), .D (signal_988), .Q (signal_4079) ) ;
    buf_clk cell_2542 ( .C (clk), .D (signal_1951), .Q (signal_4085) ) ;
    buf_clk cell_2548 ( .C (clk), .D (signal_986), .Q (signal_4091) ) ;
    buf_clk cell_2554 ( .C (clk), .D (signal_1907), .Q (signal_4097) ) ;
    buf_clk cell_2560 ( .C (clk), .D (signal_984), .Q (signal_4103) ) ;
    buf_clk cell_2566 ( .C (clk), .D (signal_1895), .Q (signal_4109) ) ;
    buf_clk cell_2572 ( .C (clk), .D (signal_982), .Q (signal_4115) ) ;
    buf_clk cell_2578 ( .C (clk), .D (signal_1891), .Q (signal_4121) ) ;
    buf_clk cell_2584 ( .C (clk), .D (signal_980), .Q (signal_4127) ) ;
    buf_clk cell_2590 ( .C (clk), .D (signal_2013), .Q (signal_4133) ) ;
    buf_clk cell_2596 ( .C (clk), .D (signal_978), .Q (signal_4139) ) ;
    buf_clk cell_2602 ( .C (clk), .D (signal_2009), .Q (signal_4145) ) ;
    buf_clk cell_2608 ( .C (clk), .D (signal_976), .Q (signal_4151) ) ;
    buf_clk cell_2614 ( .C (clk), .D (signal_2005), .Q (signal_4157) ) ;
    buf_clk cell_2620 ( .C (clk), .D (signal_974), .Q (signal_4163) ) ;
    buf_clk cell_2626 ( .C (clk), .D (signal_2001), .Q (signal_4169) ) ;
    buf_clk cell_2632 ( .C (clk), .D (signal_972), .Q (signal_4175) ) ;
    buf_clk cell_2638 ( .C (clk), .D (signal_1997), .Q (signal_4181) ) ;
    buf_clk cell_2644 ( .C (clk), .D (signal_970), .Q (signal_4187) ) ;
    buf_clk cell_2650 ( .C (clk), .D (signal_1991), .Q (signal_4193) ) ;
    buf_clk cell_2656 ( .C (clk), .D (signal_968), .Q (signal_4199) ) ;
    buf_clk cell_2662 ( .C (clk), .D (signal_1987), .Q (signal_4205) ) ;
    buf_clk cell_2668 ( .C (clk), .D (signal_966), .Q (signal_4211) ) ;
    buf_clk cell_2674 ( .C (clk), .D (signal_1983), .Q (signal_4217) ) ;
    buf_clk cell_2680 ( .C (clk), .D (signal_964), .Q (signal_4223) ) ;
    buf_clk cell_2686 ( .C (clk), .D (signal_1979), .Q (signal_4229) ) ;
    buf_clk cell_2692 ( .C (clk), .D (signal_962), .Q (signal_4235) ) ;
    buf_clk cell_2698 ( .C (clk), .D (signal_1975), .Q (signal_4241) ) ;
    buf_clk cell_2704 ( .C (clk), .D (signal_960), .Q (signal_4247) ) ;
    buf_clk cell_2710 ( .C (clk), .D (signal_1969), .Q (signal_4253) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_958), .Q (signal_4259) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_1965), .Q (signal_4265) ) ;
    buf_clk cell_2728 ( .C (clk), .D (signal_956), .Q (signal_4271) ) ;
    buf_clk cell_2734 ( .C (clk), .D (signal_1961), .Q (signal_4277) ) ;
    buf_clk cell_2740 ( .C (clk), .D (signal_954), .Q (signal_4283) ) ;
    buf_clk cell_2746 ( .C (clk), .D (signal_1957), .Q (signal_4289) ) ;
    buf_clk cell_2752 ( .C (clk), .D (signal_952), .Q (signal_4295) ) ;
    buf_clk cell_2758 ( .C (clk), .D (signal_1953), .Q (signal_4301) ) ;
    buf_clk cell_2764 ( .C (clk), .D (signal_950), .Q (signal_4307) ) ;
    buf_clk cell_2770 ( .C (clk), .D (signal_1947), .Q (signal_4313) ) ;
    buf_clk cell_2776 ( .C (clk), .D (signal_948), .Q (signal_4319) ) ;
    buf_clk cell_2782 ( .C (clk), .D (signal_1943), .Q (signal_4325) ) ;
    buf_clk cell_2788 ( .C (clk), .D (signal_946), .Q (signal_4331) ) ;
    buf_clk cell_2794 ( .C (clk), .D (signal_1939), .Q (signal_4337) ) ;
    buf_clk cell_2800 ( .C (clk), .D (signal_944), .Q (signal_4343) ) ;
    buf_clk cell_2806 ( .C (clk), .D (signal_1935), .Q (signal_4349) ) ;
    buf_clk cell_2812 ( .C (clk), .D (signal_942), .Q (signal_4355) ) ;
    buf_clk cell_2818 ( .C (clk), .D (signal_1931), .Q (signal_4361) ) ;
    buf_clk cell_2824 ( .C (clk), .D (signal_940), .Q (signal_4367) ) ;
    buf_clk cell_2830 ( .C (clk), .D (signal_1925), .Q (signal_4373) ) ;
    buf_clk cell_2836 ( .C (clk), .D (signal_938), .Q (signal_4379) ) ;
    buf_clk cell_2842 ( .C (clk), .D (signal_1921), .Q (signal_4385) ) ;
    buf_clk cell_2848 ( .C (clk), .D (signal_936), .Q (signal_4391) ) ;
    buf_clk cell_2854 ( .C (clk), .D (signal_1917), .Q (signal_4397) ) ;
    buf_clk cell_2860 ( .C (clk), .D (signal_934), .Q (signal_4403) ) ;
    buf_clk cell_2866 ( .C (clk), .D (signal_1913), .Q (signal_4409) ) ;
    buf_clk cell_2872 ( .C (clk), .D (signal_932), .Q (signal_4415) ) ;
    buf_clk cell_2878 ( .C (clk), .D (signal_1909), .Q (signal_4421) ) ;
    buf_clk cell_2884 ( .C (clk), .D (signal_930), .Q (signal_4427) ) ;
    buf_clk cell_2890 ( .C (clk), .D (signal_1903), .Q (signal_4433) ) ;
    buf_clk cell_2896 ( .C (clk), .D (signal_928), .Q (signal_4439) ) ;
    buf_clk cell_2902 ( .C (clk), .D (signal_1899), .Q (signal_4445) ) ;
    buf_clk cell_2908 ( .C (clk), .D (enc_dec), .Q (signal_4451) ) ;
    buf_clk cell_2918 ( .C (clk), .D (signal_1334), .Q (signal_4461) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_2191), .Q (signal_4465) ) ;
    buf_clk cell_2954 ( .C (clk), .D (signal_1330), .Q (signal_4497) ) ;
    buf_clk cell_2958 ( .C (clk), .D (signal_2202), .Q (signal_4501) ) ;
    buf_clk cell_2962 ( .C (clk), .D (signal_1326), .Q (signal_4505) ) ;
    buf_clk cell_2966 ( .C (clk), .D (signal_2205), .Q (signal_4509) ) ;
    buf_clk cell_2974 ( .C (clk), .D (signal_1338), .Q (signal_4517) ) ;
    buf_clk cell_2978 ( .C (clk), .D (signal_2211), .Q (signal_4521) ) ;
    buf_clk cell_2982 ( .C (clk), .D (signal_1314), .Q (signal_4525) ) ;
    buf_clk cell_2986 ( .C (clk), .D (signal_2217), .Q (signal_4529) ) ;
    buf_clk cell_2990 ( .C (clk), .D (signal_1342), .Q (signal_4533) ) ;
    buf_clk cell_2994 ( .C (clk), .D (signal_2219), .Q (signal_4537) ) ;
    buf_clk cell_3002 ( .C (clk), .D (signal_1374), .Q (signal_4545) ) ;
    buf_clk cell_3006 ( .C (clk), .D (signal_2224), .Q (signal_4549) ) ;
    buf_clk cell_3010 ( .C (clk), .D (signal_1318), .Q (signal_4553) ) ;
    buf_clk cell_3014 ( .C (clk), .D (signal_2226), .Q (signal_4557) ) ;
    buf_clk cell_3018 ( .C (clk), .D (signal_1322), .Q (signal_4561) ) ;
    buf_clk cell_3022 ( .C (clk), .D (signal_2230), .Q (signal_4565) ) ;
    buf_clk cell_3026 ( .C (clk), .D (signal_1370), .Q (signal_4569) ) ;
    buf_clk cell_3030 ( .C (clk), .D (signal_2233), .Q (signal_4573) ) ;
    buf_clk cell_3034 ( .C (clk), .D (signal_1346), .Q (signal_4577) ) ;
    buf_clk cell_3038 ( .C (clk), .D (signal_2239), .Q (signal_4581) ) ;
    buf_clk cell_3050 ( .C (clk), .D (signal_1350), .Q (signal_4593) ) ;
    buf_clk cell_3054 ( .C (clk), .D (signal_2245), .Q (signal_4597) ) ;
    buf_clk cell_3062 ( .C (clk), .D (signal_1354), .Q (signal_4605) ) ;
    buf_clk cell_3066 ( .C (clk), .D (signal_2250), .Q (signal_4609) ) ;
    buf_clk cell_3074 ( .C (clk), .D (signal_1358), .Q (signal_4617) ) ;
    buf_clk cell_3078 ( .C (clk), .D (signal_2256), .Q (signal_4621) ) ;
    buf_clk cell_3086 ( .C (clk), .D (signal_1362), .Q (signal_4629) ) ;
    buf_clk cell_3090 ( .C (clk), .D (signal_2261), .Q (signal_4633) ) ;
    buf_clk cell_3098 ( .C (clk), .D (signal_1366), .Q (signal_4641) ) ;
    buf_clk cell_3102 ( .C (clk), .D (signal_2266), .Q (signal_4645) ) ;
    buf_clk cell_3106 ( .C (clk), .D (signal_915), .Q (signal_4649) ) ;
    buf_clk cell_3114 ( .C (clk), .D (signal_1628), .Q (signal_4657) ) ;
    buf_clk cell_3122 ( .C (clk), .D (signal_917), .Q (signal_4665) ) ;
    buf_clk cell_3130 ( .C (clk), .D (signal_1634), .Q (signal_4673) ) ;
    buf_clk cell_3138 ( .C (clk), .D (signal_861), .Q (signal_4681) ) ;
    buf_clk cell_3146 ( .C (clk), .D (signal_1640), .Q (signal_4689) ) ;
    buf_clk cell_3154 ( .C (clk), .D (signal_863), .Q (signal_4697) ) ;
    buf_clk cell_3162 ( .C (clk), .D (signal_1646), .Q (signal_4705) ) ;
    buf_clk cell_3170 ( .C (clk), .D (signal_865), .Q (signal_4713) ) ;
    buf_clk cell_3178 ( .C (clk), .D (signal_1655), .Q (signal_4721) ) ;
    buf_clk cell_3186 ( .C (clk), .D (signal_867), .Q (signal_4729) ) ;
    buf_clk cell_3194 ( .C (clk), .D (signal_1661), .Q (signal_4737) ) ;
    buf_clk cell_3202 ( .C (clk), .D (signal_869), .Q (signal_4745) ) ;
    buf_clk cell_3210 ( .C (clk), .D (signal_1667), .Q (signal_4753) ) ;
    buf_clk cell_3218 ( .C (clk), .D (signal_871), .Q (signal_4761) ) ;
    buf_clk cell_3226 ( .C (clk), .D (signal_1673), .Q (signal_4769) ) ;
    buf_clk cell_3234 ( .C (clk), .D (signal_873), .Q (signal_4777) ) ;
    buf_clk cell_3242 ( .C (clk), .D (signal_1679), .Q (signal_4785) ) ;
    buf_clk cell_3250 ( .C (clk), .D (signal_919), .Q (signal_4793) ) ;
    buf_clk cell_3258 ( .C (clk), .D (signal_1682), .Q (signal_4801) ) ;
    buf_clk cell_3266 ( .C (clk), .D (signal_875), .Q (signal_4809) ) ;
    buf_clk cell_3274 ( .C (clk), .D (signal_1688), .Q (signal_4817) ) ;
    buf_clk cell_3282 ( .C (clk), .D (signal_877), .Q (signal_4825) ) ;
    buf_clk cell_3290 ( .C (clk), .D (signal_1694), .Q (signal_4833) ) ;
    buf_clk cell_3298 ( .C (clk), .D (signal_879), .Q (signal_4841) ) ;
    buf_clk cell_3306 ( .C (clk), .D (signal_1700), .Q (signal_4849) ) ;
    buf_clk cell_3314 ( .C (clk), .D (signal_881), .Q (signal_4857) ) ;
    buf_clk cell_3322 ( .C (clk), .D (signal_1706), .Q (signal_4865) ) ;
    buf_clk cell_3330 ( .C (clk), .D (signal_883), .Q (signal_4873) ) ;
    buf_clk cell_3338 ( .C (clk), .D (signal_1712), .Q (signal_4881) ) ;
    buf_clk cell_3346 ( .C (clk), .D (signal_885), .Q (signal_4889) ) ;
    buf_clk cell_3354 ( .C (clk), .D (signal_1721), .Q (signal_4897) ) ;
    buf_clk cell_3362 ( .C (clk), .D (signal_887), .Q (signal_4905) ) ;
    buf_clk cell_3370 ( .C (clk), .D (signal_1727), .Q (signal_4913) ) ;
    buf_clk cell_3378 ( .C (clk), .D (signal_889), .Q (signal_4921) ) ;
    buf_clk cell_3386 ( .C (clk), .D (signal_1733), .Q (signal_4929) ) ;
    buf_clk cell_3394 ( .C (clk), .D (signal_891), .Q (signal_4937) ) ;
    buf_clk cell_3402 ( .C (clk), .D (signal_1739), .Q (signal_4945) ) ;
    buf_clk cell_3410 ( .C (clk), .D (signal_893), .Q (signal_4953) ) ;
    buf_clk cell_3418 ( .C (clk), .D (signal_1745), .Q (signal_4961) ) ;
    buf_clk cell_3426 ( .C (clk), .D (signal_921), .Q (signal_4969) ) ;
    buf_clk cell_3434 ( .C (clk), .D (signal_1748), .Q (signal_4977) ) ;
    buf_clk cell_3442 ( .C (clk), .D (signal_895), .Q (signal_4985) ) ;
    buf_clk cell_3450 ( .C (clk), .D (signal_1754), .Q (signal_4993) ) ;
    buf_clk cell_3458 ( .C (clk), .D (signal_897), .Q (signal_5001) ) ;
    buf_clk cell_3466 ( .C (clk), .D (signal_1760), .Q (signal_5009) ) ;
    buf_clk cell_3474 ( .C (clk), .D (signal_899), .Q (signal_5017) ) ;
    buf_clk cell_3482 ( .C (clk), .D (signal_1766), .Q (signal_5025) ) ;
    buf_clk cell_3490 ( .C (clk), .D (signal_901), .Q (signal_5033) ) ;
    buf_clk cell_3498 ( .C (clk), .D (signal_1772), .Q (signal_5041) ) ;
    buf_clk cell_3506 ( .C (clk), .D (signal_903), .Q (signal_5049) ) ;
    buf_clk cell_3514 ( .C (clk), .D (signal_1778), .Q (signal_5057) ) ;
    buf_clk cell_3522 ( .C (clk), .D (signal_905), .Q (signal_5065) ) ;
    buf_clk cell_3530 ( .C (clk), .D (signal_1787), .Q (signal_5073) ) ;
    buf_clk cell_3538 ( .C (clk), .D (signal_907), .Q (signal_5081) ) ;
    buf_clk cell_3546 ( .C (clk), .D (signal_1793), .Q (signal_5089) ) ;
    buf_clk cell_3554 ( .C (clk), .D (signal_909), .Q (signal_5097) ) ;
    buf_clk cell_3562 ( .C (clk), .D (signal_1799), .Q (signal_5105) ) ;
    buf_clk cell_3570 ( .C (clk), .D (signal_911), .Q (signal_5113) ) ;
    buf_clk cell_3578 ( .C (clk), .D (signal_1805), .Q (signal_5121) ) ;
    buf_clk cell_3586 ( .C (clk), .D (signal_913), .Q (signal_5129) ) ;
    buf_clk cell_3594 ( .C (clk), .D (signal_1811), .Q (signal_5137) ) ;
    buf_clk cell_3602 ( .C (clk), .D (signal_923), .Q (signal_5145) ) ;
    buf_clk cell_3610 ( .C (clk), .D (signal_1814), .Q (signal_5153) ) ;
    buf_clk cell_3618 ( .C (clk), .D (signal_286), .Q (signal_5161) ) ;
    buf_clk cell_3626 ( .C (clk), .D (signal_2566), .Q (signal_5169) ) ;
    buf_clk cell_3634 ( .C (clk), .D (signal_308), .Q (signal_5177) ) ;
    buf_clk cell_3642 ( .C (clk), .D (signal_2140), .Q (signal_5185) ) ;
    buf_clk cell_3650 ( .C (clk), .D (signal_364), .Q (signal_5193) ) ;
    buf_clk cell_3658 ( .C (clk), .D (signal_2188), .Q (signal_5201) ) ;
    buf_clk cell_3666 ( .C (clk), .D (signal_287), .Q (signal_5209) ) ;
    buf_clk cell_3674 ( .C (clk), .D (signal_2622), .Q (signal_5217) ) ;
    buf_clk cell_3682 ( .C (clk), .D (signal_360), .Q (signal_5225) ) ;
    buf_clk cell_3690 ( .C (clk), .D (signal_2184), .Q (signal_5233) ) ;
    buf_clk cell_3698 ( .C (clk), .D (signal_288), .Q (signal_5241) ) ;
    buf_clk cell_3706 ( .C (clk), .D (signal_2623), .Q (signal_5249) ) ;
    buf_clk cell_3714 ( .C (clk), .D (signal_356), .Q (signal_5257) ) ;
    buf_clk cell_3722 ( .C (clk), .D (signal_2180), .Q (signal_5265) ) ;
    buf_clk cell_3730 ( .C (clk), .D (signal_289), .Q (signal_5273) ) ;
    buf_clk cell_3738 ( .C (clk), .D (signal_2624), .Q (signal_5281) ) ;
    buf_clk cell_3746 ( .C (clk), .D (signal_352), .Q (signal_5289) ) ;
    buf_clk cell_3754 ( .C (clk), .D (signal_2176), .Q (signal_5297) ) ;
    buf_clk cell_3762 ( .C (clk), .D (signal_290), .Q (signal_5305) ) ;
    buf_clk cell_3770 ( .C (clk), .D (signal_2625), .Q (signal_5313) ) ;
    buf_clk cell_3778 ( .C (clk), .D (signal_291), .Q (signal_5321) ) ;
    buf_clk cell_3786 ( .C (clk), .D (signal_2712), .Q (signal_5329) ) ;
    buf_clk cell_3794 ( .C (clk), .D (signal_348), .Q (signal_5337) ) ;
    buf_clk cell_3802 ( .C (clk), .D (signal_2172), .Q (signal_5345) ) ;
    buf_clk cell_3810 ( .C (clk), .D (signal_292), .Q (signal_5353) ) ;
    buf_clk cell_3818 ( .C (clk), .D (signal_2573), .Q (signal_5361) ) ;
    buf_clk cell_3826 ( .C (clk), .D (signal_344), .Q (signal_5369) ) ;
    buf_clk cell_3834 ( .C (clk), .D (signal_2168), .Q (signal_5377) ) ;
    buf_clk cell_3842 ( .C (clk), .D (signal_293), .Q (signal_5385) ) ;
    buf_clk cell_3850 ( .C (clk), .D (signal_2626), .Q (signal_5393) ) ;
    buf_clk cell_3858 ( .C (clk), .D (signal_340), .Q (signal_5401) ) ;
    buf_clk cell_3866 ( .C (clk), .D (signal_2164), .Q (signal_5409) ) ;
    buf_clk cell_3874 ( .C (clk), .D (signal_294), .Q (signal_5417) ) ;
    buf_clk cell_3882 ( .C (clk), .D (signal_2576), .Q (signal_5425) ) ;
    buf_clk cell_3890 ( .C (clk), .D (signal_336), .Q (signal_5433) ) ;
    buf_clk cell_3898 ( .C (clk), .D (signal_2160), .Q (signal_5441) ) ;
    buf_clk cell_3906 ( .C (clk), .D (signal_295), .Q (signal_5449) ) ;
    buf_clk cell_3914 ( .C (clk), .D (signal_2627), .Q (signal_5457) ) ;
    buf_clk cell_3922 ( .C (clk), .D (signal_332), .Q (signal_5465) ) ;
    buf_clk cell_3930 ( .C (clk), .D (signal_2156), .Q (signal_5473) ) ;
    buf_clk cell_3938 ( .C (clk), .D (signal_304), .Q (signal_5481) ) ;
    buf_clk cell_3946 ( .C (clk), .D (signal_1817), .Q (signal_5489) ) ;
    buf_clk cell_3954 ( .C (clk), .D (signal_296), .Q (signal_5497) ) ;
    buf_clk cell_3962 ( .C (clk), .D (signal_2690), .Q (signal_5505) ) ;
    buf_clk cell_3970 ( .C (clk), .D (signal_328), .Q (signal_5513) ) ;
    buf_clk cell_3978 ( .C (clk), .D (signal_1827), .Q (signal_5521) ) ;
    buf_clk cell_3986 ( .C (clk), .D (signal_297), .Q (signal_5529) ) ;
    buf_clk cell_3994 ( .C (clk), .D (signal_2628), .Q (signal_5537) ) ;
    buf_clk cell_4002 ( .C (clk), .D (signal_324), .Q (signal_5545) ) ;
    buf_clk cell_4010 ( .C (clk), .D (signal_2149), .Q (signal_5553) ) ;
    buf_clk cell_4018 ( .C (clk), .D (signal_298), .Q (signal_5561) ) ;
    buf_clk cell_4026 ( .C (clk), .D (signal_2582), .Q (signal_5569) ) ;
    buf_clk cell_4034 ( .C (clk), .D (signal_320), .Q (signal_5577) ) ;
    buf_clk cell_4042 ( .C (clk), .D (signal_2145), .Q (signal_5585) ) ;
    buf_clk cell_4050 ( .C (clk), .D (signal_299), .Q (signal_5593) ) ;
    buf_clk cell_4058 ( .C (clk), .D (signal_2629), .Q (signal_5601) ) ;
    buf_clk cell_4066 ( .C (clk), .D (signal_316), .Q (signal_5609) ) ;
    buf_clk cell_4074 ( .C (clk), .D (signal_1825), .Q (signal_5617) ) ;
    buf_clk cell_4082 ( .C (clk), .D (signal_300), .Q (signal_5625) ) ;
    buf_clk cell_4090 ( .C (clk), .D (signal_2630), .Q (signal_5633) ) ;
    buf_clk cell_4098 ( .C (clk), .D (signal_312), .Q (signal_5641) ) ;
    buf_clk cell_4106 ( .C (clk), .D (signal_1822), .Q (signal_5649) ) ;
    buf_clk cell_4114 ( .C (clk), .D (signal_301), .Q (signal_5657) ) ;
    buf_clk cell_4122 ( .C (clk), .D (signal_2631), .Q (signal_5665) ) ;
    buf_clk cell_4132 ( .C (clk), .D (signal_991), .Q (signal_5675) ) ;
    buf_clk cell_4140 ( .C (clk), .D (signal_2017), .Q (signal_5683) ) ;
    buf_clk cell_4148 ( .C (clk), .D (signal_989), .Q (signal_5691) ) ;
    buf_clk cell_4156 ( .C (clk), .D (signal_1973), .Q (signal_5699) ) ;
    buf_clk cell_4164 ( .C (clk), .D (signal_987), .Q (signal_5707) ) ;
    buf_clk cell_4172 ( .C (clk), .D (signal_1929), .Q (signal_5715) ) ;
    buf_clk cell_4180 ( .C (clk), .D (signal_985), .Q (signal_5723) ) ;
    buf_clk cell_4188 ( .C (clk), .D (signal_1897), .Q (signal_5731) ) ;
    buf_clk cell_4196 ( .C (clk), .D (signal_983), .Q (signal_5739) ) ;
    buf_clk cell_4204 ( .C (clk), .D (signal_1893), .Q (signal_5747) ) ;
    buf_clk cell_4212 ( .C (clk), .D (signal_981), .Q (signal_5755) ) ;
    buf_clk cell_4220 ( .C (clk), .D (signal_2015), .Q (signal_5763) ) ;
    buf_clk cell_4228 ( .C (clk), .D (signal_979), .Q (signal_5771) ) ;
    buf_clk cell_4236 ( .C (clk), .D (signal_2011), .Q (signal_5779) ) ;
    buf_clk cell_4244 ( .C (clk), .D (signal_977), .Q (signal_5787) ) ;
    buf_clk cell_4252 ( .C (clk), .D (signal_2007), .Q (signal_5795) ) ;
    buf_clk cell_4260 ( .C (clk), .D (signal_975), .Q (signal_5803) ) ;
    buf_clk cell_4268 ( .C (clk), .D (signal_2003), .Q (signal_5811) ) ;
    buf_clk cell_4276 ( .C (clk), .D (signal_973), .Q (signal_5819) ) ;
    buf_clk cell_4284 ( .C (clk), .D (signal_1999), .Q (signal_5827) ) ;
    buf_clk cell_4292 ( .C (clk), .D (signal_971), .Q (signal_5835) ) ;
    buf_clk cell_4300 ( .C (clk), .D (signal_1993), .Q (signal_5843) ) ;
    buf_clk cell_4308 ( .C (clk), .D (signal_969), .Q (signal_5851) ) ;
    buf_clk cell_4316 ( .C (clk), .D (signal_1989), .Q (signal_5859) ) ;
    buf_clk cell_4324 ( .C (clk), .D (signal_967), .Q (signal_5867) ) ;
    buf_clk cell_4332 ( .C (clk), .D (signal_1985), .Q (signal_5875) ) ;
    buf_clk cell_4340 ( .C (clk), .D (signal_965), .Q (signal_5883) ) ;
    buf_clk cell_4348 ( .C (clk), .D (signal_1981), .Q (signal_5891) ) ;
    buf_clk cell_4356 ( .C (clk), .D (signal_963), .Q (signal_5899) ) ;
    buf_clk cell_4364 ( .C (clk), .D (signal_1977), .Q (signal_5907) ) ;
    buf_clk cell_4372 ( .C (clk), .D (signal_961), .Q (signal_5915) ) ;
    buf_clk cell_4380 ( .C (clk), .D (signal_1971), .Q (signal_5923) ) ;
    buf_clk cell_4388 ( .C (clk), .D (signal_959), .Q (signal_5931) ) ;
    buf_clk cell_4396 ( .C (clk), .D (signal_1967), .Q (signal_5939) ) ;
    buf_clk cell_4404 ( .C (clk), .D (signal_957), .Q (signal_5947) ) ;
    buf_clk cell_4412 ( .C (clk), .D (signal_1963), .Q (signal_5955) ) ;
    buf_clk cell_4420 ( .C (clk), .D (signal_955), .Q (signal_5963) ) ;
    buf_clk cell_4428 ( .C (clk), .D (signal_1959), .Q (signal_5971) ) ;
    buf_clk cell_4436 ( .C (clk), .D (signal_953), .Q (signal_5979) ) ;
    buf_clk cell_4444 ( .C (clk), .D (signal_1955), .Q (signal_5987) ) ;
    buf_clk cell_4452 ( .C (clk), .D (signal_951), .Q (signal_5995) ) ;
    buf_clk cell_4460 ( .C (clk), .D (signal_1949), .Q (signal_6003) ) ;
    buf_clk cell_4468 ( .C (clk), .D (signal_949), .Q (signal_6011) ) ;
    buf_clk cell_4476 ( .C (clk), .D (signal_1945), .Q (signal_6019) ) ;
    buf_clk cell_4484 ( .C (clk), .D (signal_947), .Q (signal_6027) ) ;
    buf_clk cell_4492 ( .C (clk), .D (signal_1941), .Q (signal_6035) ) ;
    buf_clk cell_4500 ( .C (clk), .D (signal_945), .Q (signal_6043) ) ;
    buf_clk cell_4508 ( .C (clk), .D (signal_1937), .Q (signal_6051) ) ;
    buf_clk cell_4516 ( .C (clk), .D (signal_943), .Q (signal_6059) ) ;
    buf_clk cell_4524 ( .C (clk), .D (signal_1933), .Q (signal_6067) ) ;
    buf_clk cell_4532 ( .C (clk), .D (signal_941), .Q (signal_6075) ) ;
    buf_clk cell_4540 ( .C (clk), .D (signal_1927), .Q (signal_6083) ) ;
    buf_clk cell_4548 ( .C (clk), .D (signal_939), .Q (signal_6091) ) ;
    buf_clk cell_4556 ( .C (clk), .D (signal_1923), .Q (signal_6099) ) ;
    buf_clk cell_4564 ( .C (clk), .D (signal_937), .Q (signal_6107) ) ;
    buf_clk cell_4572 ( .C (clk), .D (signal_1919), .Q (signal_6115) ) ;
    buf_clk cell_4580 ( .C (clk), .D (signal_935), .Q (signal_6123) ) ;
    buf_clk cell_4588 ( .C (clk), .D (signal_1915), .Q (signal_6131) ) ;
    buf_clk cell_4596 ( .C (clk), .D (signal_933), .Q (signal_6139) ) ;
    buf_clk cell_4604 ( .C (clk), .D (signal_1911), .Q (signal_6147) ) ;
    buf_clk cell_4612 ( .C (clk), .D (signal_931), .Q (signal_6155) ) ;
    buf_clk cell_4620 ( .C (clk), .D (signal_1905), .Q (signal_6163) ) ;
    buf_clk cell_4628 ( .C (clk), .D (signal_929), .Q (signal_6171) ) ;
    buf_clk cell_4636 ( .C (clk), .D (signal_1901), .Q (signal_6179) ) ;
    buf_clk cell_4838 ( .C (clk), .D (signal_283), .Q (signal_6381) ) ;
    buf_clk cell_4846 ( .C (clk), .D (signal_282), .Q (signal_6389) ) ;
    buf_clk cell_4854 ( .C (clk), .D (signal_278), .Q (signal_6397) ) ;
    buf_clk cell_4862 ( .C (clk), .D (signal_280), .Q (signal_6405) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1255 ( .s ({signal_1828, signal_1368}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_1829, signal_1456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1256 ( .s ({signal_1830, signal_1332}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[1]), .c ({signal_1831, signal_1457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1257 ( .s ({signal_1832, signal_1316}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_1833, signal_1458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1258 ( .s ({signal_1834, signal_1344}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[3]), .c ({signal_1835, signal_1459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1259 ( .s ({signal_1836, signal_1369}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[4]), .c ({signal_1837, signal_1460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1260 ( .s ({signal_1836, signal_1369}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[5]), .c ({signal_1838, signal_1461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1261 ( .s ({signal_1839, signal_1365}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[6]), .c ({signal_1840, signal_1462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1262 ( .s ({signal_1841, signal_1373}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[7]), .c ({signal_1842, signal_1463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1263 ( .s ({signal_1843, signal_1340}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[8]), .c ({signal_1844, signal_1464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1264 ( .s ({signal_1839, signal_1365}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[9]), .c ({signal_1845, signal_1465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1265 ( .s ({signal_1846, signal_1372}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[10]), .c ({signal_1847, signal_1466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1266 ( .s ({signal_1841, signal_1373}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[11]), .c ({signal_1848, signal_1467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1267 ( .s ({signal_1843, signal_1340}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[12]), .c ({signal_1849, signal_1468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1268 ( .s ({signal_1850, signal_1320}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[13]), .c ({signal_1851, signal_1469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1269 ( .s ({signal_1832, signal_1316}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[14]), .c ({signal_1852, signal_1470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1270 ( .s ({signal_1830, signal_1332}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[15]), .c ({signal_1853, signal_1471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1271 ( .s ({signal_1854, signal_1328}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[16]), .c ({signal_1855, signal_1472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1272 ( .s ({signal_1856, signal_1324}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[17]), .c ({signal_1857, signal_1473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1273 ( .s ({signal_1854, signal_1328}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[18]), .c ({signal_1858, signal_1474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1274 ( .s ({signal_1850, signal_1320}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[19]), .c ({signal_1859, signal_1475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1275 ( .s ({signal_1860, signal_1336}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[20]), .c ({signal_1861, signal_1476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1276 ( .s ({signal_1862, signal_1312}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[21]), .c ({signal_1863, signal_1477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1277 ( .s ({signal_1834, signal_1344}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[22]), .c ({signal_1864, signal_1478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1278 ( .s ({signal_1856, signal_1324}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[23]), .c ({signal_1865, signal_1479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1279 ( .s ({signal_1860, signal_1336}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[24]), .c ({signal_1866, signal_1480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1280 ( .s ({signal_1862, signal_1312}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[25]), .c ({signal_1867, signal_1481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1281 ( .s ({signal_1868, signal_1349}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[26]), .c ({signal_1869, signal_1482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1282 ( .s ({signal_1870, signal_1348}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[27]), .c ({signal_1871, signal_1483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1283 ( .s ({signal_1868, signal_1349}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[28]), .c ({signal_1872, signal_1484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1284 ( .s ({signal_1873, signal_1353}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[29]), .c ({signal_1874, signal_1485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1285 ( .s ({signal_1875, signal_1352}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[30]), .c ({signal_1876, signal_1486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1286 ( .s ({signal_1873, signal_1353}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[31]), .c ({signal_1877, signal_1487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1287 ( .s ({signal_1878, signal_1357}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[32]), .c ({signal_1879, signal_1488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1288 ( .s ({signal_1880, signal_1356}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[33]), .c ({signal_1881, signal_1489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1289 ( .s ({signal_1878, signal_1357}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[34]), .c ({signal_1882, signal_1490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1290 ( .s ({signal_1883, signal_1361}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[35]), .c ({signal_1884, signal_1491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1291 ( .s ({signal_1885, signal_1360}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[36]), .c ({signal_1886, signal_1492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1292 ( .s ({signal_1883, signal_1361}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[37]), .c ({signal_1887, signal_1493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1293 ( .s ({signal_1888, signal_1364}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[38]), .c ({signal_1889, signal_1494}) ) ;
    buf_clk cell_1551 ( .C (clk), .D (signal_3093), .Q (signal_3094) ) ;
    buf_clk cell_1623 ( .C (clk), .D (signal_3165), .Q (signal_3166) ) ;
    buf_clk cell_1625 ( .C (clk), .D (signal_3167), .Q (signal_3168) ) ;
    buf_clk cell_1627 ( .C (clk), .D (signal_3169), .Q (signal_3170) ) ;
    buf_clk cell_1629 ( .C (clk), .D (signal_3171), .Q (signal_3172) ) ;
    buf_clk cell_1631 ( .C (clk), .D (signal_3173), .Q (signal_3174) ) ;
    buf_clk cell_1633 ( .C (clk), .D (signal_3175), .Q (signal_3176) ) ;
    buf_clk cell_1635 ( .C (clk), .D (signal_3177), .Q (signal_3178) ) ;
    buf_clk cell_1637 ( .C (clk), .D (signal_3179), .Q (signal_3180) ) ;
    buf_clk cell_1639 ( .C (clk), .D (signal_3181), .Q (signal_3182) ) ;
    buf_clk cell_1641 ( .C (clk), .D (signal_3183), .Q (signal_3184) ) ;
    buf_clk cell_1643 ( .C (clk), .D (signal_3185), .Q (signal_3186) ) ;
    buf_clk cell_1645 ( .C (clk), .D (signal_3187), .Q (signal_3188) ) ;
    buf_clk cell_1647 ( .C (clk), .D (signal_3189), .Q (signal_3190) ) ;
    buf_clk cell_1649 ( .C (clk), .D (signal_3191), .Q (signal_3192) ) ;
    buf_clk cell_1651 ( .C (clk), .D (signal_3193), .Q (signal_3194) ) ;
    buf_clk cell_1653 ( .C (clk), .D (signal_3195), .Q (signal_3196) ) ;
    buf_clk cell_1655 ( .C (clk), .D (signal_3197), .Q (signal_3198) ) ;
    buf_clk cell_1657 ( .C (clk), .D (signal_3199), .Q (signal_3200) ) ;
    buf_clk cell_1659 ( .C (clk), .D (signal_3201), .Q (signal_3202) ) ;
    buf_clk cell_1661 ( .C (clk), .D (signal_3203), .Q (signal_3204) ) ;
    buf_clk cell_1663 ( .C (clk), .D (signal_3205), .Q (signal_3206) ) ;
    buf_clk cell_1665 ( .C (clk), .D (signal_3207), .Q (signal_3208) ) ;
    buf_clk cell_1667 ( .C (clk), .D (signal_3209), .Q (signal_3210) ) ;
    buf_clk cell_1669 ( .C (clk), .D (signal_3211), .Q (signal_3212) ) ;
    buf_clk cell_1671 ( .C (clk), .D (signal_3213), .Q (signal_3214) ) ;
    buf_clk cell_1673 ( .C (clk), .D (signal_3215), .Q (signal_3216) ) ;
    buf_clk cell_1675 ( .C (clk), .D (signal_3217), .Q (signal_3218) ) ;
    buf_clk cell_1677 ( .C (clk), .D (signal_3219), .Q (signal_3220) ) ;
    buf_clk cell_1679 ( .C (clk), .D (signal_3221), .Q (signal_3222) ) ;
    buf_clk cell_1681 ( .C (clk), .D (signal_3223), .Q (signal_3224) ) ;
    buf_clk cell_1683 ( .C (clk), .D (signal_3225), .Q (signal_3226) ) ;
    buf_clk cell_1685 ( .C (clk), .D (signal_3227), .Q (signal_3228) ) ;
    buf_clk cell_1687 ( .C (clk), .D (signal_3229), .Q (signal_3230) ) ;
    buf_clk cell_1689 ( .C (clk), .D (signal_3231), .Q (signal_3232) ) ;
    buf_clk cell_1691 ( .C (clk), .D (signal_3233), .Q (signal_3234) ) ;
    buf_clk cell_1693 ( .C (clk), .D (signal_3235), .Q (signal_3236) ) ;
    buf_clk cell_1695 ( .C (clk), .D (signal_3237), .Q (signal_3238) ) ;
    buf_clk cell_1697 ( .C (clk), .D (signal_3239), .Q (signal_3240) ) ;
    buf_clk cell_1699 ( .C (clk), .D (signal_3241), .Q (signal_3242) ) ;
    buf_clk cell_1701 ( .C (clk), .D (signal_3243), .Q (signal_3244) ) ;
    buf_clk cell_1703 ( .C (clk), .D (signal_3245), .Q (signal_3246) ) ;
    buf_clk cell_1705 ( .C (clk), .D (signal_3247), .Q (signal_3248) ) ;
    buf_clk cell_1707 ( .C (clk), .D (signal_3249), .Q (signal_3250) ) ;
    buf_clk cell_1709 ( .C (clk), .D (signal_3251), .Q (signal_3252) ) ;
    buf_clk cell_1711 ( .C (clk), .D (signal_3253), .Q (signal_3254) ) ;
    buf_clk cell_1713 ( .C (clk), .D (signal_3255), .Q (signal_3256) ) ;
    buf_clk cell_1715 ( .C (clk), .D (signal_3257), .Q (signal_3258) ) ;
    buf_clk cell_1717 ( .C (clk), .D (signal_3259), .Q (signal_3260) ) ;
    buf_clk cell_1719 ( .C (clk), .D (signal_3261), .Q (signal_3262) ) ;
    buf_clk cell_1721 ( .C (clk), .D (signal_3263), .Q (signal_3264) ) ;
    buf_clk cell_1723 ( .C (clk), .D (signal_3265), .Q (signal_3266) ) ;
    buf_clk cell_1725 ( .C (clk), .D (signal_3267), .Q (signal_3268) ) ;
    buf_clk cell_1727 ( .C (clk), .D (signal_3269), .Q (signal_3270) ) ;
    buf_clk cell_1729 ( .C (clk), .D (signal_3271), .Q (signal_3272) ) ;
    buf_clk cell_1731 ( .C (clk), .D (signal_3273), .Q (signal_3274) ) ;
    buf_clk cell_1733 ( .C (clk), .D (signal_3275), .Q (signal_3276) ) ;
    buf_clk cell_1735 ( .C (clk), .D (signal_3277), .Q (signal_3278) ) ;
    buf_clk cell_1737 ( .C (clk), .D (signal_3279), .Q (signal_3280) ) ;
    buf_clk cell_1739 ( .C (clk), .D (signal_3281), .Q (signal_3282) ) ;
    buf_clk cell_1741 ( .C (clk), .D (signal_3283), .Q (signal_3284) ) ;
    buf_clk cell_1743 ( .C (clk), .D (signal_3285), .Q (signal_3286) ) ;
    buf_clk cell_1745 ( .C (clk), .D (signal_3287), .Q (signal_3288) ) ;
    buf_clk cell_1747 ( .C (clk), .D (signal_3289), .Q (signal_3290) ) ;
    buf_clk cell_1749 ( .C (clk), .D (signal_3291), .Q (signal_3292) ) ;
    buf_clk cell_1751 ( .C (clk), .D (signal_3293), .Q (signal_3294) ) ;
    buf_clk cell_1757 ( .C (clk), .D (signal_3299), .Q (signal_3300) ) ;
    buf_clk cell_1763 ( .C (clk), .D (signal_3305), .Q (signal_3306) ) ;
    buf_clk cell_1769 ( .C (clk), .D (signal_3311), .Q (signal_3312) ) ;
    buf_clk cell_1775 ( .C (clk), .D (signal_3317), .Q (signal_3318) ) ;
    buf_clk cell_1781 ( .C (clk), .D (signal_3323), .Q (signal_3324) ) ;
    buf_clk cell_1787 ( .C (clk), .D (signal_3329), .Q (signal_3330) ) ;
    buf_clk cell_1793 ( .C (clk), .D (signal_3335), .Q (signal_3336) ) ;
    buf_clk cell_1799 ( .C (clk), .D (signal_3341), .Q (signal_3342) ) ;
    buf_clk cell_1805 ( .C (clk), .D (signal_3347), .Q (signal_3348) ) ;
    buf_clk cell_1811 ( .C (clk), .D (signal_3353), .Q (signal_3354) ) ;
    buf_clk cell_1817 ( .C (clk), .D (signal_3359), .Q (signal_3360) ) ;
    buf_clk cell_1823 ( .C (clk), .D (signal_3365), .Q (signal_3366) ) ;
    buf_clk cell_1829 ( .C (clk), .D (signal_3371), .Q (signal_3372) ) ;
    buf_clk cell_1835 ( .C (clk), .D (signal_3377), .Q (signal_3378) ) ;
    buf_clk cell_1841 ( .C (clk), .D (signal_3383), .Q (signal_3384) ) ;
    buf_clk cell_1847 ( .C (clk), .D (signal_3389), .Q (signal_3390) ) ;
    buf_clk cell_1853 ( .C (clk), .D (signal_3395), .Q (signal_3396) ) ;
    buf_clk cell_1859 ( .C (clk), .D (signal_3401), .Q (signal_3402) ) ;
    buf_clk cell_1865 ( .C (clk), .D (signal_3407), .Q (signal_3408) ) ;
    buf_clk cell_1871 ( .C (clk), .D (signal_3413), .Q (signal_3414) ) ;
    buf_clk cell_1877 ( .C (clk), .D (signal_3419), .Q (signal_3420) ) ;
    buf_clk cell_1883 ( .C (clk), .D (signal_3425), .Q (signal_3426) ) ;
    buf_clk cell_1889 ( .C (clk), .D (signal_3431), .Q (signal_3432) ) ;
    buf_clk cell_1895 ( .C (clk), .D (signal_3437), .Q (signal_3438) ) ;
    buf_clk cell_1901 ( .C (clk), .D (signal_3443), .Q (signal_3444) ) ;
    buf_clk cell_1907 ( .C (clk), .D (signal_3449), .Q (signal_3450) ) ;
    buf_clk cell_1913 ( .C (clk), .D (signal_3455), .Q (signal_3456) ) ;
    buf_clk cell_1919 ( .C (clk), .D (signal_3461), .Q (signal_3462) ) ;
    buf_clk cell_1925 ( .C (clk), .D (signal_3467), .Q (signal_3468) ) ;
    buf_clk cell_1931 ( .C (clk), .D (signal_3473), .Q (signal_3474) ) ;
    buf_clk cell_1937 ( .C (clk), .D (signal_3479), .Q (signal_3480) ) ;
    buf_clk cell_1943 ( .C (clk), .D (signal_3485), .Q (signal_3486) ) ;
    buf_clk cell_1949 ( .C (clk), .D (signal_3491), .Q (signal_3492) ) ;
    buf_clk cell_1955 ( .C (clk), .D (signal_3497), .Q (signal_3498) ) ;
    buf_clk cell_1961 ( .C (clk), .D (signal_3503), .Q (signal_3504) ) ;
    buf_clk cell_1967 ( .C (clk), .D (signal_3509), .Q (signal_3510) ) ;
    buf_clk cell_1973 ( .C (clk), .D (signal_3515), .Q (signal_3516) ) ;
    buf_clk cell_1979 ( .C (clk), .D (signal_3521), .Q (signal_3522) ) ;
    buf_clk cell_1985 ( .C (clk), .D (signal_3527), .Q (signal_3528) ) ;
    buf_clk cell_1991 ( .C (clk), .D (signal_3533), .Q (signal_3534) ) ;
    buf_clk cell_1997 ( .C (clk), .D (signal_3539), .Q (signal_3540) ) ;
    buf_clk cell_2003 ( .C (clk), .D (signal_3545), .Q (signal_3546) ) ;
    buf_clk cell_2009 ( .C (clk), .D (signal_3551), .Q (signal_3552) ) ;
    buf_clk cell_2015 ( .C (clk), .D (signal_3557), .Q (signal_3558) ) ;
    buf_clk cell_2021 ( .C (clk), .D (signal_3563), .Q (signal_3564) ) ;
    buf_clk cell_2027 ( .C (clk), .D (signal_3569), .Q (signal_3570) ) ;
    buf_clk cell_2033 ( .C (clk), .D (signal_3575), .Q (signal_3576) ) ;
    buf_clk cell_2039 ( .C (clk), .D (signal_3581), .Q (signal_3582) ) ;
    buf_clk cell_2045 ( .C (clk), .D (signal_3587), .Q (signal_3588) ) ;
    buf_clk cell_2051 ( .C (clk), .D (signal_3593), .Q (signal_3594) ) ;
    buf_clk cell_2057 ( .C (clk), .D (signal_3599), .Q (signal_3600) ) ;
    buf_clk cell_2063 ( .C (clk), .D (signal_3605), .Q (signal_3606) ) ;
    buf_clk cell_2069 ( .C (clk), .D (signal_3611), .Q (signal_3612) ) ;
    buf_clk cell_2075 ( .C (clk), .D (signal_3617), .Q (signal_3618) ) ;
    buf_clk cell_2081 ( .C (clk), .D (signal_3623), .Q (signal_3624) ) ;
    buf_clk cell_2087 ( .C (clk), .D (signal_3629), .Q (signal_3630) ) ;
    buf_clk cell_2093 ( .C (clk), .D (signal_3635), .Q (signal_3636) ) ;
    buf_clk cell_2099 ( .C (clk), .D (signal_3641), .Q (signal_3642) ) ;
    buf_clk cell_2105 ( .C (clk), .D (signal_3647), .Q (signal_3648) ) ;
    buf_clk cell_2111 ( .C (clk), .D (signal_3653), .Q (signal_3654) ) ;
    buf_clk cell_2117 ( .C (clk), .D (signal_3659), .Q (signal_3660) ) ;
    buf_clk cell_2123 ( .C (clk), .D (signal_3665), .Q (signal_3666) ) ;
    buf_clk cell_2129 ( .C (clk), .D (signal_3671), .Q (signal_3672) ) ;
    buf_clk cell_2135 ( .C (clk), .D (signal_3677), .Q (signal_3678) ) ;
    buf_clk cell_2141 ( .C (clk), .D (signal_3683), .Q (signal_3684) ) ;
    buf_clk cell_2147 ( .C (clk), .D (signal_3689), .Q (signal_3690) ) ;
    buf_clk cell_2153 ( .C (clk), .D (signal_3695), .Q (signal_3696) ) ;
    buf_clk cell_2159 ( .C (clk), .D (signal_3701), .Q (signal_3702) ) ;
    buf_clk cell_2165 ( .C (clk), .D (signal_3707), .Q (signal_3708) ) ;
    buf_clk cell_2171 ( .C (clk), .D (signal_3713), .Q (signal_3714) ) ;
    buf_clk cell_2177 ( .C (clk), .D (signal_3719), .Q (signal_3720) ) ;
    buf_clk cell_2183 ( .C (clk), .D (signal_3725), .Q (signal_3726) ) ;
    buf_clk cell_2189 ( .C (clk), .D (signal_3731), .Q (signal_3732) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_3737), .Q (signal_3738) ) ;
    buf_clk cell_2201 ( .C (clk), .D (signal_3743), .Q (signal_3744) ) ;
    buf_clk cell_2207 ( .C (clk), .D (signal_3749), .Q (signal_3750) ) ;
    buf_clk cell_2213 ( .C (clk), .D (signal_3755), .Q (signal_3756) ) ;
    buf_clk cell_2219 ( .C (clk), .D (signal_3761), .Q (signal_3762) ) ;
    buf_clk cell_2225 ( .C (clk), .D (signal_3767), .Q (signal_3768) ) ;
    buf_clk cell_2231 ( .C (clk), .D (signal_3773), .Q (signal_3774) ) ;
    buf_clk cell_2237 ( .C (clk), .D (signal_3779), .Q (signal_3780) ) ;
    buf_clk cell_2243 ( .C (clk), .D (signal_3785), .Q (signal_3786) ) ;
    buf_clk cell_2249 ( .C (clk), .D (signal_3791), .Q (signal_3792) ) ;
    buf_clk cell_2255 ( .C (clk), .D (signal_3797), .Q (signal_3798) ) ;
    buf_clk cell_2261 ( .C (clk), .D (signal_3803), .Q (signal_3804) ) ;
    buf_clk cell_2267 ( .C (clk), .D (signal_3809), .Q (signal_3810) ) ;
    buf_clk cell_2273 ( .C (clk), .D (signal_3815), .Q (signal_3816) ) ;
    buf_clk cell_2279 ( .C (clk), .D (signal_3821), .Q (signal_3822) ) ;
    buf_clk cell_2285 ( .C (clk), .D (signal_3827), .Q (signal_3828) ) ;
    buf_clk cell_2291 ( .C (clk), .D (signal_3833), .Q (signal_3834) ) ;
    buf_clk cell_2297 ( .C (clk), .D (signal_3839), .Q (signal_3840) ) ;
    buf_clk cell_2303 ( .C (clk), .D (signal_3845), .Q (signal_3846) ) ;
    buf_clk cell_2309 ( .C (clk), .D (signal_3851), .Q (signal_3852) ) ;
    buf_clk cell_2315 ( .C (clk), .D (signal_3857), .Q (signal_3858) ) ;
    buf_clk cell_2321 ( .C (clk), .D (signal_3863), .Q (signal_3864) ) ;
    buf_clk cell_2327 ( .C (clk), .D (signal_3869), .Q (signal_3870) ) ;
    buf_clk cell_2333 ( .C (clk), .D (signal_3875), .Q (signal_3876) ) ;
    buf_clk cell_2339 ( .C (clk), .D (signal_3881), .Q (signal_3882) ) ;
    buf_clk cell_2345 ( .C (clk), .D (signal_3887), .Q (signal_3888) ) ;
    buf_clk cell_2351 ( .C (clk), .D (signal_3893), .Q (signal_3894) ) ;
    buf_clk cell_2357 ( .C (clk), .D (signal_3899), .Q (signal_3900) ) ;
    buf_clk cell_2363 ( .C (clk), .D (signal_3905), .Q (signal_3906) ) ;
    buf_clk cell_2369 ( .C (clk), .D (signal_3911), .Q (signal_3912) ) ;
    buf_clk cell_2375 ( .C (clk), .D (signal_3917), .Q (signal_3918) ) ;
    buf_clk cell_2381 ( .C (clk), .D (signal_3923), .Q (signal_3924) ) ;
    buf_clk cell_2387 ( .C (clk), .D (signal_3929), .Q (signal_3930) ) ;
    buf_clk cell_2393 ( .C (clk), .D (signal_3935), .Q (signal_3936) ) ;
    buf_clk cell_2399 ( .C (clk), .D (signal_3941), .Q (signal_3942) ) ;
    buf_clk cell_2405 ( .C (clk), .D (signal_3947), .Q (signal_3948) ) ;
    buf_clk cell_2411 ( .C (clk), .D (signal_3953), .Q (signal_3954) ) ;
    buf_clk cell_2417 ( .C (clk), .D (signal_3959), .Q (signal_3960) ) ;
    buf_clk cell_2423 ( .C (clk), .D (signal_3965), .Q (signal_3966) ) ;
    buf_clk cell_2429 ( .C (clk), .D (signal_3971), .Q (signal_3972) ) ;
    buf_clk cell_2435 ( .C (clk), .D (signal_3977), .Q (signal_3978) ) ;
    buf_clk cell_2441 ( .C (clk), .D (signal_3983), .Q (signal_3984) ) ;
    buf_clk cell_2447 ( .C (clk), .D (signal_3989), .Q (signal_3990) ) ;
    buf_clk cell_2453 ( .C (clk), .D (signal_3995), .Q (signal_3996) ) ;
    buf_clk cell_2459 ( .C (clk), .D (signal_4001), .Q (signal_4002) ) ;
    buf_clk cell_2465 ( .C (clk), .D (signal_4007), .Q (signal_4008) ) ;
    buf_clk cell_2471 ( .C (clk), .D (signal_4013), .Q (signal_4014) ) ;
    buf_clk cell_2477 ( .C (clk), .D (signal_4019), .Q (signal_4020) ) ;
    buf_clk cell_2483 ( .C (clk), .D (signal_4025), .Q (signal_4026) ) ;
    buf_clk cell_2489 ( .C (clk), .D (signal_4031), .Q (signal_4032) ) ;
    buf_clk cell_2495 ( .C (clk), .D (signal_4037), .Q (signal_4038) ) ;
    buf_clk cell_2501 ( .C (clk), .D (signal_4043), .Q (signal_4044) ) ;
    buf_clk cell_2507 ( .C (clk), .D (signal_4049), .Q (signal_4050) ) ;
    buf_clk cell_2513 ( .C (clk), .D (signal_4055), .Q (signal_4056) ) ;
    buf_clk cell_2519 ( .C (clk), .D (signal_4061), .Q (signal_4062) ) ;
    buf_clk cell_2525 ( .C (clk), .D (signal_4067), .Q (signal_4068) ) ;
    buf_clk cell_2531 ( .C (clk), .D (signal_4073), .Q (signal_4074) ) ;
    buf_clk cell_2537 ( .C (clk), .D (signal_4079), .Q (signal_4080) ) ;
    buf_clk cell_2543 ( .C (clk), .D (signal_4085), .Q (signal_4086) ) ;
    buf_clk cell_2549 ( .C (clk), .D (signal_4091), .Q (signal_4092) ) ;
    buf_clk cell_2555 ( .C (clk), .D (signal_4097), .Q (signal_4098) ) ;
    buf_clk cell_2561 ( .C (clk), .D (signal_4103), .Q (signal_4104) ) ;
    buf_clk cell_2567 ( .C (clk), .D (signal_4109), .Q (signal_4110) ) ;
    buf_clk cell_2573 ( .C (clk), .D (signal_4115), .Q (signal_4116) ) ;
    buf_clk cell_2579 ( .C (clk), .D (signal_4121), .Q (signal_4122) ) ;
    buf_clk cell_2585 ( .C (clk), .D (signal_4127), .Q (signal_4128) ) ;
    buf_clk cell_2591 ( .C (clk), .D (signal_4133), .Q (signal_4134) ) ;
    buf_clk cell_2597 ( .C (clk), .D (signal_4139), .Q (signal_4140) ) ;
    buf_clk cell_2603 ( .C (clk), .D (signal_4145), .Q (signal_4146) ) ;
    buf_clk cell_2609 ( .C (clk), .D (signal_4151), .Q (signal_4152) ) ;
    buf_clk cell_2615 ( .C (clk), .D (signal_4157), .Q (signal_4158) ) ;
    buf_clk cell_2621 ( .C (clk), .D (signal_4163), .Q (signal_4164) ) ;
    buf_clk cell_2627 ( .C (clk), .D (signal_4169), .Q (signal_4170) ) ;
    buf_clk cell_2633 ( .C (clk), .D (signal_4175), .Q (signal_4176) ) ;
    buf_clk cell_2639 ( .C (clk), .D (signal_4181), .Q (signal_4182) ) ;
    buf_clk cell_2645 ( .C (clk), .D (signal_4187), .Q (signal_4188) ) ;
    buf_clk cell_2651 ( .C (clk), .D (signal_4193), .Q (signal_4194) ) ;
    buf_clk cell_2657 ( .C (clk), .D (signal_4199), .Q (signal_4200) ) ;
    buf_clk cell_2663 ( .C (clk), .D (signal_4205), .Q (signal_4206) ) ;
    buf_clk cell_2669 ( .C (clk), .D (signal_4211), .Q (signal_4212) ) ;
    buf_clk cell_2675 ( .C (clk), .D (signal_4217), .Q (signal_4218) ) ;
    buf_clk cell_2681 ( .C (clk), .D (signal_4223), .Q (signal_4224) ) ;
    buf_clk cell_2687 ( .C (clk), .D (signal_4229), .Q (signal_4230) ) ;
    buf_clk cell_2693 ( .C (clk), .D (signal_4235), .Q (signal_4236) ) ;
    buf_clk cell_2699 ( .C (clk), .D (signal_4241), .Q (signal_4242) ) ;
    buf_clk cell_2705 ( .C (clk), .D (signal_4247), .Q (signal_4248) ) ;
    buf_clk cell_2711 ( .C (clk), .D (signal_4253), .Q (signal_4254) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_4259), .Q (signal_4260) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_4265), .Q (signal_4266) ) ;
    buf_clk cell_2729 ( .C (clk), .D (signal_4271), .Q (signal_4272) ) ;
    buf_clk cell_2735 ( .C (clk), .D (signal_4277), .Q (signal_4278) ) ;
    buf_clk cell_2741 ( .C (clk), .D (signal_4283), .Q (signal_4284) ) ;
    buf_clk cell_2747 ( .C (clk), .D (signal_4289), .Q (signal_4290) ) ;
    buf_clk cell_2753 ( .C (clk), .D (signal_4295), .Q (signal_4296) ) ;
    buf_clk cell_2759 ( .C (clk), .D (signal_4301), .Q (signal_4302) ) ;
    buf_clk cell_2765 ( .C (clk), .D (signal_4307), .Q (signal_4308) ) ;
    buf_clk cell_2771 ( .C (clk), .D (signal_4313), .Q (signal_4314) ) ;
    buf_clk cell_2777 ( .C (clk), .D (signal_4319), .Q (signal_4320) ) ;
    buf_clk cell_2783 ( .C (clk), .D (signal_4325), .Q (signal_4326) ) ;
    buf_clk cell_2789 ( .C (clk), .D (signal_4331), .Q (signal_4332) ) ;
    buf_clk cell_2795 ( .C (clk), .D (signal_4337), .Q (signal_4338) ) ;
    buf_clk cell_2801 ( .C (clk), .D (signal_4343), .Q (signal_4344) ) ;
    buf_clk cell_2807 ( .C (clk), .D (signal_4349), .Q (signal_4350) ) ;
    buf_clk cell_2813 ( .C (clk), .D (signal_4355), .Q (signal_4356) ) ;
    buf_clk cell_2819 ( .C (clk), .D (signal_4361), .Q (signal_4362) ) ;
    buf_clk cell_2825 ( .C (clk), .D (signal_4367), .Q (signal_4368) ) ;
    buf_clk cell_2831 ( .C (clk), .D (signal_4373), .Q (signal_4374) ) ;
    buf_clk cell_2837 ( .C (clk), .D (signal_4379), .Q (signal_4380) ) ;
    buf_clk cell_2843 ( .C (clk), .D (signal_4385), .Q (signal_4386) ) ;
    buf_clk cell_2849 ( .C (clk), .D (signal_4391), .Q (signal_4392) ) ;
    buf_clk cell_2855 ( .C (clk), .D (signal_4397), .Q (signal_4398) ) ;
    buf_clk cell_2861 ( .C (clk), .D (signal_4403), .Q (signal_4404) ) ;
    buf_clk cell_2867 ( .C (clk), .D (signal_4409), .Q (signal_4410) ) ;
    buf_clk cell_2873 ( .C (clk), .D (signal_4415), .Q (signal_4416) ) ;
    buf_clk cell_2879 ( .C (clk), .D (signal_4421), .Q (signal_4422) ) ;
    buf_clk cell_2885 ( .C (clk), .D (signal_4427), .Q (signal_4428) ) ;
    buf_clk cell_2891 ( .C (clk), .D (signal_4433), .Q (signal_4434) ) ;
    buf_clk cell_2897 ( .C (clk), .D (signal_4439), .Q (signal_4440) ) ;
    buf_clk cell_2903 ( .C (clk), .D (signal_4445), .Q (signal_4446) ) ;
    buf_clk cell_2909 ( .C (clk), .D (signal_4451), .Q (signal_4452) ) ;
    buf_clk cell_2919 ( .C (clk), .D (signal_4461), .Q (signal_4462) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_4465), .Q (signal_4466) ) ;
    buf_clk cell_2955 ( .C (clk), .D (signal_4497), .Q (signal_4498) ) ;
    buf_clk cell_2959 ( .C (clk), .D (signal_4501), .Q (signal_4502) ) ;
    buf_clk cell_2963 ( .C (clk), .D (signal_4505), .Q (signal_4506) ) ;
    buf_clk cell_2967 ( .C (clk), .D (signal_4509), .Q (signal_4510) ) ;
    buf_clk cell_2975 ( .C (clk), .D (signal_4517), .Q (signal_4518) ) ;
    buf_clk cell_2979 ( .C (clk), .D (signal_4521), .Q (signal_4522) ) ;
    buf_clk cell_2983 ( .C (clk), .D (signal_4525), .Q (signal_4526) ) ;
    buf_clk cell_2987 ( .C (clk), .D (signal_4529), .Q (signal_4530) ) ;
    buf_clk cell_2991 ( .C (clk), .D (signal_4533), .Q (signal_4534) ) ;
    buf_clk cell_2995 ( .C (clk), .D (signal_4537), .Q (signal_4538) ) ;
    buf_clk cell_3003 ( .C (clk), .D (signal_4545), .Q (signal_4546) ) ;
    buf_clk cell_3007 ( .C (clk), .D (signal_4549), .Q (signal_4550) ) ;
    buf_clk cell_3011 ( .C (clk), .D (signal_4553), .Q (signal_4554) ) ;
    buf_clk cell_3015 ( .C (clk), .D (signal_4557), .Q (signal_4558) ) ;
    buf_clk cell_3019 ( .C (clk), .D (signal_4561), .Q (signal_4562) ) ;
    buf_clk cell_3023 ( .C (clk), .D (signal_4565), .Q (signal_4566) ) ;
    buf_clk cell_3027 ( .C (clk), .D (signal_4569), .Q (signal_4570) ) ;
    buf_clk cell_3031 ( .C (clk), .D (signal_4573), .Q (signal_4574) ) ;
    buf_clk cell_3035 ( .C (clk), .D (signal_4577), .Q (signal_4578) ) ;
    buf_clk cell_3039 ( .C (clk), .D (signal_4581), .Q (signal_4582) ) ;
    buf_clk cell_3051 ( .C (clk), .D (signal_4593), .Q (signal_4594) ) ;
    buf_clk cell_3055 ( .C (clk), .D (signal_4597), .Q (signal_4598) ) ;
    buf_clk cell_3063 ( .C (clk), .D (signal_4605), .Q (signal_4606) ) ;
    buf_clk cell_3067 ( .C (clk), .D (signal_4609), .Q (signal_4610) ) ;
    buf_clk cell_3075 ( .C (clk), .D (signal_4617), .Q (signal_4618) ) ;
    buf_clk cell_3079 ( .C (clk), .D (signal_4621), .Q (signal_4622) ) ;
    buf_clk cell_3087 ( .C (clk), .D (signal_4629), .Q (signal_4630) ) ;
    buf_clk cell_3091 ( .C (clk), .D (signal_4633), .Q (signal_4634) ) ;
    buf_clk cell_3099 ( .C (clk), .D (signal_4641), .Q (signal_4642) ) ;
    buf_clk cell_3103 ( .C (clk), .D (signal_4645), .Q (signal_4646) ) ;
    buf_clk cell_3107 ( .C (clk), .D (signal_4649), .Q (signal_4650) ) ;
    buf_clk cell_3115 ( .C (clk), .D (signal_4657), .Q (signal_4658) ) ;
    buf_clk cell_3123 ( .C (clk), .D (signal_4665), .Q (signal_4666) ) ;
    buf_clk cell_3131 ( .C (clk), .D (signal_4673), .Q (signal_4674) ) ;
    buf_clk cell_3139 ( .C (clk), .D (signal_4681), .Q (signal_4682) ) ;
    buf_clk cell_3147 ( .C (clk), .D (signal_4689), .Q (signal_4690) ) ;
    buf_clk cell_3155 ( .C (clk), .D (signal_4697), .Q (signal_4698) ) ;
    buf_clk cell_3163 ( .C (clk), .D (signal_4705), .Q (signal_4706) ) ;
    buf_clk cell_3171 ( .C (clk), .D (signal_4713), .Q (signal_4714) ) ;
    buf_clk cell_3179 ( .C (clk), .D (signal_4721), .Q (signal_4722) ) ;
    buf_clk cell_3187 ( .C (clk), .D (signal_4729), .Q (signal_4730) ) ;
    buf_clk cell_3195 ( .C (clk), .D (signal_4737), .Q (signal_4738) ) ;
    buf_clk cell_3203 ( .C (clk), .D (signal_4745), .Q (signal_4746) ) ;
    buf_clk cell_3211 ( .C (clk), .D (signal_4753), .Q (signal_4754) ) ;
    buf_clk cell_3219 ( .C (clk), .D (signal_4761), .Q (signal_4762) ) ;
    buf_clk cell_3227 ( .C (clk), .D (signal_4769), .Q (signal_4770) ) ;
    buf_clk cell_3235 ( .C (clk), .D (signal_4777), .Q (signal_4778) ) ;
    buf_clk cell_3243 ( .C (clk), .D (signal_4785), .Q (signal_4786) ) ;
    buf_clk cell_3251 ( .C (clk), .D (signal_4793), .Q (signal_4794) ) ;
    buf_clk cell_3259 ( .C (clk), .D (signal_4801), .Q (signal_4802) ) ;
    buf_clk cell_3267 ( .C (clk), .D (signal_4809), .Q (signal_4810) ) ;
    buf_clk cell_3275 ( .C (clk), .D (signal_4817), .Q (signal_4818) ) ;
    buf_clk cell_3283 ( .C (clk), .D (signal_4825), .Q (signal_4826) ) ;
    buf_clk cell_3291 ( .C (clk), .D (signal_4833), .Q (signal_4834) ) ;
    buf_clk cell_3299 ( .C (clk), .D (signal_4841), .Q (signal_4842) ) ;
    buf_clk cell_3307 ( .C (clk), .D (signal_4849), .Q (signal_4850) ) ;
    buf_clk cell_3315 ( .C (clk), .D (signal_4857), .Q (signal_4858) ) ;
    buf_clk cell_3323 ( .C (clk), .D (signal_4865), .Q (signal_4866) ) ;
    buf_clk cell_3331 ( .C (clk), .D (signal_4873), .Q (signal_4874) ) ;
    buf_clk cell_3339 ( .C (clk), .D (signal_4881), .Q (signal_4882) ) ;
    buf_clk cell_3347 ( .C (clk), .D (signal_4889), .Q (signal_4890) ) ;
    buf_clk cell_3355 ( .C (clk), .D (signal_4897), .Q (signal_4898) ) ;
    buf_clk cell_3363 ( .C (clk), .D (signal_4905), .Q (signal_4906) ) ;
    buf_clk cell_3371 ( .C (clk), .D (signal_4913), .Q (signal_4914) ) ;
    buf_clk cell_3379 ( .C (clk), .D (signal_4921), .Q (signal_4922) ) ;
    buf_clk cell_3387 ( .C (clk), .D (signal_4929), .Q (signal_4930) ) ;
    buf_clk cell_3395 ( .C (clk), .D (signal_4937), .Q (signal_4938) ) ;
    buf_clk cell_3403 ( .C (clk), .D (signal_4945), .Q (signal_4946) ) ;
    buf_clk cell_3411 ( .C (clk), .D (signal_4953), .Q (signal_4954) ) ;
    buf_clk cell_3419 ( .C (clk), .D (signal_4961), .Q (signal_4962) ) ;
    buf_clk cell_3427 ( .C (clk), .D (signal_4969), .Q (signal_4970) ) ;
    buf_clk cell_3435 ( .C (clk), .D (signal_4977), .Q (signal_4978) ) ;
    buf_clk cell_3443 ( .C (clk), .D (signal_4985), .Q (signal_4986) ) ;
    buf_clk cell_3451 ( .C (clk), .D (signal_4993), .Q (signal_4994) ) ;
    buf_clk cell_3459 ( .C (clk), .D (signal_5001), .Q (signal_5002) ) ;
    buf_clk cell_3467 ( .C (clk), .D (signal_5009), .Q (signal_5010) ) ;
    buf_clk cell_3475 ( .C (clk), .D (signal_5017), .Q (signal_5018) ) ;
    buf_clk cell_3483 ( .C (clk), .D (signal_5025), .Q (signal_5026) ) ;
    buf_clk cell_3491 ( .C (clk), .D (signal_5033), .Q (signal_5034) ) ;
    buf_clk cell_3499 ( .C (clk), .D (signal_5041), .Q (signal_5042) ) ;
    buf_clk cell_3507 ( .C (clk), .D (signal_5049), .Q (signal_5050) ) ;
    buf_clk cell_3515 ( .C (clk), .D (signal_5057), .Q (signal_5058) ) ;
    buf_clk cell_3523 ( .C (clk), .D (signal_5065), .Q (signal_5066) ) ;
    buf_clk cell_3531 ( .C (clk), .D (signal_5073), .Q (signal_5074) ) ;
    buf_clk cell_3539 ( .C (clk), .D (signal_5081), .Q (signal_5082) ) ;
    buf_clk cell_3547 ( .C (clk), .D (signal_5089), .Q (signal_5090) ) ;
    buf_clk cell_3555 ( .C (clk), .D (signal_5097), .Q (signal_5098) ) ;
    buf_clk cell_3563 ( .C (clk), .D (signal_5105), .Q (signal_5106) ) ;
    buf_clk cell_3571 ( .C (clk), .D (signal_5113), .Q (signal_5114) ) ;
    buf_clk cell_3579 ( .C (clk), .D (signal_5121), .Q (signal_5122) ) ;
    buf_clk cell_3587 ( .C (clk), .D (signal_5129), .Q (signal_5130) ) ;
    buf_clk cell_3595 ( .C (clk), .D (signal_5137), .Q (signal_5138) ) ;
    buf_clk cell_3603 ( .C (clk), .D (signal_5145), .Q (signal_5146) ) ;
    buf_clk cell_3611 ( .C (clk), .D (signal_5153), .Q (signal_5154) ) ;
    buf_clk cell_3619 ( .C (clk), .D (signal_5161), .Q (signal_5162) ) ;
    buf_clk cell_3627 ( .C (clk), .D (signal_5169), .Q (signal_5170) ) ;
    buf_clk cell_3635 ( .C (clk), .D (signal_5177), .Q (signal_5178) ) ;
    buf_clk cell_3643 ( .C (clk), .D (signal_5185), .Q (signal_5186) ) ;
    buf_clk cell_3651 ( .C (clk), .D (signal_5193), .Q (signal_5194) ) ;
    buf_clk cell_3659 ( .C (clk), .D (signal_5201), .Q (signal_5202) ) ;
    buf_clk cell_3667 ( .C (clk), .D (signal_5209), .Q (signal_5210) ) ;
    buf_clk cell_3675 ( .C (clk), .D (signal_5217), .Q (signal_5218) ) ;
    buf_clk cell_3683 ( .C (clk), .D (signal_5225), .Q (signal_5226) ) ;
    buf_clk cell_3691 ( .C (clk), .D (signal_5233), .Q (signal_5234) ) ;
    buf_clk cell_3699 ( .C (clk), .D (signal_5241), .Q (signal_5242) ) ;
    buf_clk cell_3707 ( .C (clk), .D (signal_5249), .Q (signal_5250) ) ;
    buf_clk cell_3715 ( .C (clk), .D (signal_5257), .Q (signal_5258) ) ;
    buf_clk cell_3723 ( .C (clk), .D (signal_5265), .Q (signal_5266) ) ;
    buf_clk cell_3731 ( .C (clk), .D (signal_5273), .Q (signal_5274) ) ;
    buf_clk cell_3739 ( .C (clk), .D (signal_5281), .Q (signal_5282) ) ;
    buf_clk cell_3747 ( .C (clk), .D (signal_5289), .Q (signal_5290) ) ;
    buf_clk cell_3755 ( .C (clk), .D (signal_5297), .Q (signal_5298) ) ;
    buf_clk cell_3763 ( .C (clk), .D (signal_5305), .Q (signal_5306) ) ;
    buf_clk cell_3771 ( .C (clk), .D (signal_5313), .Q (signal_5314) ) ;
    buf_clk cell_3779 ( .C (clk), .D (signal_5321), .Q (signal_5322) ) ;
    buf_clk cell_3787 ( .C (clk), .D (signal_5329), .Q (signal_5330) ) ;
    buf_clk cell_3795 ( .C (clk), .D (signal_5337), .Q (signal_5338) ) ;
    buf_clk cell_3803 ( .C (clk), .D (signal_5345), .Q (signal_5346) ) ;
    buf_clk cell_3811 ( .C (clk), .D (signal_5353), .Q (signal_5354) ) ;
    buf_clk cell_3819 ( .C (clk), .D (signal_5361), .Q (signal_5362) ) ;
    buf_clk cell_3827 ( .C (clk), .D (signal_5369), .Q (signal_5370) ) ;
    buf_clk cell_3835 ( .C (clk), .D (signal_5377), .Q (signal_5378) ) ;
    buf_clk cell_3843 ( .C (clk), .D (signal_5385), .Q (signal_5386) ) ;
    buf_clk cell_3851 ( .C (clk), .D (signal_5393), .Q (signal_5394) ) ;
    buf_clk cell_3859 ( .C (clk), .D (signal_5401), .Q (signal_5402) ) ;
    buf_clk cell_3867 ( .C (clk), .D (signal_5409), .Q (signal_5410) ) ;
    buf_clk cell_3875 ( .C (clk), .D (signal_5417), .Q (signal_5418) ) ;
    buf_clk cell_3883 ( .C (clk), .D (signal_5425), .Q (signal_5426) ) ;
    buf_clk cell_3891 ( .C (clk), .D (signal_5433), .Q (signal_5434) ) ;
    buf_clk cell_3899 ( .C (clk), .D (signal_5441), .Q (signal_5442) ) ;
    buf_clk cell_3907 ( .C (clk), .D (signal_5449), .Q (signal_5450) ) ;
    buf_clk cell_3915 ( .C (clk), .D (signal_5457), .Q (signal_5458) ) ;
    buf_clk cell_3923 ( .C (clk), .D (signal_5465), .Q (signal_5466) ) ;
    buf_clk cell_3931 ( .C (clk), .D (signal_5473), .Q (signal_5474) ) ;
    buf_clk cell_3939 ( .C (clk), .D (signal_5481), .Q (signal_5482) ) ;
    buf_clk cell_3947 ( .C (clk), .D (signal_5489), .Q (signal_5490) ) ;
    buf_clk cell_3955 ( .C (clk), .D (signal_5497), .Q (signal_5498) ) ;
    buf_clk cell_3963 ( .C (clk), .D (signal_5505), .Q (signal_5506) ) ;
    buf_clk cell_3971 ( .C (clk), .D (signal_5513), .Q (signal_5514) ) ;
    buf_clk cell_3979 ( .C (clk), .D (signal_5521), .Q (signal_5522) ) ;
    buf_clk cell_3987 ( .C (clk), .D (signal_5529), .Q (signal_5530) ) ;
    buf_clk cell_3995 ( .C (clk), .D (signal_5537), .Q (signal_5538) ) ;
    buf_clk cell_4003 ( .C (clk), .D (signal_5545), .Q (signal_5546) ) ;
    buf_clk cell_4011 ( .C (clk), .D (signal_5553), .Q (signal_5554) ) ;
    buf_clk cell_4019 ( .C (clk), .D (signal_5561), .Q (signal_5562) ) ;
    buf_clk cell_4027 ( .C (clk), .D (signal_5569), .Q (signal_5570) ) ;
    buf_clk cell_4035 ( .C (clk), .D (signal_5577), .Q (signal_5578) ) ;
    buf_clk cell_4043 ( .C (clk), .D (signal_5585), .Q (signal_5586) ) ;
    buf_clk cell_4051 ( .C (clk), .D (signal_5593), .Q (signal_5594) ) ;
    buf_clk cell_4059 ( .C (clk), .D (signal_5601), .Q (signal_5602) ) ;
    buf_clk cell_4067 ( .C (clk), .D (signal_5609), .Q (signal_5610) ) ;
    buf_clk cell_4075 ( .C (clk), .D (signal_5617), .Q (signal_5618) ) ;
    buf_clk cell_4083 ( .C (clk), .D (signal_5625), .Q (signal_5626) ) ;
    buf_clk cell_4091 ( .C (clk), .D (signal_5633), .Q (signal_5634) ) ;
    buf_clk cell_4099 ( .C (clk), .D (signal_5641), .Q (signal_5642) ) ;
    buf_clk cell_4107 ( .C (clk), .D (signal_5649), .Q (signal_5650) ) ;
    buf_clk cell_4115 ( .C (clk), .D (signal_5657), .Q (signal_5658) ) ;
    buf_clk cell_4123 ( .C (clk), .D (signal_5665), .Q (signal_5666) ) ;
    buf_clk cell_4133 ( .C (clk), .D (signal_5675), .Q (signal_5676) ) ;
    buf_clk cell_4141 ( .C (clk), .D (signal_5683), .Q (signal_5684) ) ;
    buf_clk cell_4149 ( .C (clk), .D (signal_5691), .Q (signal_5692) ) ;
    buf_clk cell_4157 ( .C (clk), .D (signal_5699), .Q (signal_5700) ) ;
    buf_clk cell_4165 ( .C (clk), .D (signal_5707), .Q (signal_5708) ) ;
    buf_clk cell_4173 ( .C (clk), .D (signal_5715), .Q (signal_5716) ) ;
    buf_clk cell_4181 ( .C (clk), .D (signal_5723), .Q (signal_5724) ) ;
    buf_clk cell_4189 ( .C (clk), .D (signal_5731), .Q (signal_5732) ) ;
    buf_clk cell_4197 ( .C (clk), .D (signal_5739), .Q (signal_5740) ) ;
    buf_clk cell_4205 ( .C (clk), .D (signal_5747), .Q (signal_5748) ) ;
    buf_clk cell_4213 ( .C (clk), .D (signal_5755), .Q (signal_5756) ) ;
    buf_clk cell_4221 ( .C (clk), .D (signal_5763), .Q (signal_5764) ) ;
    buf_clk cell_4229 ( .C (clk), .D (signal_5771), .Q (signal_5772) ) ;
    buf_clk cell_4237 ( .C (clk), .D (signal_5779), .Q (signal_5780) ) ;
    buf_clk cell_4245 ( .C (clk), .D (signal_5787), .Q (signal_5788) ) ;
    buf_clk cell_4253 ( .C (clk), .D (signal_5795), .Q (signal_5796) ) ;
    buf_clk cell_4261 ( .C (clk), .D (signal_5803), .Q (signal_5804) ) ;
    buf_clk cell_4269 ( .C (clk), .D (signal_5811), .Q (signal_5812) ) ;
    buf_clk cell_4277 ( .C (clk), .D (signal_5819), .Q (signal_5820) ) ;
    buf_clk cell_4285 ( .C (clk), .D (signal_5827), .Q (signal_5828) ) ;
    buf_clk cell_4293 ( .C (clk), .D (signal_5835), .Q (signal_5836) ) ;
    buf_clk cell_4301 ( .C (clk), .D (signal_5843), .Q (signal_5844) ) ;
    buf_clk cell_4309 ( .C (clk), .D (signal_5851), .Q (signal_5852) ) ;
    buf_clk cell_4317 ( .C (clk), .D (signal_5859), .Q (signal_5860) ) ;
    buf_clk cell_4325 ( .C (clk), .D (signal_5867), .Q (signal_5868) ) ;
    buf_clk cell_4333 ( .C (clk), .D (signal_5875), .Q (signal_5876) ) ;
    buf_clk cell_4341 ( .C (clk), .D (signal_5883), .Q (signal_5884) ) ;
    buf_clk cell_4349 ( .C (clk), .D (signal_5891), .Q (signal_5892) ) ;
    buf_clk cell_4357 ( .C (clk), .D (signal_5899), .Q (signal_5900) ) ;
    buf_clk cell_4365 ( .C (clk), .D (signal_5907), .Q (signal_5908) ) ;
    buf_clk cell_4373 ( .C (clk), .D (signal_5915), .Q (signal_5916) ) ;
    buf_clk cell_4381 ( .C (clk), .D (signal_5923), .Q (signal_5924) ) ;
    buf_clk cell_4389 ( .C (clk), .D (signal_5931), .Q (signal_5932) ) ;
    buf_clk cell_4397 ( .C (clk), .D (signal_5939), .Q (signal_5940) ) ;
    buf_clk cell_4405 ( .C (clk), .D (signal_5947), .Q (signal_5948) ) ;
    buf_clk cell_4413 ( .C (clk), .D (signal_5955), .Q (signal_5956) ) ;
    buf_clk cell_4421 ( .C (clk), .D (signal_5963), .Q (signal_5964) ) ;
    buf_clk cell_4429 ( .C (clk), .D (signal_5971), .Q (signal_5972) ) ;
    buf_clk cell_4437 ( .C (clk), .D (signal_5979), .Q (signal_5980) ) ;
    buf_clk cell_4445 ( .C (clk), .D (signal_5987), .Q (signal_5988) ) ;
    buf_clk cell_4453 ( .C (clk), .D (signal_5995), .Q (signal_5996) ) ;
    buf_clk cell_4461 ( .C (clk), .D (signal_6003), .Q (signal_6004) ) ;
    buf_clk cell_4469 ( .C (clk), .D (signal_6011), .Q (signal_6012) ) ;
    buf_clk cell_4477 ( .C (clk), .D (signal_6019), .Q (signal_6020) ) ;
    buf_clk cell_4485 ( .C (clk), .D (signal_6027), .Q (signal_6028) ) ;
    buf_clk cell_4493 ( .C (clk), .D (signal_6035), .Q (signal_6036) ) ;
    buf_clk cell_4501 ( .C (clk), .D (signal_6043), .Q (signal_6044) ) ;
    buf_clk cell_4509 ( .C (clk), .D (signal_6051), .Q (signal_6052) ) ;
    buf_clk cell_4517 ( .C (clk), .D (signal_6059), .Q (signal_6060) ) ;
    buf_clk cell_4525 ( .C (clk), .D (signal_6067), .Q (signal_6068) ) ;
    buf_clk cell_4533 ( .C (clk), .D (signal_6075), .Q (signal_6076) ) ;
    buf_clk cell_4541 ( .C (clk), .D (signal_6083), .Q (signal_6084) ) ;
    buf_clk cell_4549 ( .C (clk), .D (signal_6091), .Q (signal_6092) ) ;
    buf_clk cell_4557 ( .C (clk), .D (signal_6099), .Q (signal_6100) ) ;
    buf_clk cell_4565 ( .C (clk), .D (signal_6107), .Q (signal_6108) ) ;
    buf_clk cell_4573 ( .C (clk), .D (signal_6115), .Q (signal_6116) ) ;
    buf_clk cell_4581 ( .C (clk), .D (signal_6123), .Q (signal_6124) ) ;
    buf_clk cell_4589 ( .C (clk), .D (signal_6131), .Q (signal_6132) ) ;
    buf_clk cell_4597 ( .C (clk), .D (signal_6139), .Q (signal_6140) ) ;
    buf_clk cell_4605 ( .C (clk), .D (signal_6147), .Q (signal_6148) ) ;
    buf_clk cell_4613 ( .C (clk), .D (signal_6155), .Q (signal_6156) ) ;
    buf_clk cell_4621 ( .C (clk), .D (signal_6163), .Q (signal_6164) ) ;
    buf_clk cell_4629 ( .C (clk), .D (signal_6171), .Q (signal_6172) ) ;
    buf_clk cell_4637 ( .C (clk), .D (signal_6179), .Q (signal_6180) ) ;
    buf_clk cell_4839 ( .C (clk), .D (signal_6381), .Q (signal_6382) ) ;
    buf_clk cell_4847 ( .C (clk), .D (signal_6389), .Q (signal_6390) ) ;
    buf_clk cell_4855 ( .C (clk), .D (signal_6397), .Q (signal_6398) ) ;
    buf_clk cell_4863 ( .C (clk), .D (signal_6405), .Q (signal_6406) ) ;

    /* cells in depth 3 */
    buf_clk cell_1552 ( .C (clk), .D (signal_3094), .Q (signal_3095) ) ;
    buf_clk cell_1752 ( .C (clk), .D (signal_3294), .Q (signal_3295) ) ;
    buf_clk cell_1758 ( .C (clk), .D (signal_3300), .Q (signal_3301) ) ;
    buf_clk cell_1764 ( .C (clk), .D (signal_3306), .Q (signal_3307) ) ;
    buf_clk cell_1770 ( .C (clk), .D (signal_3312), .Q (signal_3313) ) ;
    buf_clk cell_1776 ( .C (clk), .D (signal_3318), .Q (signal_3319) ) ;
    buf_clk cell_1782 ( .C (clk), .D (signal_3324), .Q (signal_3325) ) ;
    buf_clk cell_1788 ( .C (clk), .D (signal_3330), .Q (signal_3331) ) ;
    buf_clk cell_1794 ( .C (clk), .D (signal_3336), .Q (signal_3337) ) ;
    buf_clk cell_1800 ( .C (clk), .D (signal_3342), .Q (signal_3343) ) ;
    buf_clk cell_1806 ( .C (clk), .D (signal_3348), .Q (signal_3349) ) ;
    buf_clk cell_1812 ( .C (clk), .D (signal_3354), .Q (signal_3355) ) ;
    buf_clk cell_1818 ( .C (clk), .D (signal_3360), .Q (signal_3361) ) ;
    buf_clk cell_1824 ( .C (clk), .D (signal_3366), .Q (signal_3367) ) ;
    buf_clk cell_1830 ( .C (clk), .D (signal_3372), .Q (signal_3373) ) ;
    buf_clk cell_1836 ( .C (clk), .D (signal_3378), .Q (signal_3379) ) ;
    buf_clk cell_1842 ( .C (clk), .D (signal_3384), .Q (signal_3385) ) ;
    buf_clk cell_1848 ( .C (clk), .D (signal_3390), .Q (signal_3391) ) ;
    buf_clk cell_1854 ( .C (clk), .D (signal_3396), .Q (signal_3397) ) ;
    buf_clk cell_1860 ( .C (clk), .D (signal_3402), .Q (signal_3403) ) ;
    buf_clk cell_1866 ( .C (clk), .D (signal_3408), .Q (signal_3409) ) ;
    buf_clk cell_1872 ( .C (clk), .D (signal_3414), .Q (signal_3415) ) ;
    buf_clk cell_1878 ( .C (clk), .D (signal_3420), .Q (signal_3421) ) ;
    buf_clk cell_1884 ( .C (clk), .D (signal_3426), .Q (signal_3427) ) ;
    buf_clk cell_1890 ( .C (clk), .D (signal_3432), .Q (signal_3433) ) ;
    buf_clk cell_1896 ( .C (clk), .D (signal_3438), .Q (signal_3439) ) ;
    buf_clk cell_1902 ( .C (clk), .D (signal_3444), .Q (signal_3445) ) ;
    buf_clk cell_1908 ( .C (clk), .D (signal_3450), .Q (signal_3451) ) ;
    buf_clk cell_1914 ( .C (clk), .D (signal_3456), .Q (signal_3457) ) ;
    buf_clk cell_1920 ( .C (clk), .D (signal_3462), .Q (signal_3463) ) ;
    buf_clk cell_1926 ( .C (clk), .D (signal_3468), .Q (signal_3469) ) ;
    buf_clk cell_1932 ( .C (clk), .D (signal_3474), .Q (signal_3475) ) ;
    buf_clk cell_1938 ( .C (clk), .D (signal_3480), .Q (signal_3481) ) ;
    buf_clk cell_1944 ( .C (clk), .D (signal_3486), .Q (signal_3487) ) ;
    buf_clk cell_1950 ( .C (clk), .D (signal_3492), .Q (signal_3493) ) ;
    buf_clk cell_1956 ( .C (clk), .D (signal_3498), .Q (signal_3499) ) ;
    buf_clk cell_1962 ( .C (clk), .D (signal_3504), .Q (signal_3505) ) ;
    buf_clk cell_1968 ( .C (clk), .D (signal_3510), .Q (signal_3511) ) ;
    buf_clk cell_1974 ( .C (clk), .D (signal_3516), .Q (signal_3517) ) ;
    buf_clk cell_1980 ( .C (clk), .D (signal_3522), .Q (signal_3523) ) ;
    buf_clk cell_1986 ( .C (clk), .D (signal_3528), .Q (signal_3529) ) ;
    buf_clk cell_1992 ( .C (clk), .D (signal_3534), .Q (signal_3535) ) ;
    buf_clk cell_1998 ( .C (clk), .D (signal_3540), .Q (signal_3541) ) ;
    buf_clk cell_2004 ( .C (clk), .D (signal_3546), .Q (signal_3547) ) ;
    buf_clk cell_2010 ( .C (clk), .D (signal_3552), .Q (signal_3553) ) ;
    buf_clk cell_2016 ( .C (clk), .D (signal_3558), .Q (signal_3559) ) ;
    buf_clk cell_2022 ( .C (clk), .D (signal_3564), .Q (signal_3565) ) ;
    buf_clk cell_2028 ( .C (clk), .D (signal_3570), .Q (signal_3571) ) ;
    buf_clk cell_2034 ( .C (clk), .D (signal_3576), .Q (signal_3577) ) ;
    buf_clk cell_2040 ( .C (clk), .D (signal_3582), .Q (signal_3583) ) ;
    buf_clk cell_2046 ( .C (clk), .D (signal_3588), .Q (signal_3589) ) ;
    buf_clk cell_2052 ( .C (clk), .D (signal_3594), .Q (signal_3595) ) ;
    buf_clk cell_2058 ( .C (clk), .D (signal_3600), .Q (signal_3601) ) ;
    buf_clk cell_2064 ( .C (clk), .D (signal_3606), .Q (signal_3607) ) ;
    buf_clk cell_2070 ( .C (clk), .D (signal_3612), .Q (signal_3613) ) ;
    buf_clk cell_2076 ( .C (clk), .D (signal_3618), .Q (signal_3619) ) ;
    buf_clk cell_2082 ( .C (clk), .D (signal_3624), .Q (signal_3625) ) ;
    buf_clk cell_2088 ( .C (clk), .D (signal_3630), .Q (signal_3631) ) ;
    buf_clk cell_2094 ( .C (clk), .D (signal_3636), .Q (signal_3637) ) ;
    buf_clk cell_2100 ( .C (clk), .D (signal_3642), .Q (signal_3643) ) ;
    buf_clk cell_2106 ( .C (clk), .D (signal_3648), .Q (signal_3649) ) ;
    buf_clk cell_2112 ( .C (clk), .D (signal_3654), .Q (signal_3655) ) ;
    buf_clk cell_2118 ( .C (clk), .D (signal_3660), .Q (signal_3661) ) ;
    buf_clk cell_2124 ( .C (clk), .D (signal_3666), .Q (signal_3667) ) ;
    buf_clk cell_2130 ( .C (clk), .D (signal_3672), .Q (signal_3673) ) ;
    buf_clk cell_2136 ( .C (clk), .D (signal_3678), .Q (signal_3679) ) ;
    buf_clk cell_2142 ( .C (clk), .D (signal_3684), .Q (signal_3685) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_3690), .Q (signal_3691) ) ;
    buf_clk cell_2154 ( .C (clk), .D (signal_3696), .Q (signal_3697) ) ;
    buf_clk cell_2160 ( .C (clk), .D (signal_3702), .Q (signal_3703) ) ;
    buf_clk cell_2166 ( .C (clk), .D (signal_3708), .Q (signal_3709) ) ;
    buf_clk cell_2172 ( .C (clk), .D (signal_3714), .Q (signal_3715) ) ;
    buf_clk cell_2178 ( .C (clk), .D (signal_3720), .Q (signal_3721) ) ;
    buf_clk cell_2184 ( .C (clk), .D (signal_3726), .Q (signal_3727) ) ;
    buf_clk cell_2190 ( .C (clk), .D (signal_3732), .Q (signal_3733) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_3738), .Q (signal_3739) ) ;
    buf_clk cell_2202 ( .C (clk), .D (signal_3744), .Q (signal_3745) ) ;
    buf_clk cell_2208 ( .C (clk), .D (signal_3750), .Q (signal_3751) ) ;
    buf_clk cell_2214 ( .C (clk), .D (signal_3756), .Q (signal_3757) ) ;
    buf_clk cell_2220 ( .C (clk), .D (signal_3762), .Q (signal_3763) ) ;
    buf_clk cell_2226 ( .C (clk), .D (signal_3768), .Q (signal_3769) ) ;
    buf_clk cell_2232 ( .C (clk), .D (signal_3774), .Q (signal_3775) ) ;
    buf_clk cell_2238 ( .C (clk), .D (signal_3780), .Q (signal_3781) ) ;
    buf_clk cell_2244 ( .C (clk), .D (signal_3786), .Q (signal_3787) ) ;
    buf_clk cell_2250 ( .C (clk), .D (signal_3792), .Q (signal_3793) ) ;
    buf_clk cell_2256 ( .C (clk), .D (signal_3798), .Q (signal_3799) ) ;
    buf_clk cell_2262 ( .C (clk), .D (signal_3804), .Q (signal_3805) ) ;
    buf_clk cell_2268 ( .C (clk), .D (signal_3810), .Q (signal_3811) ) ;
    buf_clk cell_2274 ( .C (clk), .D (signal_3816), .Q (signal_3817) ) ;
    buf_clk cell_2280 ( .C (clk), .D (signal_3822), .Q (signal_3823) ) ;
    buf_clk cell_2286 ( .C (clk), .D (signal_3828), .Q (signal_3829) ) ;
    buf_clk cell_2292 ( .C (clk), .D (signal_3834), .Q (signal_3835) ) ;
    buf_clk cell_2298 ( .C (clk), .D (signal_3840), .Q (signal_3841) ) ;
    buf_clk cell_2304 ( .C (clk), .D (signal_3846), .Q (signal_3847) ) ;
    buf_clk cell_2310 ( .C (clk), .D (signal_3852), .Q (signal_3853) ) ;
    buf_clk cell_2316 ( .C (clk), .D (signal_3858), .Q (signal_3859) ) ;
    buf_clk cell_2322 ( .C (clk), .D (signal_3864), .Q (signal_3865) ) ;
    buf_clk cell_2328 ( .C (clk), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_2334 ( .C (clk), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_2340 ( .C (clk), .D (signal_3882), .Q (signal_3883) ) ;
    buf_clk cell_2346 ( .C (clk), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_2352 ( .C (clk), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_2358 ( .C (clk), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_2364 ( .C (clk), .D (signal_3906), .Q (signal_3907) ) ;
    buf_clk cell_2370 ( .C (clk), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_2376 ( .C (clk), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_2382 ( .C (clk), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_2388 ( .C (clk), .D (signal_3930), .Q (signal_3931) ) ;
    buf_clk cell_2394 ( .C (clk), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_2400 ( .C (clk), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_2406 ( .C (clk), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_2412 ( .C (clk), .D (signal_3954), .Q (signal_3955) ) ;
    buf_clk cell_2418 ( .C (clk), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_2424 ( .C (clk), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_2430 ( .C (clk), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_2436 ( .C (clk), .D (signal_3978), .Q (signal_3979) ) ;
    buf_clk cell_2442 ( .C (clk), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_2448 ( .C (clk), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_2454 ( .C (clk), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_2460 ( .C (clk), .D (signal_4002), .Q (signal_4003) ) ;
    buf_clk cell_2466 ( .C (clk), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_2472 ( .C (clk), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_2478 ( .C (clk), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_2484 ( .C (clk), .D (signal_4026), .Q (signal_4027) ) ;
    buf_clk cell_2490 ( .C (clk), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_2496 ( .C (clk), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_2502 ( .C (clk), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_2508 ( .C (clk), .D (signal_4050), .Q (signal_4051) ) ;
    buf_clk cell_2514 ( .C (clk), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_2520 ( .C (clk), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_2526 ( .C (clk), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_2532 ( .C (clk), .D (signal_4074), .Q (signal_4075) ) ;
    buf_clk cell_2538 ( .C (clk), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_2544 ( .C (clk), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_2550 ( .C (clk), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_2556 ( .C (clk), .D (signal_4098), .Q (signal_4099) ) ;
    buf_clk cell_2562 ( .C (clk), .D (signal_4104), .Q (signal_4105) ) ;
    buf_clk cell_2568 ( .C (clk), .D (signal_4110), .Q (signal_4111) ) ;
    buf_clk cell_2574 ( .C (clk), .D (signal_4116), .Q (signal_4117) ) ;
    buf_clk cell_2580 ( .C (clk), .D (signal_4122), .Q (signal_4123) ) ;
    buf_clk cell_2586 ( .C (clk), .D (signal_4128), .Q (signal_4129) ) ;
    buf_clk cell_2592 ( .C (clk), .D (signal_4134), .Q (signal_4135) ) ;
    buf_clk cell_2598 ( .C (clk), .D (signal_4140), .Q (signal_4141) ) ;
    buf_clk cell_2604 ( .C (clk), .D (signal_4146), .Q (signal_4147) ) ;
    buf_clk cell_2610 ( .C (clk), .D (signal_4152), .Q (signal_4153) ) ;
    buf_clk cell_2616 ( .C (clk), .D (signal_4158), .Q (signal_4159) ) ;
    buf_clk cell_2622 ( .C (clk), .D (signal_4164), .Q (signal_4165) ) ;
    buf_clk cell_2628 ( .C (clk), .D (signal_4170), .Q (signal_4171) ) ;
    buf_clk cell_2634 ( .C (clk), .D (signal_4176), .Q (signal_4177) ) ;
    buf_clk cell_2640 ( .C (clk), .D (signal_4182), .Q (signal_4183) ) ;
    buf_clk cell_2646 ( .C (clk), .D (signal_4188), .Q (signal_4189) ) ;
    buf_clk cell_2652 ( .C (clk), .D (signal_4194), .Q (signal_4195) ) ;
    buf_clk cell_2658 ( .C (clk), .D (signal_4200), .Q (signal_4201) ) ;
    buf_clk cell_2664 ( .C (clk), .D (signal_4206), .Q (signal_4207) ) ;
    buf_clk cell_2670 ( .C (clk), .D (signal_4212), .Q (signal_4213) ) ;
    buf_clk cell_2676 ( .C (clk), .D (signal_4218), .Q (signal_4219) ) ;
    buf_clk cell_2682 ( .C (clk), .D (signal_4224), .Q (signal_4225) ) ;
    buf_clk cell_2688 ( .C (clk), .D (signal_4230), .Q (signal_4231) ) ;
    buf_clk cell_2694 ( .C (clk), .D (signal_4236), .Q (signal_4237) ) ;
    buf_clk cell_2700 ( .C (clk), .D (signal_4242), .Q (signal_4243) ) ;
    buf_clk cell_2706 ( .C (clk), .D (signal_4248), .Q (signal_4249) ) ;
    buf_clk cell_2712 ( .C (clk), .D (signal_4254), .Q (signal_4255) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_4260), .Q (signal_4261) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_4266), .Q (signal_4267) ) ;
    buf_clk cell_2730 ( .C (clk), .D (signal_4272), .Q (signal_4273) ) ;
    buf_clk cell_2736 ( .C (clk), .D (signal_4278), .Q (signal_4279) ) ;
    buf_clk cell_2742 ( .C (clk), .D (signal_4284), .Q (signal_4285) ) ;
    buf_clk cell_2748 ( .C (clk), .D (signal_4290), .Q (signal_4291) ) ;
    buf_clk cell_2754 ( .C (clk), .D (signal_4296), .Q (signal_4297) ) ;
    buf_clk cell_2760 ( .C (clk), .D (signal_4302), .Q (signal_4303) ) ;
    buf_clk cell_2766 ( .C (clk), .D (signal_4308), .Q (signal_4309) ) ;
    buf_clk cell_2772 ( .C (clk), .D (signal_4314), .Q (signal_4315) ) ;
    buf_clk cell_2778 ( .C (clk), .D (signal_4320), .Q (signal_4321) ) ;
    buf_clk cell_2784 ( .C (clk), .D (signal_4326), .Q (signal_4327) ) ;
    buf_clk cell_2790 ( .C (clk), .D (signal_4332), .Q (signal_4333) ) ;
    buf_clk cell_2796 ( .C (clk), .D (signal_4338), .Q (signal_4339) ) ;
    buf_clk cell_2802 ( .C (clk), .D (signal_4344), .Q (signal_4345) ) ;
    buf_clk cell_2808 ( .C (clk), .D (signal_4350), .Q (signal_4351) ) ;
    buf_clk cell_2814 ( .C (clk), .D (signal_4356), .Q (signal_4357) ) ;
    buf_clk cell_2820 ( .C (clk), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_2826 ( .C (clk), .D (signal_4368), .Q (signal_4369) ) ;
    buf_clk cell_2832 ( .C (clk), .D (signal_4374), .Q (signal_4375) ) ;
    buf_clk cell_2838 ( .C (clk), .D (signal_4380), .Q (signal_4381) ) ;
    buf_clk cell_2844 ( .C (clk), .D (signal_4386), .Q (signal_4387) ) ;
    buf_clk cell_2850 ( .C (clk), .D (signal_4392), .Q (signal_4393) ) ;
    buf_clk cell_2856 ( .C (clk), .D (signal_4398), .Q (signal_4399) ) ;
    buf_clk cell_2862 ( .C (clk), .D (signal_4404), .Q (signal_4405) ) ;
    buf_clk cell_2868 ( .C (clk), .D (signal_4410), .Q (signal_4411) ) ;
    buf_clk cell_2874 ( .C (clk), .D (signal_4416), .Q (signal_4417) ) ;
    buf_clk cell_2880 ( .C (clk), .D (signal_4422), .Q (signal_4423) ) ;
    buf_clk cell_2886 ( .C (clk), .D (signal_4428), .Q (signal_4429) ) ;
    buf_clk cell_2892 ( .C (clk), .D (signal_4434), .Q (signal_4435) ) ;
    buf_clk cell_2898 ( .C (clk), .D (signal_4440), .Q (signal_4441) ) ;
    buf_clk cell_2904 ( .C (clk), .D (signal_4446), .Q (signal_4447) ) ;
    buf_clk cell_2910 ( .C (clk), .D (signal_4452), .Q (signal_4453) ) ;
    buf_clk cell_2914 ( .C (clk), .D (signal_3250), .Q (signal_4457) ) ;
    buf_clk cell_2916 ( .C (clk), .D (signal_3252), .Q (signal_4459) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_4462), .Q (signal_4463) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_4466), .Q (signal_4467) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_3290), .Q (signal_4469) ) ;
    buf_clk cell_2928 ( .C (clk), .D (signal_3292), .Q (signal_4471) ) ;
    buf_clk cell_2930 ( .C (clk), .D (signal_3182), .Q (signal_4473) ) ;
    buf_clk cell_2932 ( .C (clk), .D (signal_3184), .Q (signal_4475) ) ;
    buf_clk cell_2934 ( .C (clk), .D (signal_3222), .Q (signal_4477) ) ;
    buf_clk cell_2936 ( .C (clk), .D (signal_3224), .Q (signal_4479) ) ;
    buf_clk cell_2938 ( .C (clk), .D (signal_3214), .Q (signal_4481) ) ;
    buf_clk cell_2940 ( .C (clk), .D (signal_3216), .Q (signal_4483) ) ;
    buf_clk cell_2942 ( .C (clk), .D (signal_3246), .Q (signal_4485) ) ;
    buf_clk cell_2944 ( .C (clk), .D (signal_3248), .Q (signal_4487) ) ;
    buf_clk cell_2946 ( .C (clk), .D (signal_3230), .Q (signal_4489) ) ;
    buf_clk cell_2948 ( .C (clk), .D (signal_3232), .Q (signal_4491) ) ;
    buf_clk cell_2950 ( .C (clk), .D (signal_3238), .Q (signal_4493) ) ;
    buf_clk cell_2952 ( .C (clk), .D (signal_3240), .Q (signal_4495) ) ;
    buf_clk cell_2956 ( .C (clk), .D (signal_4498), .Q (signal_4499) ) ;
    buf_clk cell_2960 ( .C (clk), .D (signal_4502), .Q (signal_4503) ) ;
    buf_clk cell_2964 ( .C (clk), .D (signal_4506), .Q (signal_4507) ) ;
    buf_clk cell_2968 ( .C (clk), .D (signal_4510), .Q (signal_4511) ) ;
    buf_clk cell_2970 ( .C (clk), .D (signal_3242), .Q (signal_4513) ) ;
    buf_clk cell_2972 ( .C (clk), .D (signal_3244), .Q (signal_4515) ) ;
    buf_clk cell_2976 ( .C (clk), .D (signal_4518), .Q (signal_4519) ) ;
    buf_clk cell_2980 ( .C (clk), .D (signal_4522), .Q (signal_4523) ) ;
    buf_clk cell_2984 ( .C (clk), .D (signal_4526), .Q (signal_4527) ) ;
    buf_clk cell_2988 ( .C (clk), .D (signal_4530), .Q (signal_4531) ) ;
    buf_clk cell_2992 ( .C (clk), .D (signal_4534), .Q (signal_4535) ) ;
    buf_clk cell_2996 ( .C (clk), .D (signal_4538), .Q (signal_4539) ) ;
    buf_clk cell_2998 ( .C (clk), .D (signal_3210), .Q (signal_4541) ) ;
    buf_clk cell_3000 ( .C (clk), .D (signal_3212), .Q (signal_4543) ) ;
    buf_clk cell_3004 ( .C (clk), .D (signal_4546), .Q (signal_4547) ) ;
    buf_clk cell_3008 ( .C (clk), .D (signal_4550), .Q (signal_4551) ) ;
    buf_clk cell_3012 ( .C (clk), .D (signal_4554), .Q (signal_4555) ) ;
    buf_clk cell_3016 ( .C (clk), .D (signal_4558), .Q (signal_4559) ) ;
    buf_clk cell_3020 ( .C (clk), .D (signal_4562), .Q (signal_4563) ) ;
    buf_clk cell_3024 ( .C (clk), .D (signal_4566), .Q (signal_4567) ) ;
    buf_clk cell_3028 ( .C (clk), .D (signal_4570), .Q (signal_4571) ) ;
    buf_clk cell_3032 ( .C (clk), .D (signal_4574), .Q (signal_4575) ) ;
    buf_clk cell_3036 ( .C (clk), .D (signal_4578), .Q (signal_4579) ) ;
    buf_clk cell_3040 ( .C (clk), .D (signal_4582), .Q (signal_4583) ) ;
    buf_clk cell_3042 ( .C (clk), .D (signal_3234), .Q (signal_4585) ) ;
    buf_clk cell_3044 ( .C (clk), .D (signal_3236), .Q (signal_4587) ) ;
    buf_clk cell_3046 ( .C (clk), .D (signal_3218), .Q (signal_4589) ) ;
    buf_clk cell_3048 ( .C (clk), .D (signal_3220), .Q (signal_4591) ) ;
    buf_clk cell_3052 ( .C (clk), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_3056 ( .C (clk), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_3058 ( .C (clk), .D (signal_3258), .Q (signal_4601) ) ;
    buf_clk cell_3060 ( .C (clk), .D (signal_3260), .Q (signal_4603) ) ;
    buf_clk cell_3064 ( .C (clk), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_3068 ( .C (clk), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_3070 ( .C (clk), .D (signal_3266), .Q (signal_4613) ) ;
    buf_clk cell_3072 ( .C (clk), .D (signal_3268), .Q (signal_4615) ) ;
    buf_clk cell_3076 ( .C (clk), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_3080 ( .C (clk), .D (signal_4622), .Q (signal_4623) ) ;
    buf_clk cell_3082 ( .C (clk), .D (signal_3274), .Q (signal_4625) ) ;
    buf_clk cell_3084 ( .C (clk), .D (signal_3276), .Q (signal_4627) ) ;
    buf_clk cell_3088 ( .C (clk), .D (signal_4630), .Q (signal_4631) ) ;
    buf_clk cell_3092 ( .C (clk), .D (signal_4634), .Q (signal_4635) ) ;
    buf_clk cell_3094 ( .C (clk), .D (signal_3282), .Q (signal_4637) ) ;
    buf_clk cell_3096 ( .C (clk), .D (signal_3284), .Q (signal_4639) ) ;
    buf_clk cell_3100 ( .C (clk), .D (signal_4642), .Q (signal_4643) ) ;
    buf_clk cell_3104 ( .C (clk), .D (signal_4646), .Q (signal_4647) ) ;
    buf_clk cell_3108 ( .C (clk), .D (signal_4650), .Q (signal_4651) ) ;
    buf_clk cell_3116 ( .C (clk), .D (signal_4658), .Q (signal_4659) ) ;
    buf_clk cell_3124 ( .C (clk), .D (signal_4666), .Q (signal_4667) ) ;
    buf_clk cell_3132 ( .C (clk), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_3140 ( .C (clk), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_3148 ( .C (clk), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_3156 ( .C (clk), .D (signal_4698), .Q (signal_4699) ) ;
    buf_clk cell_3164 ( .C (clk), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_3172 ( .C (clk), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_3180 ( .C (clk), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_3188 ( .C (clk), .D (signal_4730), .Q (signal_4731) ) ;
    buf_clk cell_3196 ( .C (clk), .D (signal_4738), .Q (signal_4739) ) ;
    buf_clk cell_3204 ( .C (clk), .D (signal_4746), .Q (signal_4747) ) ;
    buf_clk cell_3212 ( .C (clk), .D (signal_4754), .Q (signal_4755) ) ;
    buf_clk cell_3220 ( .C (clk), .D (signal_4762), .Q (signal_4763) ) ;
    buf_clk cell_3228 ( .C (clk), .D (signal_4770), .Q (signal_4771) ) ;
    buf_clk cell_3236 ( .C (clk), .D (signal_4778), .Q (signal_4779) ) ;
    buf_clk cell_3244 ( .C (clk), .D (signal_4786), .Q (signal_4787) ) ;
    buf_clk cell_3252 ( .C (clk), .D (signal_4794), .Q (signal_4795) ) ;
    buf_clk cell_3260 ( .C (clk), .D (signal_4802), .Q (signal_4803) ) ;
    buf_clk cell_3268 ( .C (clk), .D (signal_4810), .Q (signal_4811) ) ;
    buf_clk cell_3276 ( .C (clk), .D (signal_4818), .Q (signal_4819) ) ;
    buf_clk cell_3284 ( .C (clk), .D (signal_4826), .Q (signal_4827) ) ;
    buf_clk cell_3292 ( .C (clk), .D (signal_4834), .Q (signal_4835) ) ;
    buf_clk cell_3300 ( .C (clk), .D (signal_4842), .Q (signal_4843) ) ;
    buf_clk cell_3308 ( .C (clk), .D (signal_4850), .Q (signal_4851) ) ;
    buf_clk cell_3316 ( .C (clk), .D (signal_4858), .Q (signal_4859) ) ;
    buf_clk cell_3324 ( .C (clk), .D (signal_4866), .Q (signal_4867) ) ;
    buf_clk cell_3332 ( .C (clk), .D (signal_4874), .Q (signal_4875) ) ;
    buf_clk cell_3340 ( .C (clk), .D (signal_4882), .Q (signal_4883) ) ;
    buf_clk cell_3348 ( .C (clk), .D (signal_4890), .Q (signal_4891) ) ;
    buf_clk cell_3356 ( .C (clk), .D (signal_4898), .Q (signal_4899) ) ;
    buf_clk cell_3364 ( .C (clk), .D (signal_4906), .Q (signal_4907) ) ;
    buf_clk cell_3372 ( .C (clk), .D (signal_4914), .Q (signal_4915) ) ;
    buf_clk cell_3380 ( .C (clk), .D (signal_4922), .Q (signal_4923) ) ;
    buf_clk cell_3388 ( .C (clk), .D (signal_4930), .Q (signal_4931) ) ;
    buf_clk cell_3396 ( .C (clk), .D (signal_4938), .Q (signal_4939) ) ;
    buf_clk cell_3404 ( .C (clk), .D (signal_4946), .Q (signal_4947) ) ;
    buf_clk cell_3412 ( .C (clk), .D (signal_4954), .Q (signal_4955) ) ;
    buf_clk cell_3420 ( .C (clk), .D (signal_4962), .Q (signal_4963) ) ;
    buf_clk cell_3428 ( .C (clk), .D (signal_4970), .Q (signal_4971) ) ;
    buf_clk cell_3436 ( .C (clk), .D (signal_4978), .Q (signal_4979) ) ;
    buf_clk cell_3444 ( .C (clk), .D (signal_4986), .Q (signal_4987) ) ;
    buf_clk cell_3452 ( .C (clk), .D (signal_4994), .Q (signal_4995) ) ;
    buf_clk cell_3460 ( .C (clk), .D (signal_5002), .Q (signal_5003) ) ;
    buf_clk cell_3468 ( .C (clk), .D (signal_5010), .Q (signal_5011) ) ;
    buf_clk cell_3476 ( .C (clk), .D (signal_5018), .Q (signal_5019) ) ;
    buf_clk cell_3484 ( .C (clk), .D (signal_5026), .Q (signal_5027) ) ;
    buf_clk cell_3492 ( .C (clk), .D (signal_5034), .Q (signal_5035) ) ;
    buf_clk cell_3500 ( .C (clk), .D (signal_5042), .Q (signal_5043) ) ;
    buf_clk cell_3508 ( .C (clk), .D (signal_5050), .Q (signal_5051) ) ;
    buf_clk cell_3516 ( .C (clk), .D (signal_5058), .Q (signal_5059) ) ;
    buf_clk cell_3524 ( .C (clk), .D (signal_5066), .Q (signal_5067) ) ;
    buf_clk cell_3532 ( .C (clk), .D (signal_5074), .Q (signal_5075) ) ;
    buf_clk cell_3540 ( .C (clk), .D (signal_5082), .Q (signal_5083) ) ;
    buf_clk cell_3548 ( .C (clk), .D (signal_5090), .Q (signal_5091) ) ;
    buf_clk cell_3556 ( .C (clk), .D (signal_5098), .Q (signal_5099) ) ;
    buf_clk cell_3564 ( .C (clk), .D (signal_5106), .Q (signal_5107) ) ;
    buf_clk cell_3572 ( .C (clk), .D (signal_5114), .Q (signal_5115) ) ;
    buf_clk cell_3580 ( .C (clk), .D (signal_5122), .Q (signal_5123) ) ;
    buf_clk cell_3588 ( .C (clk), .D (signal_5130), .Q (signal_5131) ) ;
    buf_clk cell_3596 ( .C (clk), .D (signal_5138), .Q (signal_5139) ) ;
    buf_clk cell_3604 ( .C (clk), .D (signal_5146), .Q (signal_5147) ) ;
    buf_clk cell_3612 ( .C (clk), .D (signal_5154), .Q (signal_5155) ) ;
    buf_clk cell_3620 ( .C (clk), .D (signal_5162), .Q (signal_5163) ) ;
    buf_clk cell_3628 ( .C (clk), .D (signal_5170), .Q (signal_5171) ) ;
    buf_clk cell_3636 ( .C (clk), .D (signal_5178), .Q (signal_5179) ) ;
    buf_clk cell_3644 ( .C (clk), .D (signal_5186), .Q (signal_5187) ) ;
    buf_clk cell_3652 ( .C (clk), .D (signal_5194), .Q (signal_5195) ) ;
    buf_clk cell_3660 ( .C (clk), .D (signal_5202), .Q (signal_5203) ) ;
    buf_clk cell_3668 ( .C (clk), .D (signal_5210), .Q (signal_5211) ) ;
    buf_clk cell_3676 ( .C (clk), .D (signal_5218), .Q (signal_5219) ) ;
    buf_clk cell_3684 ( .C (clk), .D (signal_5226), .Q (signal_5227) ) ;
    buf_clk cell_3692 ( .C (clk), .D (signal_5234), .Q (signal_5235) ) ;
    buf_clk cell_3700 ( .C (clk), .D (signal_5242), .Q (signal_5243) ) ;
    buf_clk cell_3708 ( .C (clk), .D (signal_5250), .Q (signal_5251) ) ;
    buf_clk cell_3716 ( .C (clk), .D (signal_5258), .Q (signal_5259) ) ;
    buf_clk cell_3724 ( .C (clk), .D (signal_5266), .Q (signal_5267) ) ;
    buf_clk cell_3732 ( .C (clk), .D (signal_5274), .Q (signal_5275) ) ;
    buf_clk cell_3740 ( .C (clk), .D (signal_5282), .Q (signal_5283) ) ;
    buf_clk cell_3748 ( .C (clk), .D (signal_5290), .Q (signal_5291) ) ;
    buf_clk cell_3756 ( .C (clk), .D (signal_5298), .Q (signal_5299) ) ;
    buf_clk cell_3764 ( .C (clk), .D (signal_5306), .Q (signal_5307) ) ;
    buf_clk cell_3772 ( .C (clk), .D (signal_5314), .Q (signal_5315) ) ;
    buf_clk cell_3780 ( .C (clk), .D (signal_5322), .Q (signal_5323) ) ;
    buf_clk cell_3788 ( .C (clk), .D (signal_5330), .Q (signal_5331) ) ;
    buf_clk cell_3796 ( .C (clk), .D (signal_5338), .Q (signal_5339) ) ;
    buf_clk cell_3804 ( .C (clk), .D (signal_5346), .Q (signal_5347) ) ;
    buf_clk cell_3812 ( .C (clk), .D (signal_5354), .Q (signal_5355) ) ;
    buf_clk cell_3820 ( .C (clk), .D (signal_5362), .Q (signal_5363) ) ;
    buf_clk cell_3828 ( .C (clk), .D (signal_5370), .Q (signal_5371) ) ;
    buf_clk cell_3836 ( .C (clk), .D (signal_5378), .Q (signal_5379) ) ;
    buf_clk cell_3844 ( .C (clk), .D (signal_5386), .Q (signal_5387) ) ;
    buf_clk cell_3852 ( .C (clk), .D (signal_5394), .Q (signal_5395) ) ;
    buf_clk cell_3860 ( .C (clk), .D (signal_5402), .Q (signal_5403) ) ;
    buf_clk cell_3868 ( .C (clk), .D (signal_5410), .Q (signal_5411) ) ;
    buf_clk cell_3876 ( .C (clk), .D (signal_5418), .Q (signal_5419) ) ;
    buf_clk cell_3884 ( .C (clk), .D (signal_5426), .Q (signal_5427) ) ;
    buf_clk cell_3892 ( .C (clk), .D (signal_5434), .Q (signal_5435) ) ;
    buf_clk cell_3900 ( .C (clk), .D (signal_5442), .Q (signal_5443) ) ;
    buf_clk cell_3908 ( .C (clk), .D (signal_5450), .Q (signal_5451) ) ;
    buf_clk cell_3916 ( .C (clk), .D (signal_5458), .Q (signal_5459) ) ;
    buf_clk cell_3924 ( .C (clk), .D (signal_5466), .Q (signal_5467) ) ;
    buf_clk cell_3932 ( .C (clk), .D (signal_5474), .Q (signal_5475) ) ;
    buf_clk cell_3940 ( .C (clk), .D (signal_5482), .Q (signal_5483) ) ;
    buf_clk cell_3948 ( .C (clk), .D (signal_5490), .Q (signal_5491) ) ;
    buf_clk cell_3956 ( .C (clk), .D (signal_5498), .Q (signal_5499) ) ;
    buf_clk cell_3964 ( .C (clk), .D (signal_5506), .Q (signal_5507) ) ;
    buf_clk cell_3972 ( .C (clk), .D (signal_5514), .Q (signal_5515) ) ;
    buf_clk cell_3980 ( .C (clk), .D (signal_5522), .Q (signal_5523) ) ;
    buf_clk cell_3988 ( .C (clk), .D (signal_5530), .Q (signal_5531) ) ;
    buf_clk cell_3996 ( .C (clk), .D (signal_5538), .Q (signal_5539) ) ;
    buf_clk cell_4004 ( .C (clk), .D (signal_5546), .Q (signal_5547) ) ;
    buf_clk cell_4012 ( .C (clk), .D (signal_5554), .Q (signal_5555) ) ;
    buf_clk cell_4020 ( .C (clk), .D (signal_5562), .Q (signal_5563) ) ;
    buf_clk cell_4028 ( .C (clk), .D (signal_5570), .Q (signal_5571) ) ;
    buf_clk cell_4036 ( .C (clk), .D (signal_5578), .Q (signal_5579) ) ;
    buf_clk cell_4044 ( .C (clk), .D (signal_5586), .Q (signal_5587) ) ;
    buf_clk cell_4052 ( .C (clk), .D (signal_5594), .Q (signal_5595) ) ;
    buf_clk cell_4060 ( .C (clk), .D (signal_5602), .Q (signal_5603) ) ;
    buf_clk cell_4068 ( .C (clk), .D (signal_5610), .Q (signal_5611) ) ;
    buf_clk cell_4076 ( .C (clk), .D (signal_5618), .Q (signal_5619) ) ;
    buf_clk cell_4084 ( .C (clk), .D (signal_5626), .Q (signal_5627) ) ;
    buf_clk cell_4092 ( .C (clk), .D (signal_5634), .Q (signal_5635) ) ;
    buf_clk cell_4100 ( .C (clk), .D (signal_5642), .Q (signal_5643) ) ;
    buf_clk cell_4108 ( .C (clk), .D (signal_5650), .Q (signal_5651) ) ;
    buf_clk cell_4116 ( .C (clk), .D (signal_5658), .Q (signal_5659) ) ;
    buf_clk cell_4124 ( .C (clk), .D (signal_5666), .Q (signal_5667) ) ;
    buf_clk cell_4134 ( .C (clk), .D (signal_5676), .Q (signal_5677) ) ;
    buf_clk cell_4142 ( .C (clk), .D (signal_5684), .Q (signal_5685) ) ;
    buf_clk cell_4150 ( .C (clk), .D (signal_5692), .Q (signal_5693) ) ;
    buf_clk cell_4158 ( .C (clk), .D (signal_5700), .Q (signal_5701) ) ;
    buf_clk cell_4166 ( .C (clk), .D (signal_5708), .Q (signal_5709) ) ;
    buf_clk cell_4174 ( .C (clk), .D (signal_5716), .Q (signal_5717) ) ;
    buf_clk cell_4182 ( .C (clk), .D (signal_5724), .Q (signal_5725) ) ;
    buf_clk cell_4190 ( .C (clk), .D (signal_5732), .Q (signal_5733) ) ;
    buf_clk cell_4198 ( .C (clk), .D (signal_5740), .Q (signal_5741) ) ;
    buf_clk cell_4206 ( .C (clk), .D (signal_5748), .Q (signal_5749) ) ;
    buf_clk cell_4214 ( .C (clk), .D (signal_5756), .Q (signal_5757) ) ;
    buf_clk cell_4222 ( .C (clk), .D (signal_5764), .Q (signal_5765) ) ;
    buf_clk cell_4230 ( .C (clk), .D (signal_5772), .Q (signal_5773) ) ;
    buf_clk cell_4238 ( .C (clk), .D (signal_5780), .Q (signal_5781) ) ;
    buf_clk cell_4246 ( .C (clk), .D (signal_5788), .Q (signal_5789) ) ;
    buf_clk cell_4254 ( .C (clk), .D (signal_5796), .Q (signal_5797) ) ;
    buf_clk cell_4262 ( .C (clk), .D (signal_5804), .Q (signal_5805) ) ;
    buf_clk cell_4270 ( .C (clk), .D (signal_5812), .Q (signal_5813) ) ;
    buf_clk cell_4278 ( .C (clk), .D (signal_5820), .Q (signal_5821) ) ;
    buf_clk cell_4286 ( .C (clk), .D (signal_5828), .Q (signal_5829) ) ;
    buf_clk cell_4294 ( .C (clk), .D (signal_5836), .Q (signal_5837) ) ;
    buf_clk cell_4302 ( .C (clk), .D (signal_5844), .Q (signal_5845) ) ;
    buf_clk cell_4310 ( .C (clk), .D (signal_5852), .Q (signal_5853) ) ;
    buf_clk cell_4318 ( .C (clk), .D (signal_5860), .Q (signal_5861) ) ;
    buf_clk cell_4326 ( .C (clk), .D (signal_5868), .Q (signal_5869) ) ;
    buf_clk cell_4334 ( .C (clk), .D (signal_5876), .Q (signal_5877) ) ;
    buf_clk cell_4342 ( .C (clk), .D (signal_5884), .Q (signal_5885) ) ;
    buf_clk cell_4350 ( .C (clk), .D (signal_5892), .Q (signal_5893) ) ;
    buf_clk cell_4358 ( .C (clk), .D (signal_5900), .Q (signal_5901) ) ;
    buf_clk cell_4366 ( .C (clk), .D (signal_5908), .Q (signal_5909) ) ;
    buf_clk cell_4374 ( .C (clk), .D (signal_5916), .Q (signal_5917) ) ;
    buf_clk cell_4382 ( .C (clk), .D (signal_5924), .Q (signal_5925) ) ;
    buf_clk cell_4390 ( .C (clk), .D (signal_5932), .Q (signal_5933) ) ;
    buf_clk cell_4398 ( .C (clk), .D (signal_5940), .Q (signal_5941) ) ;
    buf_clk cell_4406 ( .C (clk), .D (signal_5948), .Q (signal_5949) ) ;
    buf_clk cell_4414 ( .C (clk), .D (signal_5956), .Q (signal_5957) ) ;
    buf_clk cell_4422 ( .C (clk), .D (signal_5964), .Q (signal_5965) ) ;
    buf_clk cell_4430 ( .C (clk), .D (signal_5972), .Q (signal_5973) ) ;
    buf_clk cell_4438 ( .C (clk), .D (signal_5980), .Q (signal_5981) ) ;
    buf_clk cell_4446 ( .C (clk), .D (signal_5988), .Q (signal_5989) ) ;
    buf_clk cell_4454 ( .C (clk), .D (signal_5996), .Q (signal_5997) ) ;
    buf_clk cell_4462 ( .C (clk), .D (signal_6004), .Q (signal_6005) ) ;
    buf_clk cell_4470 ( .C (clk), .D (signal_6012), .Q (signal_6013) ) ;
    buf_clk cell_4478 ( .C (clk), .D (signal_6020), .Q (signal_6021) ) ;
    buf_clk cell_4486 ( .C (clk), .D (signal_6028), .Q (signal_6029) ) ;
    buf_clk cell_4494 ( .C (clk), .D (signal_6036), .Q (signal_6037) ) ;
    buf_clk cell_4502 ( .C (clk), .D (signal_6044), .Q (signal_6045) ) ;
    buf_clk cell_4510 ( .C (clk), .D (signal_6052), .Q (signal_6053) ) ;
    buf_clk cell_4518 ( .C (clk), .D (signal_6060), .Q (signal_6061) ) ;
    buf_clk cell_4526 ( .C (clk), .D (signal_6068), .Q (signal_6069) ) ;
    buf_clk cell_4534 ( .C (clk), .D (signal_6076), .Q (signal_6077) ) ;
    buf_clk cell_4542 ( .C (clk), .D (signal_6084), .Q (signal_6085) ) ;
    buf_clk cell_4550 ( .C (clk), .D (signal_6092), .Q (signal_6093) ) ;
    buf_clk cell_4558 ( .C (clk), .D (signal_6100), .Q (signal_6101) ) ;
    buf_clk cell_4566 ( .C (clk), .D (signal_6108), .Q (signal_6109) ) ;
    buf_clk cell_4574 ( .C (clk), .D (signal_6116), .Q (signal_6117) ) ;
    buf_clk cell_4582 ( .C (clk), .D (signal_6124), .Q (signal_6125) ) ;
    buf_clk cell_4590 ( .C (clk), .D (signal_6132), .Q (signal_6133) ) ;
    buf_clk cell_4598 ( .C (clk), .D (signal_6140), .Q (signal_6141) ) ;
    buf_clk cell_4606 ( .C (clk), .D (signal_6148), .Q (signal_6149) ) ;
    buf_clk cell_4614 ( .C (clk), .D (signal_6156), .Q (signal_6157) ) ;
    buf_clk cell_4622 ( .C (clk), .D (signal_6164), .Q (signal_6165) ) ;
    buf_clk cell_4630 ( .C (clk), .D (signal_6172), .Q (signal_6173) ) ;
    buf_clk cell_4638 ( .C (clk), .D (signal_6180), .Q (signal_6181) ) ;
    buf_clk cell_4840 ( .C (clk), .D (signal_6382), .Q (signal_6383) ) ;
    buf_clk cell_4848 ( .C (clk), .D (signal_6390), .Q (signal_6391) ) ;
    buf_clk cell_4856 ( .C (clk), .D (signal_6398), .Q (signal_6399) ) ;
    buf_clk cell_4864 ( .C (clk), .D (signal_6406), .Q (signal_6407) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1294 ( .s ({signal_3168, signal_3166}), .b ({signal_1849, signal_1468}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[39]), .c ({signal_2019, signal_1495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1295 ( .s ({signal_3172, signal_3170}), .b ({1'b0, 1'b1}), .a ({signal_1842, signal_1463}), .clk (clk), .r (Fresh[40]), .c ({signal_2020, signal_1496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1296 ( .s ({signal_3176, signal_3174}), .b ({1'b0, 1'b1}), .a ({signal_1837, signal_1460}), .clk (clk), .r (Fresh[41]), .c ({signal_2021, signal_1497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1297 ( .s ({signal_3180, signal_3178}), .b ({1'b0, 1'b0}), .a ({signal_1865, signal_1479}), .clk (clk), .r (Fresh[42]), .c ({signal_2023, signal_1498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1298 ( .s ({signal_3184, signal_3182}), .b ({signal_1851, signal_1469}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[43]), .c ({signal_2025, signal_1499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1299 ( .s ({signal_3188, signal_3186}), .b ({1'b0, 1'b0}), .a ({signal_1863, signal_1477}), .clk (clk), .r (Fresh[44]), .c ({signal_2027, signal_1500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1300 ( .s ({signal_3180, signal_3178}), .b ({signal_1857, signal_1473}), .a ({signal_1865, signal_1479}), .clk (clk), .r (Fresh[45]), .c ({signal_2028, signal_1501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1301 ( .s ({signal_3168, signal_3166}), .b ({1'b0, 1'b0}), .a ({signal_1844, signal_1464}), .clk (clk), .r (Fresh[46]), .c ({signal_2029, signal_1502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1302 ( .s ({signal_3192, signal_3190}), .b ({signal_1859, signal_1475}), .a ({signal_1851, signal_1469}), .clk (clk), .r (Fresh[47]), .c ({signal_2031, signal_1503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1303 ( .s ({signal_3196, signal_3194}), .b ({1'b0, 1'b1}), .a ({signal_1840, signal_1462}), .clk (clk), .r (Fresh[48]), .c ({signal_2032, signal_1504}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1304 ( .s ({signal_3200, signal_3198}), .b ({signal_1853, signal_1471}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[49]), .c ({signal_2034, signal_1505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1305 ( .s ({signal_3204, signal_3202}), .b ({1'b0, 1'b0}), .a ({signal_1866, signal_1480}), .clk (clk), .r (Fresh[50]), .c ({signal_2036, signal_1506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1306 ( .s ({signal_3180, signal_3178}), .b ({signal_1865, signal_1479}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[51]), .c ({signal_2037, signal_1507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1307 ( .s ({signal_3208, signal_3206}), .b ({signal_1852, signal_1470}), .a ({signal_1833, signal_1458}), .clk (clk), .r (Fresh[52]), .c ({signal_2039, signal_1508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1308 ( .s ({signal_3208, signal_3206}), .b ({signal_1833, signal_1458}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[53]), .c ({signal_2040, signal_1509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1309 ( .s ({signal_3204, signal_3202}), .b ({signal_1866, signal_1480}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[54]), .c ({signal_2041, signal_1510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1310 ( .s ({signal_3168, signal_3166}), .b ({signal_1849, signal_1468}), .a ({signal_1844, signal_1464}), .clk (clk), .r (Fresh[55]), .c ({signal_2042, signal_1511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1311 ( .s ({signal_3212, signal_3210}), .b ({signal_1858, signal_1474}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[56]), .c ({signal_2044, signal_1512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1312 ( .s ({signal_3216, signal_3214}), .b ({signal_1833, signal_1458}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[57]), .c ({signal_2046, signal_1513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1313 ( .s ({signal_3196, signal_3194}), .b ({signal_1840, signal_1462}), .a ({signal_1845, signal_1465}), .clk (clk), .r (Fresh[58]), .c ({signal_2047, signal_1514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1314 ( .s ({signal_3176, signal_3174}), .b ({signal_1837, signal_1460}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[59]), .c ({signal_2048, signal_1515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1315 ( .s ({signal_3176, signal_3174}), .b ({signal_1837, signal_1460}), .a ({signal_1838, signal_1461}), .clk (clk), .r (Fresh[60]), .c ({signal_2049, signal_1516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1316 ( .s ({signal_3208, signal_3206}), .b ({1'b0, 1'b1}), .a ({signal_1833, signal_1458}), .clk (clk), .r (Fresh[61]), .c ({signal_2050, signal_1517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1317 ( .s ({signal_3200, signal_3198}), .b ({1'b0, 1'b1}), .a ({signal_1831, signal_1457}), .clk (clk), .r (Fresh[62]), .c ({signal_2051, signal_1518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1318 ( .s ({signal_3220, signal_3218}), .b ({signal_1847, signal_1466}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[63]), .c ({signal_2053, signal_1519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1319 ( .s ({signal_3180, signal_3178}), .b ({signal_1857, signal_1473}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[64]), .c ({signal_2054, signal_1520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1320 ( .s ({signal_3192, signal_3190}), .b ({1'b0, 1'b0}), .a ({signal_1851, signal_1469}), .clk (clk), .r (Fresh[65]), .c ({signal_2055, signal_1521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1321 ( .s ({signal_3224, signal_3222}), .b ({signal_1866, signal_1480}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[66]), .c ({signal_2057, signal_1522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1322 ( .s ({signal_3196, signal_3194}), .b ({1'b0, 1'b1}), .a ({signal_1845, signal_1465}), .clk (clk), .r (Fresh[67]), .c ({signal_2058, signal_1523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1323 ( .s ({signal_3228, signal_3226}), .b ({1'b0, 1'b0}), .a ({signal_1858, signal_1474}), .clk (clk), .r (Fresh[68]), .c ({signal_2060, signal_1524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1324 ( .s ({signal_3168, signal_3166}), .b ({1'b0, 1'b1}), .a ({signal_1844, signal_1464}), .clk (clk), .r (Fresh[69]), .c ({signal_2061, signal_1525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1325 ( .s ({signal_3200, signal_3198}), .b ({signal_1831, signal_1457}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[70]), .c ({signal_2062, signal_1526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1326 ( .s ({signal_3180, signal_3178}), .b ({1'b0, 1'b1}), .a ({signal_1865, signal_1479}), .clk (clk), .r (Fresh[71]), .c ({signal_2063, signal_1527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1327 ( .s ({signal_3232, signal_3230}), .b ({signal_1831, signal_1457}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[72]), .c ({signal_2065, signal_1528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1328 ( .s ({signal_3204, signal_3202}), .b ({signal_1861, signal_1476}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[73]), .c ({signal_2066, signal_1529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1329 ( .s ({signal_3236, signal_3234}), .b ({signal_1835, signal_1459}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[74]), .c ({signal_2068, signal_1530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1330 ( .s ({signal_3228, signal_3226}), .b ({signal_1858, signal_1474}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[75]), .c ({signal_2069, signal_1531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1331 ( .s ({signal_3240, signal_3238}), .b ({signal_1844, signal_1464}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[76]), .c ({signal_2071, signal_1532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1332 ( .s ({signal_3244, signal_3242}), .b ({signal_1829, signal_1456}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[77]), .c ({signal_2073, signal_1533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1333 ( .s ({signal_3188, signal_3186}), .b ({1'b0, 1'b1}), .a ({signal_1863, signal_1477}), .clk (clk), .r (Fresh[78]), .c ({signal_2074, signal_1534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1334 ( .s ({signal_3248, signal_3246}), .b ({signal_1863, signal_1477}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[79]), .c ({signal_2076, signal_1535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1335 ( .s ({signal_3192, signal_3190}), .b ({signal_1851, signal_1469}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[80]), .c ({signal_2077, signal_1536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1336 ( .s ({signal_3228, signal_3226}), .b ({signal_1855, signal_1472}), .a ({signal_1858, signal_1474}), .clk (clk), .r (Fresh[81]), .c ({signal_2078, signal_1537}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1337 ( .s ({signal_3192, signal_3190}), .b ({1'b0, 1'b1}), .a ({signal_1851, signal_1469}), .clk (clk), .r (Fresh[82]), .c ({signal_2079, signal_1538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1338 ( .s ({signal_3228, signal_3226}), .b ({1'b0, 1'b1}), .a ({signal_1858, signal_1474}), .clk (clk), .r (Fresh[83]), .c ({signal_2080, signal_1539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1339 ( .s ({signal_3188, signal_3186}), .b ({signal_1863, signal_1477}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[84]), .c ({signal_2081, signal_1540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1340 ( .s ({signal_3228, signal_3226}), .b ({signal_1855, signal_1472}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[85]), .c ({signal_2082, signal_1541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1341 ( .s ({signal_3208, signal_3206}), .b ({1'b0, 1'b0}), .a ({signal_1833, signal_1458}), .clk (clk), .r (Fresh[86]), .c ({signal_2083, signal_1542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1342 ( .s ({signal_3176, signal_3174}), .b ({signal_1837, signal_1460}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[87]), .c ({signal_2084, signal_1543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1343 ( .s ({signal_3200, signal_3198}), .b ({signal_1853, signal_1471}), .a ({signal_1831, signal_1457}), .clk (clk), .r (Fresh[88]), .c ({signal_2085, signal_1544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1344 ( .s ({signal_3204, signal_3202}), .b ({1'b0, 1'b1}), .a ({signal_1866, signal_1480}), .clk (clk), .r (Fresh[89]), .c ({signal_2086, signal_1545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1345 ( .s ({signal_3204, signal_3202}), .b ({signal_1861, signal_1476}), .a ({signal_1866, signal_1480}), .clk (clk), .r (Fresh[90]), .c ({signal_2087, signal_1546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1346 ( .s ({signal_3196, signal_3194}), .b ({signal_1840, signal_1462}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[91]), .c ({signal_2088, signal_1547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1347 ( .s ({signal_3168, signal_3166}), .b ({signal_1844, signal_1464}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[92]), .c ({signal_2089, signal_1548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1348 ( .s ({signal_3192, signal_3190}), .b ({signal_1859, signal_1475}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[93]), .c ({signal_2090, signal_1549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1349 ( .s ({signal_3200, signal_3198}), .b ({1'b0, 1'b0}), .a ({signal_1831, signal_1457}), .clk (clk), .r (Fresh[94]), .c ({signal_2091, signal_1550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1350 ( .s ({signal_3176, signal_3174}), .b ({1'b0, 1'b1}), .a ({signal_1838, signal_1461}), .clk (clk), .r (Fresh[95]), .c ({signal_2092, signal_1551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1351 ( .s ({signal_3188, signal_3186}), .b ({signal_1867, signal_1481}), .a ({signal_1863, signal_1477}), .clk (clk), .r (Fresh[96]), .c ({signal_2093, signal_1552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1352 ( .s ({signal_3252, signal_3250}), .b ({signal_1865, signal_1479}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[97]), .c ({signal_2095, signal_1553}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1353 ( .s ({signal_3208, signal_3206}), .b ({signal_1852, signal_1470}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[98]), .c ({signal_2096, signal_1554}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1354 ( .s ({signal_3188, signal_3186}), .b ({signal_1867, signal_1481}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[99]), .c ({signal_2097, signal_1555}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1355 ( .s ({signal_3256, signal_3254}), .b ({1'b0, 1'b1}), .a ({signal_1835, signal_1459}), .clk (clk), .r (Fresh[100]), .c ({signal_2099, signal_1556}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1356 ( .s ({signal_3256, signal_3254}), .b ({signal_1864, signal_1478}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[101]), .c ({signal_2100, signal_1557}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1357 ( .s ({signal_3256, signal_3254}), .b ({signal_1835, signal_1459}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[102]), .c ({signal_2101, signal_1558}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1358 ( .s ({signal_3172, signal_3170}), .b ({signal_1848, signal_1467}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[103]), .c ({signal_2102, signal_1559}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1359 ( .s ({signal_3172, signal_3170}), .b ({1'b0, 1'b1}), .a ({signal_1848, signal_1467}), .clk (clk), .r (Fresh[104]), .c ({signal_2103, signal_1560}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1360 ( .s ({signal_3256, signal_3254}), .b ({1'b0, 1'b0}), .a ({signal_1835, signal_1459}), .clk (clk), .r (Fresh[105]), .c ({signal_2104, signal_1561}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1361 ( .s ({signal_3256, signal_3254}), .b ({signal_1864, signal_1478}), .a ({signal_1835, signal_1459}), .clk (clk), .r (Fresh[106]), .c ({signal_2105, signal_1562}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .s ({signal_3260, signal_3258}), .b ({signal_1871, signal_1483}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[107]), .c ({signal_2107, signal_1563}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .s ({signal_3264, signal_3262}), .b ({1'b0, 1'b1}), .a ({signal_1872, signal_1484}), .clk (clk), .r (Fresh[108]), .c ({signal_2108, signal_1564}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .s ({signal_3264, signal_3262}), .b ({signal_1869, signal_1482}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[109]), .c ({signal_2109, signal_1565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .s ({signal_3264, signal_3262}), .b ({1'b0, 1'b1}), .a ({signal_1869, signal_1482}), .clk (clk), .r (Fresh[110]), .c ({signal_2110, signal_1566}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .s ({signal_3264, signal_3262}), .b ({signal_1869, signal_1482}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[111]), .c ({signal_2111, signal_1567}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .s ({signal_3264, signal_3262}), .b ({signal_1869, signal_1482}), .a ({signal_1872, signal_1484}), .clk (clk), .r (Fresh[112]), .c ({signal_2112, signal_1568}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1368 ( .s ({signal_3268, signal_3266}), .b ({signal_1876, signal_1486}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[113]), .c ({signal_2114, signal_1569}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1369 ( .s ({signal_3272, signal_3270}), .b ({1'b0, 1'b1}), .a ({signal_1877, signal_1487}), .clk (clk), .r (Fresh[114]), .c ({signal_2115, signal_1570}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1370 ( .s ({signal_3272, signal_3270}), .b ({signal_1874, signal_1485}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[115]), .c ({signal_2116, signal_1571}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1371 ( .s ({signal_3272, signal_3270}), .b ({1'b0, 1'b1}), .a ({signal_1874, signal_1485}), .clk (clk), .r (Fresh[116]), .c ({signal_2117, signal_1572}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1372 ( .s ({signal_3272, signal_3270}), .b ({signal_1874, signal_1485}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[117]), .c ({signal_2118, signal_1573}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1373 ( .s ({signal_3272, signal_3270}), .b ({signal_1874, signal_1485}), .a ({signal_1877, signal_1487}), .clk (clk), .r (Fresh[118]), .c ({signal_2119, signal_1574}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1374 ( .s ({signal_3172, signal_3170}), .b ({signal_1848, signal_1467}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[119]), .c ({signal_2120, signal_1575}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1375 ( .s ({signal_3276, signal_3274}), .b ({signal_1881, signal_1489}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[120]), .c ({signal_2122, signal_1576}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1376 ( .s ({signal_3280, signal_3278}), .b ({1'b0, 1'b1}), .a ({signal_1882, signal_1490}), .clk (clk), .r (Fresh[121]), .c ({signal_2123, signal_1577}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1377 ( .s ({signal_3280, signal_3278}), .b ({signal_1879, signal_1488}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[122]), .c ({signal_2124, signal_1578}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1378 ( .s ({signal_3280, signal_3278}), .b ({1'b0, 1'b1}), .a ({signal_1879, signal_1488}), .clk (clk), .r (Fresh[123]), .c ({signal_2125, signal_1579}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1379 ( .s ({signal_3280, signal_3278}), .b ({signal_1879, signal_1488}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[124]), .c ({signal_2126, signal_1580}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1380 ( .s ({signal_3280, signal_3278}), .b ({signal_1879, signal_1488}), .a ({signal_1882, signal_1490}), .clk (clk), .r (Fresh[125]), .c ({signal_2127, signal_1581}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1381 ( .s ({signal_3284, signal_3282}), .b ({signal_1886, signal_1492}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[126]), .c ({signal_2129, signal_1582}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1382 ( .s ({signal_3288, signal_3286}), .b ({1'b0, 1'b1}), .a ({signal_1887, signal_1493}), .clk (clk), .r (Fresh[127]), .c ({signal_2130, signal_1583}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1383 ( .s ({signal_3288, signal_3286}), .b ({signal_1884, signal_1491}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[128]), .c ({signal_2131, signal_1584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .s ({signal_3288, signal_3286}), .b ({1'b0, 1'b1}), .a ({signal_1884, signal_1491}), .clk (clk), .r (Fresh[129]), .c ({signal_2132, signal_1585}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .s ({signal_3288, signal_3286}), .b ({signal_1884, signal_1491}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[130]), .c ({signal_2133, signal_1586}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .s ({signal_3288, signal_3286}), .b ({signal_1884, signal_1491}), .a ({signal_1887, signal_1493}), .clk (clk), .r (Fresh[131]), .c ({signal_2134, signal_1587}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .s ({signal_3292, signal_3290}), .b ({signal_1889, signal_1494}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[132]), .c ({signal_2136, signal_1588}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .s ({signal_3196, signal_3194}), .b ({signal_1840, signal_1462}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[133]), .c ({signal_2137, signal_1589}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .s ({signal_3172, signal_3170}), .b ({signal_1848, signal_1467}), .a ({signal_1842, signal_1463}), .clk (clk), .r (Fresh[134]), .c ({signal_2138, signal_1590}) ) ;
    buf_clk cell_1553 ( .C (clk), .D (signal_3095), .Q (signal_3096) ) ;
    buf_clk cell_1753 ( .C (clk), .D (signal_3295), .Q (signal_3296) ) ;
    buf_clk cell_1759 ( .C (clk), .D (signal_3301), .Q (signal_3302) ) ;
    buf_clk cell_1765 ( .C (clk), .D (signal_3307), .Q (signal_3308) ) ;
    buf_clk cell_1771 ( .C (clk), .D (signal_3313), .Q (signal_3314) ) ;
    buf_clk cell_1777 ( .C (clk), .D (signal_3319), .Q (signal_3320) ) ;
    buf_clk cell_1783 ( .C (clk), .D (signal_3325), .Q (signal_3326) ) ;
    buf_clk cell_1789 ( .C (clk), .D (signal_3331), .Q (signal_3332) ) ;
    buf_clk cell_1795 ( .C (clk), .D (signal_3337), .Q (signal_3338) ) ;
    buf_clk cell_1801 ( .C (clk), .D (signal_3343), .Q (signal_3344) ) ;
    buf_clk cell_1807 ( .C (clk), .D (signal_3349), .Q (signal_3350) ) ;
    buf_clk cell_1813 ( .C (clk), .D (signal_3355), .Q (signal_3356) ) ;
    buf_clk cell_1819 ( .C (clk), .D (signal_3361), .Q (signal_3362) ) ;
    buf_clk cell_1825 ( .C (clk), .D (signal_3367), .Q (signal_3368) ) ;
    buf_clk cell_1831 ( .C (clk), .D (signal_3373), .Q (signal_3374) ) ;
    buf_clk cell_1837 ( .C (clk), .D (signal_3379), .Q (signal_3380) ) ;
    buf_clk cell_1843 ( .C (clk), .D (signal_3385), .Q (signal_3386) ) ;
    buf_clk cell_1849 ( .C (clk), .D (signal_3391), .Q (signal_3392) ) ;
    buf_clk cell_1855 ( .C (clk), .D (signal_3397), .Q (signal_3398) ) ;
    buf_clk cell_1861 ( .C (clk), .D (signal_3403), .Q (signal_3404) ) ;
    buf_clk cell_1867 ( .C (clk), .D (signal_3409), .Q (signal_3410) ) ;
    buf_clk cell_1873 ( .C (clk), .D (signal_3415), .Q (signal_3416) ) ;
    buf_clk cell_1879 ( .C (clk), .D (signal_3421), .Q (signal_3422) ) ;
    buf_clk cell_1885 ( .C (clk), .D (signal_3427), .Q (signal_3428) ) ;
    buf_clk cell_1891 ( .C (clk), .D (signal_3433), .Q (signal_3434) ) ;
    buf_clk cell_1897 ( .C (clk), .D (signal_3439), .Q (signal_3440) ) ;
    buf_clk cell_1903 ( .C (clk), .D (signal_3445), .Q (signal_3446) ) ;
    buf_clk cell_1909 ( .C (clk), .D (signal_3451), .Q (signal_3452) ) ;
    buf_clk cell_1915 ( .C (clk), .D (signal_3457), .Q (signal_3458) ) ;
    buf_clk cell_1921 ( .C (clk), .D (signal_3463), .Q (signal_3464) ) ;
    buf_clk cell_1927 ( .C (clk), .D (signal_3469), .Q (signal_3470) ) ;
    buf_clk cell_1933 ( .C (clk), .D (signal_3475), .Q (signal_3476) ) ;
    buf_clk cell_1939 ( .C (clk), .D (signal_3481), .Q (signal_3482) ) ;
    buf_clk cell_1945 ( .C (clk), .D (signal_3487), .Q (signal_3488) ) ;
    buf_clk cell_1951 ( .C (clk), .D (signal_3493), .Q (signal_3494) ) ;
    buf_clk cell_1957 ( .C (clk), .D (signal_3499), .Q (signal_3500) ) ;
    buf_clk cell_1963 ( .C (clk), .D (signal_3505), .Q (signal_3506) ) ;
    buf_clk cell_1969 ( .C (clk), .D (signal_3511), .Q (signal_3512) ) ;
    buf_clk cell_1975 ( .C (clk), .D (signal_3517), .Q (signal_3518) ) ;
    buf_clk cell_1981 ( .C (clk), .D (signal_3523), .Q (signal_3524) ) ;
    buf_clk cell_1987 ( .C (clk), .D (signal_3529), .Q (signal_3530) ) ;
    buf_clk cell_1993 ( .C (clk), .D (signal_3535), .Q (signal_3536) ) ;
    buf_clk cell_1999 ( .C (clk), .D (signal_3541), .Q (signal_3542) ) ;
    buf_clk cell_2005 ( .C (clk), .D (signal_3547), .Q (signal_3548) ) ;
    buf_clk cell_2011 ( .C (clk), .D (signal_3553), .Q (signal_3554) ) ;
    buf_clk cell_2017 ( .C (clk), .D (signal_3559), .Q (signal_3560) ) ;
    buf_clk cell_2023 ( .C (clk), .D (signal_3565), .Q (signal_3566) ) ;
    buf_clk cell_2029 ( .C (clk), .D (signal_3571), .Q (signal_3572) ) ;
    buf_clk cell_2035 ( .C (clk), .D (signal_3577), .Q (signal_3578) ) ;
    buf_clk cell_2041 ( .C (clk), .D (signal_3583), .Q (signal_3584) ) ;
    buf_clk cell_2047 ( .C (clk), .D (signal_3589), .Q (signal_3590) ) ;
    buf_clk cell_2053 ( .C (clk), .D (signal_3595), .Q (signal_3596) ) ;
    buf_clk cell_2059 ( .C (clk), .D (signal_3601), .Q (signal_3602) ) ;
    buf_clk cell_2065 ( .C (clk), .D (signal_3607), .Q (signal_3608) ) ;
    buf_clk cell_2071 ( .C (clk), .D (signal_3613), .Q (signal_3614) ) ;
    buf_clk cell_2077 ( .C (clk), .D (signal_3619), .Q (signal_3620) ) ;
    buf_clk cell_2083 ( .C (clk), .D (signal_3625), .Q (signal_3626) ) ;
    buf_clk cell_2089 ( .C (clk), .D (signal_3631), .Q (signal_3632) ) ;
    buf_clk cell_2095 ( .C (clk), .D (signal_3637), .Q (signal_3638) ) ;
    buf_clk cell_2101 ( .C (clk), .D (signal_3643), .Q (signal_3644) ) ;
    buf_clk cell_2107 ( .C (clk), .D (signal_3649), .Q (signal_3650) ) ;
    buf_clk cell_2113 ( .C (clk), .D (signal_3655), .Q (signal_3656) ) ;
    buf_clk cell_2119 ( .C (clk), .D (signal_3661), .Q (signal_3662) ) ;
    buf_clk cell_2125 ( .C (clk), .D (signal_3667), .Q (signal_3668) ) ;
    buf_clk cell_2131 ( .C (clk), .D (signal_3673), .Q (signal_3674) ) ;
    buf_clk cell_2137 ( .C (clk), .D (signal_3679), .Q (signal_3680) ) ;
    buf_clk cell_2143 ( .C (clk), .D (signal_3685), .Q (signal_3686) ) ;
    buf_clk cell_2149 ( .C (clk), .D (signal_3691), .Q (signal_3692) ) ;
    buf_clk cell_2155 ( .C (clk), .D (signal_3697), .Q (signal_3698) ) ;
    buf_clk cell_2161 ( .C (clk), .D (signal_3703), .Q (signal_3704) ) ;
    buf_clk cell_2167 ( .C (clk), .D (signal_3709), .Q (signal_3710) ) ;
    buf_clk cell_2173 ( .C (clk), .D (signal_3715), .Q (signal_3716) ) ;
    buf_clk cell_2179 ( .C (clk), .D (signal_3721), .Q (signal_3722) ) ;
    buf_clk cell_2185 ( .C (clk), .D (signal_3727), .Q (signal_3728) ) ;
    buf_clk cell_2191 ( .C (clk), .D (signal_3733), .Q (signal_3734) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_3739), .Q (signal_3740) ) ;
    buf_clk cell_2203 ( .C (clk), .D (signal_3745), .Q (signal_3746) ) ;
    buf_clk cell_2209 ( .C (clk), .D (signal_3751), .Q (signal_3752) ) ;
    buf_clk cell_2215 ( .C (clk), .D (signal_3757), .Q (signal_3758) ) ;
    buf_clk cell_2221 ( .C (clk), .D (signal_3763), .Q (signal_3764) ) ;
    buf_clk cell_2227 ( .C (clk), .D (signal_3769), .Q (signal_3770) ) ;
    buf_clk cell_2233 ( .C (clk), .D (signal_3775), .Q (signal_3776) ) ;
    buf_clk cell_2239 ( .C (clk), .D (signal_3781), .Q (signal_3782) ) ;
    buf_clk cell_2245 ( .C (clk), .D (signal_3787), .Q (signal_3788) ) ;
    buf_clk cell_2251 ( .C (clk), .D (signal_3793), .Q (signal_3794) ) ;
    buf_clk cell_2257 ( .C (clk), .D (signal_3799), .Q (signal_3800) ) ;
    buf_clk cell_2263 ( .C (clk), .D (signal_3805), .Q (signal_3806) ) ;
    buf_clk cell_2269 ( .C (clk), .D (signal_3811), .Q (signal_3812) ) ;
    buf_clk cell_2275 ( .C (clk), .D (signal_3817), .Q (signal_3818) ) ;
    buf_clk cell_2281 ( .C (clk), .D (signal_3823), .Q (signal_3824) ) ;
    buf_clk cell_2287 ( .C (clk), .D (signal_3829), .Q (signal_3830) ) ;
    buf_clk cell_2293 ( .C (clk), .D (signal_3835), .Q (signal_3836) ) ;
    buf_clk cell_2299 ( .C (clk), .D (signal_3841), .Q (signal_3842) ) ;
    buf_clk cell_2305 ( .C (clk), .D (signal_3847), .Q (signal_3848) ) ;
    buf_clk cell_2311 ( .C (clk), .D (signal_3853), .Q (signal_3854) ) ;
    buf_clk cell_2317 ( .C (clk), .D (signal_3859), .Q (signal_3860) ) ;
    buf_clk cell_2323 ( .C (clk), .D (signal_3865), .Q (signal_3866) ) ;
    buf_clk cell_2329 ( .C (clk), .D (signal_3871), .Q (signal_3872) ) ;
    buf_clk cell_2335 ( .C (clk), .D (signal_3877), .Q (signal_3878) ) ;
    buf_clk cell_2341 ( .C (clk), .D (signal_3883), .Q (signal_3884) ) ;
    buf_clk cell_2347 ( .C (clk), .D (signal_3889), .Q (signal_3890) ) ;
    buf_clk cell_2353 ( .C (clk), .D (signal_3895), .Q (signal_3896) ) ;
    buf_clk cell_2359 ( .C (clk), .D (signal_3901), .Q (signal_3902) ) ;
    buf_clk cell_2365 ( .C (clk), .D (signal_3907), .Q (signal_3908) ) ;
    buf_clk cell_2371 ( .C (clk), .D (signal_3913), .Q (signal_3914) ) ;
    buf_clk cell_2377 ( .C (clk), .D (signal_3919), .Q (signal_3920) ) ;
    buf_clk cell_2383 ( .C (clk), .D (signal_3925), .Q (signal_3926) ) ;
    buf_clk cell_2389 ( .C (clk), .D (signal_3931), .Q (signal_3932) ) ;
    buf_clk cell_2395 ( .C (clk), .D (signal_3937), .Q (signal_3938) ) ;
    buf_clk cell_2401 ( .C (clk), .D (signal_3943), .Q (signal_3944) ) ;
    buf_clk cell_2407 ( .C (clk), .D (signal_3949), .Q (signal_3950) ) ;
    buf_clk cell_2413 ( .C (clk), .D (signal_3955), .Q (signal_3956) ) ;
    buf_clk cell_2419 ( .C (clk), .D (signal_3961), .Q (signal_3962) ) ;
    buf_clk cell_2425 ( .C (clk), .D (signal_3967), .Q (signal_3968) ) ;
    buf_clk cell_2431 ( .C (clk), .D (signal_3973), .Q (signal_3974) ) ;
    buf_clk cell_2437 ( .C (clk), .D (signal_3979), .Q (signal_3980) ) ;
    buf_clk cell_2443 ( .C (clk), .D (signal_3985), .Q (signal_3986) ) ;
    buf_clk cell_2449 ( .C (clk), .D (signal_3991), .Q (signal_3992) ) ;
    buf_clk cell_2455 ( .C (clk), .D (signal_3997), .Q (signal_3998) ) ;
    buf_clk cell_2461 ( .C (clk), .D (signal_4003), .Q (signal_4004) ) ;
    buf_clk cell_2467 ( .C (clk), .D (signal_4009), .Q (signal_4010) ) ;
    buf_clk cell_2473 ( .C (clk), .D (signal_4015), .Q (signal_4016) ) ;
    buf_clk cell_2479 ( .C (clk), .D (signal_4021), .Q (signal_4022) ) ;
    buf_clk cell_2485 ( .C (clk), .D (signal_4027), .Q (signal_4028) ) ;
    buf_clk cell_2491 ( .C (clk), .D (signal_4033), .Q (signal_4034) ) ;
    buf_clk cell_2497 ( .C (clk), .D (signal_4039), .Q (signal_4040) ) ;
    buf_clk cell_2503 ( .C (clk), .D (signal_4045), .Q (signal_4046) ) ;
    buf_clk cell_2509 ( .C (clk), .D (signal_4051), .Q (signal_4052) ) ;
    buf_clk cell_2515 ( .C (clk), .D (signal_4057), .Q (signal_4058) ) ;
    buf_clk cell_2521 ( .C (clk), .D (signal_4063), .Q (signal_4064) ) ;
    buf_clk cell_2527 ( .C (clk), .D (signal_4069), .Q (signal_4070) ) ;
    buf_clk cell_2533 ( .C (clk), .D (signal_4075), .Q (signal_4076) ) ;
    buf_clk cell_2539 ( .C (clk), .D (signal_4081), .Q (signal_4082) ) ;
    buf_clk cell_2545 ( .C (clk), .D (signal_4087), .Q (signal_4088) ) ;
    buf_clk cell_2551 ( .C (clk), .D (signal_4093), .Q (signal_4094) ) ;
    buf_clk cell_2557 ( .C (clk), .D (signal_4099), .Q (signal_4100) ) ;
    buf_clk cell_2563 ( .C (clk), .D (signal_4105), .Q (signal_4106) ) ;
    buf_clk cell_2569 ( .C (clk), .D (signal_4111), .Q (signal_4112) ) ;
    buf_clk cell_2575 ( .C (clk), .D (signal_4117), .Q (signal_4118) ) ;
    buf_clk cell_2581 ( .C (clk), .D (signal_4123), .Q (signal_4124) ) ;
    buf_clk cell_2587 ( .C (clk), .D (signal_4129), .Q (signal_4130) ) ;
    buf_clk cell_2593 ( .C (clk), .D (signal_4135), .Q (signal_4136) ) ;
    buf_clk cell_2599 ( .C (clk), .D (signal_4141), .Q (signal_4142) ) ;
    buf_clk cell_2605 ( .C (clk), .D (signal_4147), .Q (signal_4148) ) ;
    buf_clk cell_2611 ( .C (clk), .D (signal_4153), .Q (signal_4154) ) ;
    buf_clk cell_2617 ( .C (clk), .D (signal_4159), .Q (signal_4160) ) ;
    buf_clk cell_2623 ( .C (clk), .D (signal_4165), .Q (signal_4166) ) ;
    buf_clk cell_2629 ( .C (clk), .D (signal_4171), .Q (signal_4172) ) ;
    buf_clk cell_2635 ( .C (clk), .D (signal_4177), .Q (signal_4178) ) ;
    buf_clk cell_2641 ( .C (clk), .D (signal_4183), .Q (signal_4184) ) ;
    buf_clk cell_2647 ( .C (clk), .D (signal_4189), .Q (signal_4190) ) ;
    buf_clk cell_2653 ( .C (clk), .D (signal_4195), .Q (signal_4196) ) ;
    buf_clk cell_2659 ( .C (clk), .D (signal_4201), .Q (signal_4202) ) ;
    buf_clk cell_2665 ( .C (clk), .D (signal_4207), .Q (signal_4208) ) ;
    buf_clk cell_2671 ( .C (clk), .D (signal_4213), .Q (signal_4214) ) ;
    buf_clk cell_2677 ( .C (clk), .D (signal_4219), .Q (signal_4220) ) ;
    buf_clk cell_2683 ( .C (clk), .D (signal_4225), .Q (signal_4226) ) ;
    buf_clk cell_2689 ( .C (clk), .D (signal_4231), .Q (signal_4232) ) ;
    buf_clk cell_2695 ( .C (clk), .D (signal_4237), .Q (signal_4238) ) ;
    buf_clk cell_2701 ( .C (clk), .D (signal_4243), .Q (signal_4244) ) ;
    buf_clk cell_2707 ( .C (clk), .D (signal_4249), .Q (signal_4250) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_4255), .Q (signal_4256) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_4261), .Q (signal_4262) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_4267), .Q (signal_4268) ) ;
    buf_clk cell_2731 ( .C (clk), .D (signal_4273), .Q (signal_4274) ) ;
    buf_clk cell_2737 ( .C (clk), .D (signal_4279), .Q (signal_4280) ) ;
    buf_clk cell_2743 ( .C (clk), .D (signal_4285), .Q (signal_4286) ) ;
    buf_clk cell_2749 ( .C (clk), .D (signal_4291), .Q (signal_4292) ) ;
    buf_clk cell_2755 ( .C (clk), .D (signal_4297), .Q (signal_4298) ) ;
    buf_clk cell_2761 ( .C (clk), .D (signal_4303), .Q (signal_4304) ) ;
    buf_clk cell_2767 ( .C (clk), .D (signal_4309), .Q (signal_4310) ) ;
    buf_clk cell_2773 ( .C (clk), .D (signal_4315), .Q (signal_4316) ) ;
    buf_clk cell_2779 ( .C (clk), .D (signal_4321), .Q (signal_4322) ) ;
    buf_clk cell_2785 ( .C (clk), .D (signal_4327), .Q (signal_4328) ) ;
    buf_clk cell_2791 ( .C (clk), .D (signal_4333), .Q (signal_4334) ) ;
    buf_clk cell_2797 ( .C (clk), .D (signal_4339), .Q (signal_4340) ) ;
    buf_clk cell_2803 ( .C (clk), .D (signal_4345), .Q (signal_4346) ) ;
    buf_clk cell_2809 ( .C (clk), .D (signal_4351), .Q (signal_4352) ) ;
    buf_clk cell_2815 ( .C (clk), .D (signal_4357), .Q (signal_4358) ) ;
    buf_clk cell_2821 ( .C (clk), .D (signal_4363), .Q (signal_4364) ) ;
    buf_clk cell_2827 ( .C (clk), .D (signal_4369), .Q (signal_4370) ) ;
    buf_clk cell_2833 ( .C (clk), .D (signal_4375), .Q (signal_4376) ) ;
    buf_clk cell_2839 ( .C (clk), .D (signal_4381), .Q (signal_4382) ) ;
    buf_clk cell_2845 ( .C (clk), .D (signal_4387), .Q (signal_4388) ) ;
    buf_clk cell_2851 ( .C (clk), .D (signal_4393), .Q (signal_4394) ) ;
    buf_clk cell_2857 ( .C (clk), .D (signal_4399), .Q (signal_4400) ) ;
    buf_clk cell_2863 ( .C (clk), .D (signal_4405), .Q (signal_4406) ) ;
    buf_clk cell_2869 ( .C (clk), .D (signal_4411), .Q (signal_4412) ) ;
    buf_clk cell_2875 ( .C (clk), .D (signal_4417), .Q (signal_4418) ) ;
    buf_clk cell_2881 ( .C (clk), .D (signal_4423), .Q (signal_4424) ) ;
    buf_clk cell_2887 ( .C (clk), .D (signal_4429), .Q (signal_4430) ) ;
    buf_clk cell_2893 ( .C (clk), .D (signal_4435), .Q (signal_4436) ) ;
    buf_clk cell_2899 ( .C (clk), .D (signal_4441), .Q (signal_4442) ) ;
    buf_clk cell_2905 ( .C (clk), .D (signal_4447), .Q (signal_4448) ) ;
    buf_clk cell_2911 ( .C (clk), .D (signal_4453), .Q (signal_4454) ) ;
    buf_clk cell_2915 ( .C (clk), .D (signal_4457), .Q (signal_4458) ) ;
    buf_clk cell_2917 ( .C (clk), .D (signal_4459), .Q (signal_4460) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_4463), .Q (signal_4464) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_4467), .Q (signal_4468) ) ;
    buf_clk cell_2927 ( .C (clk), .D (signal_4469), .Q (signal_4470) ) ;
    buf_clk cell_2929 ( .C (clk), .D (signal_4471), .Q (signal_4472) ) ;
    buf_clk cell_2931 ( .C (clk), .D (signal_4473), .Q (signal_4474) ) ;
    buf_clk cell_2933 ( .C (clk), .D (signal_4475), .Q (signal_4476) ) ;
    buf_clk cell_2935 ( .C (clk), .D (signal_4477), .Q (signal_4478) ) ;
    buf_clk cell_2937 ( .C (clk), .D (signal_4479), .Q (signal_4480) ) ;
    buf_clk cell_2939 ( .C (clk), .D (signal_4481), .Q (signal_4482) ) ;
    buf_clk cell_2941 ( .C (clk), .D (signal_4483), .Q (signal_4484) ) ;
    buf_clk cell_2943 ( .C (clk), .D (signal_4485), .Q (signal_4486) ) ;
    buf_clk cell_2945 ( .C (clk), .D (signal_4487), .Q (signal_4488) ) ;
    buf_clk cell_2947 ( .C (clk), .D (signal_4489), .Q (signal_4490) ) ;
    buf_clk cell_2949 ( .C (clk), .D (signal_4491), .Q (signal_4492) ) ;
    buf_clk cell_2951 ( .C (clk), .D (signal_4493), .Q (signal_4494) ) ;
    buf_clk cell_2953 ( .C (clk), .D (signal_4495), .Q (signal_4496) ) ;
    buf_clk cell_2957 ( .C (clk), .D (signal_4499), .Q (signal_4500) ) ;
    buf_clk cell_2961 ( .C (clk), .D (signal_4503), .Q (signal_4504) ) ;
    buf_clk cell_2965 ( .C (clk), .D (signal_4507), .Q (signal_4508) ) ;
    buf_clk cell_2969 ( .C (clk), .D (signal_4511), .Q (signal_4512) ) ;
    buf_clk cell_2971 ( .C (clk), .D (signal_4513), .Q (signal_4514) ) ;
    buf_clk cell_2973 ( .C (clk), .D (signal_4515), .Q (signal_4516) ) ;
    buf_clk cell_2977 ( .C (clk), .D (signal_4519), .Q (signal_4520) ) ;
    buf_clk cell_2981 ( .C (clk), .D (signal_4523), .Q (signal_4524) ) ;
    buf_clk cell_2985 ( .C (clk), .D (signal_4527), .Q (signal_4528) ) ;
    buf_clk cell_2989 ( .C (clk), .D (signal_4531), .Q (signal_4532) ) ;
    buf_clk cell_2993 ( .C (clk), .D (signal_4535), .Q (signal_4536) ) ;
    buf_clk cell_2997 ( .C (clk), .D (signal_4539), .Q (signal_4540) ) ;
    buf_clk cell_2999 ( .C (clk), .D (signal_4541), .Q (signal_4542) ) ;
    buf_clk cell_3001 ( .C (clk), .D (signal_4543), .Q (signal_4544) ) ;
    buf_clk cell_3005 ( .C (clk), .D (signal_4547), .Q (signal_4548) ) ;
    buf_clk cell_3009 ( .C (clk), .D (signal_4551), .Q (signal_4552) ) ;
    buf_clk cell_3013 ( .C (clk), .D (signal_4555), .Q (signal_4556) ) ;
    buf_clk cell_3017 ( .C (clk), .D (signal_4559), .Q (signal_4560) ) ;
    buf_clk cell_3021 ( .C (clk), .D (signal_4563), .Q (signal_4564) ) ;
    buf_clk cell_3025 ( .C (clk), .D (signal_4567), .Q (signal_4568) ) ;
    buf_clk cell_3029 ( .C (clk), .D (signal_4571), .Q (signal_4572) ) ;
    buf_clk cell_3033 ( .C (clk), .D (signal_4575), .Q (signal_4576) ) ;
    buf_clk cell_3037 ( .C (clk), .D (signal_4579), .Q (signal_4580) ) ;
    buf_clk cell_3041 ( .C (clk), .D (signal_4583), .Q (signal_4584) ) ;
    buf_clk cell_3043 ( .C (clk), .D (signal_4585), .Q (signal_4586) ) ;
    buf_clk cell_3045 ( .C (clk), .D (signal_4587), .Q (signal_4588) ) ;
    buf_clk cell_3047 ( .C (clk), .D (signal_4589), .Q (signal_4590) ) ;
    buf_clk cell_3049 ( .C (clk), .D (signal_4591), .Q (signal_4592) ) ;
    buf_clk cell_3053 ( .C (clk), .D (signal_4595), .Q (signal_4596) ) ;
    buf_clk cell_3057 ( .C (clk), .D (signal_4599), .Q (signal_4600) ) ;
    buf_clk cell_3059 ( .C (clk), .D (signal_4601), .Q (signal_4602) ) ;
    buf_clk cell_3061 ( .C (clk), .D (signal_4603), .Q (signal_4604) ) ;
    buf_clk cell_3065 ( .C (clk), .D (signal_4607), .Q (signal_4608) ) ;
    buf_clk cell_3069 ( .C (clk), .D (signal_4611), .Q (signal_4612) ) ;
    buf_clk cell_3071 ( .C (clk), .D (signal_4613), .Q (signal_4614) ) ;
    buf_clk cell_3073 ( .C (clk), .D (signal_4615), .Q (signal_4616) ) ;
    buf_clk cell_3077 ( .C (clk), .D (signal_4619), .Q (signal_4620) ) ;
    buf_clk cell_3081 ( .C (clk), .D (signal_4623), .Q (signal_4624) ) ;
    buf_clk cell_3083 ( .C (clk), .D (signal_4625), .Q (signal_4626) ) ;
    buf_clk cell_3085 ( .C (clk), .D (signal_4627), .Q (signal_4628) ) ;
    buf_clk cell_3089 ( .C (clk), .D (signal_4631), .Q (signal_4632) ) ;
    buf_clk cell_3093 ( .C (clk), .D (signal_4635), .Q (signal_4636) ) ;
    buf_clk cell_3095 ( .C (clk), .D (signal_4637), .Q (signal_4638) ) ;
    buf_clk cell_3097 ( .C (clk), .D (signal_4639), .Q (signal_4640) ) ;
    buf_clk cell_3101 ( .C (clk), .D (signal_4643), .Q (signal_4644) ) ;
    buf_clk cell_3105 ( .C (clk), .D (signal_4647), .Q (signal_4648) ) ;
    buf_clk cell_3109 ( .C (clk), .D (signal_4651), .Q (signal_4652) ) ;
    buf_clk cell_3117 ( .C (clk), .D (signal_4659), .Q (signal_4660) ) ;
    buf_clk cell_3125 ( .C (clk), .D (signal_4667), .Q (signal_4668) ) ;
    buf_clk cell_3133 ( .C (clk), .D (signal_4675), .Q (signal_4676) ) ;
    buf_clk cell_3141 ( .C (clk), .D (signal_4683), .Q (signal_4684) ) ;
    buf_clk cell_3149 ( .C (clk), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_3157 ( .C (clk), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_3165 ( .C (clk), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_3173 ( .C (clk), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_3181 ( .C (clk), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_3189 ( .C (clk), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_3197 ( .C (clk), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_3205 ( .C (clk), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_3213 ( .C (clk), .D (signal_4755), .Q (signal_4756) ) ;
    buf_clk cell_3221 ( .C (clk), .D (signal_4763), .Q (signal_4764) ) ;
    buf_clk cell_3229 ( .C (clk), .D (signal_4771), .Q (signal_4772) ) ;
    buf_clk cell_3237 ( .C (clk), .D (signal_4779), .Q (signal_4780) ) ;
    buf_clk cell_3245 ( .C (clk), .D (signal_4787), .Q (signal_4788) ) ;
    buf_clk cell_3253 ( .C (clk), .D (signal_4795), .Q (signal_4796) ) ;
    buf_clk cell_3261 ( .C (clk), .D (signal_4803), .Q (signal_4804) ) ;
    buf_clk cell_3269 ( .C (clk), .D (signal_4811), .Q (signal_4812) ) ;
    buf_clk cell_3277 ( .C (clk), .D (signal_4819), .Q (signal_4820) ) ;
    buf_clk cell_3285 ( .C (clk), .D (signal_4827), .Q (signal_4828) ) ;
    buf_clk cell_3293 ( .C (clk), .D (signal_4835), .Q (signal_4836) ) ;
    buf_clk cell_3301 ( .C (clk), .D (signal_4843), .Q (signal_4844) ) ;
    buf_clk cell_3309 ( .C (clk), .D (signal_4851), .Q (signal_4852) ) ;
    buf_clk cell_3317 ( .C (clk), .D (signal_4859), .Q (signal_4860) ) ;
    buf_clk cell_3325 ( .C (clk), .D (signal_4867), .Q (signal_4868) ) ;
    buf_clk cell_3333 ( .C (clk), .D (signal_4875), .Q (signal_4876) ) ;
    buf_clk cell_3341 ( .C (clk), .D (signal_4883), .Q (signal_4884) ) ;
    buf_clk cell_3349 ( .C (clk), .D (signal_4891), .Q (signal_4892) ) ;
    buf_clk cell_3357 ( .C (clk), .D (signal_4899), .Q (signal_4900) ) ;
    buf_clk cell_3365 ( .C (clk), .D (signal_4907), .Q (signal_4908) ) ;
    buf_clk cell_3373 ( .C (clk), .D (signal_4915), .Q (signal_4916) ) ;
    buf_clk cell_3381 ( .C (clk), .D (signal_4923), .Q (signal_4924) ) ;
    buf_clk cell_3389 ( .C (clk), .D (signal_4931), .Q (signal_4932) ) ;
    buf_clk cell_3397 ( .C (clk), .D (signal_4939), .Q (signal_4940) ) ;
    buf_clk cell_3405 ( .C (clk), .D (signal_4947), .Q (signal_4948) ) ;
    buf_clk cell_3413 ( .C (clk), .D (signal_4955), .Q (signal_4956) ) ;
    buf_clk cell_3421 ( .C (clk), .D (signal_4963), .Q (signal_4964) ) ;
    buf_clk cell_3429 ( .C (clk), .D (signal_4971), .Q (signal_4972) ) ;
    buf_clk cell_3437 ( .C (clk), .D (signal_4979), .Q (signal_4980) ) ;
    buf_clk cell_3445 ( .C (clk), .D (signal_4987), .Q (signal_4988) ) ;
    buf_clk cell_3453 ( .C (clk), .D (signal_4995), .Q (signal_4996) ) ;
    buf_clk cell_3461 ( .C (clk), .D (signal_5003), .Q (signal_5004) ) ;
    buf_clk cell_3469 ( .C (clk), .D (signal_5011), .Q (signal_5012) ) ;
    buf_clk cell_3477 ( .C (clk), .D (signal_5019), .Q (signal_5020) ) ;
    buf_clk cell_3485 ( .C (clk), .D (signal_5027), .Q (signal_5028) ) ;
    buf_clk cell_3493 ( .C (clk), .D (signal_5035), .Q (signal_5036) ) ;
    buf_clk cell_3501 ( .C (clk), .D (signal_5043), .Q (signal_5044) ) ;
    buf_clk cell_3509 ( .C (clk), .D (signal_5051), .Q (signal_5052) ) ;
    buf_clk cell_3517 ( .C (clk), .D (signal_5059), .Q (signal_5060) ) ;
    buf_clk cell_3525 ( .C (clk), .D (signal_5067), .Q (signal_5068) ) ;
    buf_clk cell_3533 ( .C (clk), .D (signal_5075), .Q (signal_5076) ) ;
    buf_clk cell_3541 ( .C (clk), .D (signal_5083), .Q (signal_5084) ) ;
    buf_clk cell_3549 ( .C (clk), .D (signal_5091), .Q (signal_5092) ) ;
    buf_clk cell_3557 ( .C (clk), .D (signal_5099), .Q (signal_5100) ) ;
    buf_clk cell_3565 ( .C (clk), .D (signal_5107), .Q (signal_5108) ) ;
    buf_clk cell_3573 ( .C (clk), .D (signal_5115), .Q (signal_5116) ) ;
    buf_clk cell_3581 ( .C (clk), .D (signal_5123), .Q (signal_5124) ) ;
    buf_clk cell_3589 ( .C (clk), .D (signal_5131), .Q (signal_5132) ) ;
    buf_clk cell_3597 ( .C (clk), .D (signal_5139), .Q (signal_5140) ) ;
    buf_clk cell_3605 ( .C (clk), .D (signal_5147), .Q (signal_5148) ) ;
    buf_clk cell_3613 ( .C (clk), .D (signal_5155), .Q (signal_5156) ) ;
    buf_clk cell_3621 ( .C (clk), .D (signal_5163), .Q (signal_5164) ) ;
    buf_clk cell_3629 ( .C (clk), .D (signal_5171), .Q (signal_5172) ) ;
    buf_clk cell_3637 ( .C (clk), .D (signal_5179), .Q (signal_5180) ) ;
    buf_clk cell_3645 ( .C (clk), .D (signal_5187), .Q (signal_5188) ) ;
    buf_clk cell_3653 ( .C (clk), .D (signal_5195), .Q (signal_5196) ) ;
    buf_clk cell_3661 ( .C (clk), .D (signal_5203), .Q (signal_5204) ) ;
    buf_clk cell_3669 ( .C (clk), .D (signal_5211), .Q (signal_5212) ) ;
    buf_clk cell_3677 ( .C (clk), .D (signal_5219), .Q (signal_5220) ) ;
    buf_clk cell_3685 ( .C (clk), .D (signal_5227), .Q (signal_5228) ) ;
    buf_clk cell_3693 ( .C (clk), .D (signal_5235), .Q (signal_5236) ) ;
    buf_clk cell_3701 ( .C (clk), .D (signal_5243), .Q (signal_5244) ) ;
    buf_clk cell_3709 ( .C (clk), .D (signal_5251), .Q (signal_5252) ) ;
    buf_clk cell_3717 ( .C (clk), .D (signal_5259), .Q (signal_5260) ) ;
    buf_clk cell_3725 ( .C (clk), .D (signal_5267), .Q (signal_5268) ) ;
    buf_clk cell_3733 ( .C (clk), .D (signal_5275), .Q (signal_5276) ) ;
    buf_clk cell_3741 ( .C (clk), .D (signal_5283), .Q (signal_5284) ) ;
    buf_clk cell_3749 ( .C (clk), .D (signal_5291), .Q (signal_5292) ) ;
    buf_clk cell_3757 ( .C (clk), .D (signal_5299), .Q (signal_5300) ) ;
    buf_clk cell_3765 ( .C (clk), .D (signal_5307), .Q (signal_5308) ) ;
    buf_clk cell_3773 ( .C (clk), .D (signal_5315), .Q (signal_5316) ) ;
    buf_clk cell_3781 ( .C (clk), .D (signal_5323), .Q (signal_5324) ) ;
    buf_clk cell_3789 ( .C (clk), .D (signal_5331), .Q (signal_5332) ) ;
    buf_clk cell_3797 ( .C (clk), .D (signal_5339), .Q (signal_5340) ) ;
    buf_clk cell_3805 ( .C (clk), .D (signal_5347), .Q (signal_5348) ) ;
    buf_clk cell_3813 ( .C (clk), .D (signal_5355), .Q (signal_5356) ) ;
    buf_clk cell_3821 ( .C (clk), .D (signal_5363), .Q (signal_5364) ) ;
    buf_clk cell_3829 ( .C (clk), .D (signal_5371), .Q (signal_5372) ) ;
    buf_clk cell_3837 ( .C (clk), .D (signal_5379), .Q (signal_5380) ) ;
    buf_clk cell_3845 ( .C (clk), .D (signal_5387), .Q (signal_5388) ) ;
    buf_clk cell_3853 ( .C (clk), .D (signal_5395), .Q (signal_5396) ) ;
    buf_clk cell_3861 ( .C (clk), .D (signal_5403), .Q (signal_5404) ) ;
    buf_clk cell_3869 ( .C (clk), .D (signal_5411), .Q (signal_5412) ) ;
    buf_clk cell_3877 ( .C (clk), .D (signal_5419), .Q (signal_5420) ) ;
    buf_clk cell_3885 ( .C (clk), .D (signal_5427), .Q (signal_5428) ) ;
    buf_clk cell_3893 ( .C (clk), .D (signal_5435), .Q (signal_5436) ) ;
    buf_clk cell_3901 ( .C (clk), .D (signal_5443), .Q (signal_5444) ) ;
    buf_clk cell_3909 ( .C (clk), .D (signal_5451), .Q (signal_5452) ) ;
    buf_clk cell_3917 ( .C (clk), .D (signal_5459), .Q (signal_5460) ) ;
    buf_clk cell_3925 ( .C (clk), .D (signal_5467), .Q (signal_5468) ) ;
    buf_clk cell_3933 ( .C (clk), .D (signal_5475), .Q (signal_5476) ) ;
    buf_clk cell_3941 ( .C (clk), .D (signal_5483), .Q (signal_5484) ) ;
    buf_clk cell_3949 ( .C (clk), .D (signal_5491), .Q (signal_5492) ) ;
    buf_clk cell_3957 ( .C (clk), .D (signal_5499), .Q (signal_5500) ) ;
    buf_clk cell_3965 ( .C (clk), .D (signal_5507), .Q (signal_5508) ) ;
    buf_clk cell_3973 ( .C (clk), .D (signal_5515), .Q (signal_5516) ) ;
    buf_clk cell_3981 ( .C (clk), .D (signal_5523), .Q (signal_5524) ) ;
    buf_clk cell_3989 ( .C (clk), .D (signal_5531), .Q (signal_5532) ) ;
    buf_clk cell_3997 ( .C (clk), .D (signal_5539), .Q (signal_5540) ) ;
    buf_clk cell_4005 ( .C (clk), .D (signal_5547), .Q (signal_5548) ) ;
    buf_clk cell_4013 ( .C (clk), .D (signal_5555), .Q (signal_5556) ) ;
    buf_clk cell_4021 ( .C (clk), .D (signal_5563), .Q (signal_5564) ) ;
    buf_clk cell_4029 ( .C (clk), .D (signal_5571), .Q (signal_5572) ) ;
    buf_clk cell_4037 ( .C (clk), .D (signal_5579), .Q (signal_5580) ) ;
    buf_clk cell_4045 ( .C (clk), .D (signal_5587), .Q (signal_5588) ) ;
    buf_clk cell_4053 ( .C (clk), .D (signal_5595), .Q (signal_5596) ) ;
    buf_clk cell_4061 ( .C (clk), .D (signal_5603), .Q (signal_5604) ) ;
    buf_clk cell_4069 ( .C (clk), .D (signal_5611), .Q (signal_5612) ) ;
    buf_clk cell_4077 ( .C (clk), .D (signal_5619), .Q (signal_5620) ) ;
    buf_clk cell_4085 ( .C (clk), .D (signal_5627), .Q (signal_5628) ) ;
    buf_clk cell_4093 ( .C (clk), .D (signal_5635), .Q (signal_5636) ) ;
    buf_clk cell_4101 ( .C (clk), .D (signal_5643), .Q (signal_5644) ) ;
    buf_clk cell_4109 ( .C (clk), .D (signal_5651), .Q (signal_5652) ) ;
    buf_clk cell_4117 ( .C (clk), .D (signal_5659), .Q (signal_5660) ) ;
    buf_clk cell_4125 ( .C (clk), .D (signal_5667), .Q (signal_5668) ) ;
    buf_clk cell_4135 ( .C (clk), .D (signal_5677), .Q (signal_5678) ) ;
    buf_clk cell_4143 ( .C (clk), .D (signal_5685), .Q (signal_5686) ) ;
    buf_clk cell_4151 ( .C (clk), .D (signal_5693), .Q (signal_5694) ) ;
    buf_clk cell_4159 ( .C (clk), .D (signal_5701), .Q (signal_5702) ) ;
    buf_clk cell_4167 ( .C (clk), .D (signal_5709), .Q (signal_5710) ) ;
    buf_clk cell_4175 ( .C (clk), .D (signal_5717), .Q (signal_5718) ) ;
    buf_clk cell_4183 ( .C (clk), .D (signal_5725), .Q (signal_5726) ) ;
    buf_clk cell_4191 ( .C (clk), .D (signal_5733), .Q (signal_5734) ) ;
    buf_clk cell_4199 ( .C (clk), .D (signal_5741), .Q (signal_5742) ) ;
    buf_clk cell_4207 ( .C (clk), .D (signal_5749), .Q (signal_5750) ) ;
    buf_clk cell_4215 ( .C (clk), .D (signal_5757), .Q (signal_5758) ) ;
    buf_clk cell_4223 ( .C (clk), .D (signal_5765), .Q (signal_5766) ) ;
    buf_clk cell_4231 ( .C (clk), .D (signal_5773), .Q (signal_5774) ) ;
    buf_clk cell_4239 ( .C (clk), .D (signal_5781), .Q (signal_5782) ) ;
    buf_clk cell_4247 ( .C (clk), .D (signal_5789), .Q (signal_5790) ) ;
    buf_clk cell_4255 ( .C (clk), .D (signal_5797), .Q (signal_5798) ) ;
    buf_clk cell_4263 ( .C (clk), .D (signal_5805), .Q (signal_5806) ) ;
    buf_clk cell_4271 ( .C (clk), .D (signal_5813), .Q (signal_5814) ) ;
    buf_clk cell_4279 ( .C (clk), .D (signal_5821), .Q (signal_5822) ) ;
    buf_clk cell_4287 ( .C (clk), .D (signal_5829), .Q (signal_5830) ) ;
    buf_clk cell_4295 ( .C (clk), .D (signal_5837), .Q (signal_5838) ) ;
    buf_clk cell_4303 ( .C (clk), .D (signal_5845), .Q (signal_5846) ) ;
    buf_clk cell_4311 ( .C (clk), .D (signal_5853), .Q (signal_5854) ) ;
    buf_clk cell_4319 ( .C (clk), .D (signal_5861), .Q (signal_5862) ) ;
    buf_clk cell_4327 ( .C (clk), .D (signal_5869), .Q (signal_5870) ) ;
    buf_clk cell_4335 ( .C (clk), .D (signal_5877), .Q (signal_5878) ) ;
    buf_clk cell_4343 ( .C (clk), .D (signal_5885), .Q (signal_5886) ) ;
    buf_clk cell_4351 ( .C (clk), .D (signal_5893), .Q (signal_5894) ) ;
    buf_clk cell_4359 ( .C (clk), .D (signal_5901), .Q (signal_5902) ) ;
    buf_clk cell_4367 ( .C (clk), .D (signal_5909), .Q (signal_5910) ) ;
    buf_clk cell_4375 ( .C (clk), .D (signal_5917), .Q (signal_5918) ) ;
    buf_clk cell_4383 ( .C (clk), .D (signal_5925), .Q (signal_5926) ) ;
    buf_clk cell_4391 ( .C (clk), .D (signal_5933), .Q (signal_5934) ) ;
    buf_clk cell_4399 ( .C (clk), .D (signal_5941), .Q (signal_5942) ) ;
    buf_clk cell_4407 ( .C (clk), .D (signal_5949), .Q (signal_5950) ) ;
    buf_clk cell_4415 ( .C (clk), .D (signal_5957), .Q (signal_5958) ) ;
    buf_clk cell_4423 ( .C (clk), .D (signal_5965), .Q (signal_5966) ) ;
    buf_clk cell_4431 ( .C (clk), .D (signal_5973), .Q (signal_5974) ) ;
    buf_clk cell_4439 ( .C (clk), .D (signal_5981), .Q (signal_5982) ) ;
    buf_clk cell_4447 ( .C (clk), .D (signal_5989), .Q (signal_5990) ) ;
    buf_clk cell_4455 ( .C (clk), .D (signal_5997), .Q (signal_5998) ) ;
    buf_clk cell_4463 ( .C (clk), .D (signal_6005), .Q (signal_6006) ) ;
    buf_clk cell_4471 ( .C (clk), .D (signal_6013), .Q (signal_6014) ) ;
    buf_clk cell_4479 ( .C (clk), .D (signal_6021), .Q (signal_6022) ) ;
    buf_clk cell_4487 ( .C (clk), .D (signal_6029), .Q (signal_6030) ) ;
    buf_clk cell_4495 ( .C (clk), .D (signal_6037), .Q (signal_6038) ) ;
    buf_clk cell_4503 ( .C (clk), .D (signal_6045), .Q (signal_6046) ) ;
    buf_clk cell_4511 ( .C (clk), .D (signal_6053), .Q (signal_6054) ) ;
    buf_clk cell_4519 ( .C (clk), .D (signal_6061), .Q (signal_6062) ) ;
    buf_clk cell_4527 ( .C (clk), .D (signal_6069), .Q (signal_6070) ) ;
    buf_clk cell_4535 ( .C (clk), .D (signal_6077), .Q (signal_6078) ) ;
    buf_clk cell_4543 ( .C (clk), .D (signal_6085), .Q (signal_6086) ) ;
    buf_clk cell_4551 ( .C (clk), .D (signal_6093), .Q (signal_6094) ) ;
    buf_clk cell_4559 ( .C (clk), .D (signal_6101), .Q (signal_6102) ) ;
    buf_clk cell_4567 ( .C (clk), .D (signal_6109), .Q (signal_6110) ) ;
    buf_clk cell_4575 ( .C (clk), .D (signal_6117), .Q (signal_6118) ) ;
    buf_clk cell_4583 ( .C (clk), .D (signal_6125), .Q (signal_6126) ) ;
    buf_clk cell_4591 ( .C (clk), .D (signal_6133), .Q (signal_6134) ) ;
    buf_clk cell_4599 ( .C (clk), .D (signal_6141), .Q (signal_6142) ) ;
    buf_clk cell_4607 ( .C (clk), .D (signal_6149), .Q (signal_6150) ) ;
    buf_clk cell_4615 ( .C (clk), .D (signal_6157), .Q (signal_6158) ) ;
    buf_clk cell_4623 ( .C (clk), .D (signal_6165), .Q (signal_6166) ) ;
    buf_clk cell_4631 ( .C (clk), .D (signal_6173), .Q (signal_6174) ) ;
    buf_clk cell_4639 ( .C (clk), .D (signal_6181), .Q (signal_6182) ) ;
    buf_clk cell_4841 ( .C (clk), .D (signal_6383), .Q (signal_6384) ) ;
    buf_clk cell_4849 ( .C (clk), .D (signal_6391), .Q (signal_6392) ) ;
    buf_clk cell_4857 ( .C (clk), .D (signal_6399), .Q (signal_6400) ) ;
    buf_clk cell_4865 ( .C (clk), .D (signal_6407), .Q (signal_6408) ) ;

    /* cells in depth 5 */
    buf_clk cell_1554 ( .C (clk), .D (signal_3096), .Q (signal_3097) ) ;
    buf_clk cell_1754 ( .C (clk), .D (signal_3296), .Q (signal_3297) ) ;
    buf_clk cell_1760 ( .C (clk), .D (signal_3302), .Q (signal_3303) ) ;
    buf_clk cell_1766 ( .C (clk), .D (signal_3308), .Q (signal_3309) ) ;
    buf_clk cell_1772 ( .C (clk), .D (signal_3314), .Q (signal_3315) ) ;
    buf_clk cell_1778 ( .C (clk), .D (signal_3320), .Q (signal_3321) ) ;
    buf_clk cell_1784 ( .C (clk), .D (signal_3326), .Q (signal_3327) ) ;
    buf_clk cell_1790 ( .C (clk), .D (signal_3332), .Q (signal_3333) ) ;
    buf_clk cell_1796 ( .C (clk), .D (signal_3338), .Q (signal_3339) ) ;
    buf_clk cell_1802 ( .C (clk), .D (signal_3344), .Q (signal_3345) ) ;
    buf_clk cell_1808 ( .C (clk), .D (signal_3350), .Q (signal_3351) ) ;
    buf_clk cell_1814 ( .C (clk), .D (signal_3356), .Q (signal_3357) ) ;
    buf_clk cell_1820 ( .C (clk), .D (signal_3362), .Q (signal_3363) ) ;
    buf_clk cell_1826 ( .C (clk), .D (signal_3368), .Q (signal_3369) ) ;
    buf_clk cell_1832 ( .C (clk), .D (signal_3374), .Q (signal_3375) ) ;
    buf_clk cell_1838 ( .C (clk), .D (signal_3380), .Q (signal_3381) ) ;
    buf_clk cell_1844 ( .C (clk), .D (signal_3386), .Q (signal_3387) ) ;
    buf_clk cell_1850 ( .C (clk), .D (signal_3392), .Q (signal_3393) ) ;
    buf_clk cell_1856 ( .C (clk), .D (signal_3398), .Q (signal_3399) ) ;
    buf_clk cell_1862 ( .C (clk), .D (signal_3404), .Q (signal_3405) ) ;
    buf_clk cell_1868 ( .C (clk), .D (signal_3410), .Q (signal_3411) ) ;
    buf_clk cell_1874 ( .C (clk), .D (signal_3416), .Q (signal_3417) ) ;
    buf_clk cell_1880 ( .C (clk), .D (signal_3422), .Q (signal_3423) ) ;
    buf_clk cell_1886 ( .C (clk), .D (signal_3428), .Q (signal_3429) ) ;
    buf_clk cell_1892 ( .C (clk), .D (signal_3434), .Q (signal_3435) ) ;
    buf_clk cell_1898 ( .C (clk), .D (signal_3440), .Q (signal_3441) ) ;
    buf_clk cell_1904 ( .C (clk), .D (signal_3446), .Q (signal_3447) ) ;
    buf_clk cell_1910 ( .C (clk), .D (signal_3452), .Q (signal_3453) ) ;
    buf_clk cell_1916 ( .C (clk), .D (signal_3458), .Q (signal_3459) ) ;
    buf_clk cell_1922 ( .C (clk), .D (signal_3464), .Q (signal_3465) ) ;
    buf_clk cell_1928 ( .C (clk), .D (signal_3470), .Q (signal_3471) ) ;
    buf_clk cell_1934 ( .C (clk), .D (signal_3476), .Q (signal_3477) ) ;
    buf_clk cell_1940 ( .C (clk), .D (signal_3482), .Q (signal_3483) ) ;
    buf_clk cell_1946 ( .C (clk), .D (signal_3488), .Q (signal_3489) ) ;
    buf_clk cell_1952 ( .C (clk), .D (signal_3494), .Q (signal_3495) ) ;
    buf_clk cell_1958 ( .C (clk), .D (signal_3500), .Q (signal_3501) ) ;
    buf_clk cell_1964 ( .C (clk), .D (signal_3506), .Q (signal_3507) ) ;
    buf_clk cell_1970 ( .C (clk), .D (signal_3512), .Q (signal_3513) ) ;
    buf_clk cell_1976 ( .C (clk), .D (signal_3518), .Q (signal_3519) ) ;
    buf_clk cell_1982 ( .C (clk), .D (signal_3524), .Q (signal_3525) ) ;
    buf_clk cell_1988 ( .C (clk), .D (signal_3530), .Q (signal_3531) ) ;
    buf_clk cell_1994 ( .C (clk), .D (signal_3536), .Q (signal_3537) ) ;
    buf_clk cell_2000 ( .C (clk), .D (signal_3542), .Q (signal_3543) ) ;
    buf_clk cell_2006 ( .C (clk), .D (signal_3548), .Q (signal_3549) ) ;
    buf_clk cell_2012 ( .C (clk), .D (signal_3554), .Q (signal_3555) ) ;
    buf_clk cell_2018 ( .C (clk), .D (signal_3560), .Q (signal_3561) ) ;
    buf_clk cell_2024 ( .C (clk), .D (signal_3566), .Q (signal_3567) ) ;
    buf_clk cell_2030 ( .C (clk), .D (signal_3572), .Q (signal_3573) ) ;
    buf_clk cell_2036 ( .C (clk), .D (signal_3578), .Q (signal_3579) ) ;
    buf_clk cell_2042 ( .C (clk), .D (signal_3584), .Q (signal_3585) ) ;
    buf_clk cell_2048 ( .C (clk), .D (signal_3590), .Q (signal_3591) ) ;
    buf_clk cell_2054 ( .C (clk), .D (signal_3596), .Q (signal_3597) ) ;
    buf_clk cell_2060 ( .C (clk), .D (signal_3602), .Q (signal_3603) ) ;
    buf_clk cell_2066 ( .C (clk), .D (signal_3608), .Q (signal_3609) ) ;
    buf_clk cell_2072 ( .C (clk), .D (signal_3614), .Q (signal_3615) ) ;
    buf_clk cell_2078 ( .C (clk), .D (signal_3620), .Q (signal_3621) ) ;
    buf_clk cell_2084 ( .C (clk), .D (signal_3626), .Q (signal_3627) ) ;
    buf_clk cell_2090 ( .C (clk), .D (signal_3632), .Q (signal_3633) ) ;
    buf_clk cell_2096 ( .C (clk), .D (signal_3638), .Q (signal_3639) ) ;
    buf_clk cell_2102 ( .C (clk), .D (signal_3644), .Q (signal_3645) ) ;
    buf_clk cell_2108 ( .C (clk), .D (signal_3650), .Q (signal_3651) ) ;
    buf_clk cell_2114 ( .C (clk), .D (signal_3656), .Q (signal_3657) ) ;
    buf_clk cell_2120 ( .C (clk), .D (signal_3662), .Q (signal_3663) ) ;
    buf_clk cell_2126 ( .C (clk), .D (signal_3668), .Q (signal_3669) ) ;
    buf_clk cell_2132 ( .C (clk), .D (signal_3674), .Q (signal_3675) ) ;
    buf_clk cell_2138 ( .C (clk), .D (signal_3680), .Q (signal_3681) ) ;
    buf_clk cell_2144 ( .C (clk), .D (signal_3686), .Q (signal_3687) ) ;
    buf_clk cell_2150 ( .C (clk), .D (signal_3692), .Q (signal_3693) ) ;
    buf_clk cell_2156 ( .C (clk), .D (signal_3698), .Q (signal_3699) ) ;
    buf_clk cell_2162 ( .C (clk), .D (signal_3704), .Q (signal_3705) ) ;
    buf_clk cell_2168 ( .C (clk), .D (signal_3710), .Q (signal_3711) ) ;
    buf_clk cell_2174 ( .C (clk), .D (signal_3716), .Q (signal_3717) ) ;
    buf_clk cell_2180 ( .C (clk), .D (signal_3722), .Q (signal_3723) ) ;
    buf_clk cell_2186 ( .C (clk), .D (signal_3728), .Q (signal_3729) ) ;
    buf_clk cell_2192 ( .C (clk), .D (signal_3734), .Q (signal_3735) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_3740), .Q (signal_3741) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_3746), .Q (signal_3747) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_3752), .Q (signal_3753) ) ;
    buf_clk cell_2216 ( .C (clk), .D (signal_3758), .Q (signal_3759) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_3764), .Q (signal_3765) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_3770), .Q (signal_3771) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_3776), .Q (signal_3777) ) ;
    buf_clk cell_2240 ( .C (clk), .D (signal_3782), .Q (signal_3783) ) ;
    buf_clk cell_2246 ( .C (clk), .D (signal_3788), .Q (signal_3789) ) ;
    buf_clk cell_2252 ( .C (clk), .D (signal_3794), .Q (signal_3795) ) ;
    buf_clk cell_2258 ( .C (clk), .D (signal_3800), .Q (signal_3801) ) ;
    buf_clk cell_2264 ( .C (clk), .D (signal_3806), .Q (signal_3807) ) ;
    buf_clk cell_2270 ( .C (clk), .D (signal_3812), .Q (signal_3813) ) ;
    buf_clk cell_2276 ( .C (clk), .D (signal_3818), .Q (signal_3819) ) ;
    buf_clk cell_2282 ( .C (clk), .D (signal_3824), .Q (signal_3825) ) ;
    buf_clk cell_2288 ( .C (clk), .D (signal_3830), .Q (signal_3831) ) ;
    buf_clk cell_2294 ( .C (clk), .D (signal_3836), .Q (signal_3837) ) ;
    buf_clk cell_2300 ( .C (clk), .D (signal_3842), .Q (signal_3843) ) ;
    buf_clk cell_2306 ( .C (clk), .D (signal_3848), .Q (signal_3849) ) ;
    buf_clk cell_2312 ( .C (clk), .D (signal_3854), .Q (signal_3855) ) ;
    buf_clk cell_2318 ( .C (clk), .D (signal_3860), .Q (signal_3861) ) ;
    buf_clk cell_2324 ( .C (clk), .D (signal_3866), .Q (signal_3867) ) ;
    buf_clk cell_2330 ( .C (clk), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_2336 ( .C (clk), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_2342 ( .C (clk), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_2348 ( .C (clk), .D (signal_3890), .Q (signal_3891) ) ;
    buf_clk cell_2354 ( .C (clk), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_2360 ( .C (clk), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_2366 ( .C (clk), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_2372 ( .C (clk), .D (signal_3914), .Q (signal_3915) ) ;
    buf_clk cell_2378 ( .C (clk), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_2384 ( .C (clk), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_2390 ( .C (clk), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_2396 ( .C (clk), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_2402 ( .C (clk), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_2408 ( .C (clk), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_2414 ( .C (clk), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_2420 ( .C (clk), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_2426 ( .C (clk), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_2432 ( .C (clk), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_2438 ( .C (clk), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_2444 ( .C (clk), .D (signal_3986), .Q (signal_3987) ) ;
    buf_clk cell_2450 ( .C (clk), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_2456 ( .C (clk), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_2462 ( .C (clk), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_2468 ( .C (clk), .D (signal_4010), .Q (signal_4011) ) ;
    buf_clk cell_2474 ( .C (clk), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_2480 ( .C (clk), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_2486 ( .C (clk), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_2492 ( .C (clk), .D (signal_4034), .Q (signal_4035) ) ;
    buf_clk cell_2498 ( .C (clk), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_2504 ( .C (clk), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_2510 ( .C (clk), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_2516 ( .C (clk), .D (signal_4058), .Q (signal_4059) ) ;
    buf_clk cell_2522 ( .C (clk), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_2528 ( .C (clk), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_2534 ( .C (clk), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_2540 ( .C (clk), .D (signal_4082), .Q (signal_4083) ) ;
    buf_clk cell_2546 ( .C (clk), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_2552 ( .C (clk), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_2558 ( .C (clk), .D (signal_4100), .Q (signal_4101) ) ;
    buf_clk cell_2564 ( .C (clk), .D (signal_4106), .Q (signal_4107) ) ;
    buf_clk cell_2570 ( .C (clk), .D (signal_4112), .Q (signal_4113) ) ;
    buf_clk cell_2576 ( .C (clk), .D (signal_4118), .Q (signal_4119) ) ;
    buf_clk cell_2582 ( .C (clk), .D (signal_4124), .Q (signal_4125) ) ;
    buf_clk cell_2588 ( .C (clk), .D (signal_4130), .Q (signal_4131) ) ;
    buf_clk cell_2594 ( .C (clk), .D (signal_4136), .Q (signal_4137) ) ;
    buf_clk cell_2600 ( .C (clk), .D (signal_4142), .Q (signal_4143) ) ;
    buf_clk cell_2606 ( .C (clk), .D (signal_4148), .Q (signal_4149) ) ;
    buf_clk cell_2612 ( .C (clk), .D (signal_4154), .Q (signal_4155) ) ;
    buf_clk cell_2618 ( .C (clk), .D (signal_4160), .Q (signal_4161) ) ;
    buf_clk cell_2624 ( .C (clk), .D (signal_4166), .Q (signal_4167) ) ;
    buf_clk cell_2630 ( .C (clk), .D (signal_4172), .Q (signal_4173) ) ;
    buf_clk cell_2636 ( .C (clk), .D (signal_4178), .Q (signal_4179) ) ;
    buf_clk cell_2642 ( .C (clk), .D (signal_4184), .Q (signal_4185) ) ;
    buf_clk cell_2648 ( .C (clk), .D (signal_4190), .Q (signal_4191) ) ;
    buf_clk cell_2654 ( .C (clk), .D (signal_4196), .Q (signal_4197) ) ;
    buf_clk cell_2660 ( .C (clk), .D (signal_4202), .Q (signal_4203) ) ;
    buf_clk cell_2666 ( .C (clk), .D (signal_4208), .Q (signal_4209) ) ;
    buf_clk cell_2672 ( .C (clk), .D (signal_4214), .Q (signal_4215) ) ;
    buf_clk cell_2678 ( .C (clk), .D (signal_4220), .Q (signal_4221) ) ;
    buf_clk cell_2684 ( .C (clk), .D (signal_4226), .Q (signal_4227) ) ;
    buf_clk cell_2690 ( .C (clk), .D (signal_4232), .Q (signal_4233) ) ;
    buf_clk cell_2696 ( .C (clk), .D (signal_4238), .Q (signal_4239) ) ;
    buf_clk cell_2702 ( .C (clk), .D (signal_4244), .Q (signal_4245) ) ;
    buf_clk cell_2708 ( .C (clk), .D (signal_4250), .Q (signal_4251) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_4256), .Q (signal_4257) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_4262), .Q (signal_4263) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_4268), .Q (signal_4269) ) ;
    buf_clk cell_2732 ( .C (clk), .D (signal_4274), .Q (signal_4275) ) ;
    buf_clk cell_2738 ( .C (clk), .D (signal_4280), .Q (signal_4281) ) ;
    buf_clk cell_2744 ( .C (clk), .D (signal_4286), .Q (signal_4287) ) ;
    buf_clk cell_2750 ( .C (clk), .D (signal_4292), .Q (signal_4293) ) ;
    buf_clk cell_2756 ( .C (clk), .D (signal_4298), .Q (signal_4299) ) ;
    buf_clk cell_2762 ( .C (clk), .D (signal_4304), .Q (signal_4305) ) ;
    buf_clk cell_2768 ( .C (clk), .D (signal_4310), .Q (signal_4311) ) ;
    buf_clk cell_2774 ( .C (clk), .D (signal_4316), .Q (signal_4317) ) ;
    buf_clk cell_2780 ( .C (clk), .D (signal_4322), .Q (signal_4323) ) ;
    buf_clk cell_2786 ( .C (clk), .D (signal_4328), .Q (signal_4329) ) ;
    buf_clk cell_2792 ( .C (clk), .D (signal_4334), .Q (signal_4335) ) ;
    buf_clk cell_2798 ( .C (clk), .D (signal_4340), .Q (signal_4341) ) ;
    buf_clk cell_2804 ( .C (clk), .D (signal_4346), .Q (signal_4347) ) ;
    buf_clk cell_2810 ( .C (clk), .D (signal_4352), .Q (signal_4353) ) ;
    buf_clk cell_2816 ( .C (clk), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_2822 ( .C (clk), .D (signal_4364), .Q (signal_4365) ) ;
    buf_clk cell_2828 ( .C (clk), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_2834 ( .C (clk), .D (signal_4376), .Q (signal_4377) ) ;
    buf_clk cell_2840 ( .C (clk), .D (signal_4382), .Q (signal_4383) ) ;
    buf_clk cell_2846 ( .C (clk), .D (signal_4388), .Q (signal_4389) ) ;
    buf_clk cell_2852 ( .C (clk), .D (signal_4394), .Q (signal_4395) ) ;
    buf_clk cell_2858 ( .C (clk), .D (signal_4400), .Q (signal_4401) ) ;
    buf_clk cell_2864 ( .C (clk), .D (signal_4406), .Q (signal_4407) ) ;
    buf_clk cell_2870 ( .C (clk), .D (signal_4412), .Q (signal_4413) ) ;
    buf_clk cell_2876 ( .C (clk), .D (signal_4418), .Q (signal_4419) ) ;
    buf_clk cell_2882 ( .C (clk), .D (signal_4424), .Q (signal_4425) ) ;
    buf_clk cell_2888 ( .C (clk), .D (signal_4430), .Q (signal_4431) ) ;
    buf_clk cell_2894 ( .C (clk), .D (signal_4436), .Q (signal_4437) ) ;
    buf_clk cell_2900 ( .C (clk), .D (signal_4442), .Q (signal_4443) ) ;
    buf_clk cell_2906 ( .C (clk), .D (signal_4448), .Q (signal_4449) ) ;
    buf_clk cell_2912 ( .C (clk), .D (signal_4454), .Q (signal_4455) ) ;
    buf_clk cell_3110 ( .C (clk), .D (signal_4652), .Q (signal_4653) ) ;
    buf_clk cell_3118 ( .C (clk), .D (signal_4660), .Q (signal_4661) ) ;
    buf_clk cell_3126 ( .C (clk), .D (signal_4668), .Q (signal_4669) ) ;
    buf_clk cell_3134 ( .C (clk), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_3142 ( .C (clk), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_3150 ( .C (clk), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_3158 ( .C (clk), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_3166 ( .C (clk), .D (signal_4708), .Q (signal_4709) ) ;
    buf_clk cell_3174 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_3182 ( .C (clk), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_3190 ( .C (clk), .D (signal_4732), .Q (signal_4733) ) ;
    buf_clk cell_3198 ( .C (clk), .D (signal_4740), .Q (signal_4741) ) ;
    buf_clk cell_3206 ( .C (clk), .D (signal_4748), .Q (signal_4749) ) ;
    buf_clk cell_3214 ( .C (clk), .D (signal_4756), .Q (signal_4757) ) ;
    buf_clk cell_3222 ( .C (clk), .D (signal_4764), .Q (signal_4765) ) ;
    buf_clk cell_3230 ( .C (clk), .D (signal_4772), .Q (signal_4773) ) ;
    buf_clk cell_3238 ( .C (clk), .D (signal_4780), .Q (signal_4781) ) ;
    buf_clk cell_3246 ( .C (clk), .D (signal_4788), .Q (signal_4789) ) ;
    buf_clk cell_3254 ( .C (clk), .D (signal_4796), .Q (signal_4797) ) ;
    buf_clk cell_3262 ( .C (clk), .D (signal_4804), .Q (signal_4805) ) ;
    buf_clk cell_3270 ( .C (clk), .D (signal_4812), .Q (signal_4813) ) ;
    buf_clk cell_3278 ( .C (clk), .D (signal_4820), .Q (signal_4821) ) ;
    buf_clk cell_3286 ( .C (clk), .D (signal_4828), .Q (signal_4829) ) ;
    buf_clk cell_3294 ( .C (clk), .D (signal_4836), .Q (signal_4837) ) ;
    buf_clk cell_3302 ( .C (clk), .D (signal_4844), .Q (signal_4845) ) ;
    buf_clk cell_3310 ( .C (clk), .D (signal_4852), .Q (signal_4853) ) ;
    buf_clk cell_3318 ( .C (clk), .D (signal_4860), .Q (signal_4861) ) ;
    buf_clk cell_3326 ( .C (clk), .D (signal_4868), .Q (signal_4869) ) ;
    buf_clk cell_3334 ( .C (clk), .D (signal_4876), .Q (signal_4877) ) ;
    buf_clk cell_3342 ( .C (clk), .D (signal_4884), .Q (signal_4885) ) ;
    buf_clk cell_3350 ( .C (clk), .D (signal_4892), .Q (signal_4893) ) ;
    buf_clk cell_3358 ( .C (clk), .D (signal_4900), .Q (signal_4901) ) ;
    buf_clk cell_3366 ( .C (clk), .D (signal_4908), .Q (signal_4909) ) ;
    buf_clk cell_3374 ( .C (clk), .D (signal_4916), .Q (signal_4917) ) ;
    buf_clk cell_3382 ( .C (clk), .D (signal_4924), .Q (signal_4925) ) ;
    buf_clk cell_3390 ( .C (clk), .D (signal_4932), .Q (signal_4933) ) ;
    buf_clk cell_3398 ( .C (clk), .D (signal_4940), .Q (signal_4941) ) ;
    buf_clk cell_3406 ( .C (clk), .D (signal_4948), .Q (signal_4949) ) ;
    buf_clk cell_3414 ( .C (clk), .D (signal_4956), .Q (signal_4957) ) ;
    buf_clk cell_3422 ( .C (clk), .D (signal_4964), .Q (signal_4965) ) ;
    buf_clk cell_3430 ( .C (clk), .D (signal_4972), .Q (signal_4973) ) ;
    buf_clk cell_3438 ( .C (clk), .D (signal_4980), .Q (signal_4981) ) ;
    buf_clk cell_3446 ( .C (clk), .D (signal_4988), .Q (signal_4989) ) ;
    buf_clk cell_3454 ( .C (clk), .D (signal_4996), .Q (signal_4997) ) ;
    buf_clk cell_3462 ( .C (clk), .D (signal_5004), .Q (signal_5005) ) ;
    buf_clk cell_3470 ( .C (clk), .D (signal_5012), .Q (signal_5013) ) ;
    buf_clk cell_3478 ( .C (clk), .D (signal_5020), .Q (signal_5021) ) ;
    buf_clk cell_3486 ( .C (clk), .D (signal_5028), .Q (signal_5029) ) ;
    buf_clk cell_3494 ( .C (clk), .D (signal_5036), .Q (signal_5037) ) ;
    buf_clk cell_3502 ( .C (clk), .D (signal_5044), .Q (signal_5045) ) ;
    buf_clk cell_3510 ( .C (clk), .D (signal_5052), .Q (signal_5053) ) ;
    buf_clk cell_3518 ( .C (clk), .D (signal_5060), .Q (signal_5061) ) ;
    buf_clk cell_3526 ( .C (clk), .D (signal_5068), .Q (signal_5069) ) ;
    buf_clk cell_3534 ( .C (clk), .D (signal_5076), .Q (signal_5077) ) ;
    buf_clk cell_3542 ( .C (clk), .D (signal_5084), .Q (signal_5085) ) ;
    buf_clk cell_3550 ( .C (clk), .D (signal_5092), .Q (signal_5093) ) ;
    buf_clk cell_3558 ( .C (clk), .D (signal_5100), .Q (signal_5101) ) ;
    buf_clk cell_3566 ( .C (clk), .D (signal_5108), .Q (signal_5109) ) ;
    buf_clk cell_3574 ( .C (clk), .D (signal_5116), .Q (signal_5117) ) ;
    buf_clk cell_3582 ( .C (clk), .D (signal_5124), .Q (signal_5125) ) ;
    buf_clk cell_3590 ( .C (clk), .D (signal_5132), .Q (signal_5133) ) ;
    buf_clk cell_3598 ( .C (clk), .D (signal_5140), .Q (signal_5141) ) ;
    buf_clk cell_3606 ( .C (clk), .D (signal_5148), .Q (signal_5149) ) ;
    buf_clk cell_3614 ( .C (clk), .D (signal_5156), .Q (signal_5157) ) ;
    buf_clk cell_3622 ( .C (clk), .D (signal_5164), .Q (signal_5165) ) ;
    buf_clk cell_3630 ( .C (clk), .D (signal_5172), .Q (signal_5173) ) ;
    buf_clk cell_3638 ( .C (clk), .D (signal_5180), .Q (signal_5181) ) ;
    buf_clk cell_3646 ( .C (clk), .D (signal_5188), .Q (signal_5189) ) ;
    buf_clk cell_3654 ( .C (clk), .D (signal_5196), .Q (signal_5197) ) ;
    buf_clk cell_3662 ( .C (clk), .D (signal_5204), .Q (signal_5205) ) ;
    buf_clk cell_3670 ( .C (clk), .D (signal_5212), .Q (signal_5213) ) ;
    buf_clk cell_3678 ( .C (clk), .D (signal_5220), .Q (signal_5221) ) ;
    buf_clk cell_3686 ( .C (clk), .D (signal_5228), .Q (signal_5229) ) ;
    buf_clk cell_3694 ( .C (clk), .D (signal_5236), .Q (signal_5237) ) ;
    buf_clk cell_3702 ( .C (clk), .D (signal_5244), .Q (signal_5245) ) ;
    buf_clk cell_3710 ( .C (clk), .D (signal_5252), .Q (signal_5253) ) ;
    buf_clk cell_3718 ( .C (clk), .D (signal_5260), .Q (signal_5261) ) ;
    buf_clk cell_3726 ( .C (clk), .D (signal_5268), .Q (signal_5269) ) ;
    buf_clk cell_3734 ( .C (clk), .D (signal_5276), .Q (signal_5277) ) ;
    buf_clk cell_3742 ( .C (clk), .D (signal_5284), .Q (signal_5285) ) ;
    buf_clk cell_3750 ( .C (clk), .D (signal_5292), .Q (signal_5293) ) ;
    buf_clk cell_3758 ( .C (clk), .D (signal_5300), .Q (signal_5301) ) ;
    buf_clk cell_3766 ( .C (clk), .D (signal_5308), .Q (signal_5309) ) ;
    buf_clk cell_3774 ( .C (clk), .D (signal_5316), .Q (signal_5317) ) ;
    buf_clk cell_3782 ( .C (clk), .D (signal_5324), .Q (signal_5325) ) ;
    buf_clk cell_3790 ( .C (clk), .D (signal_5332), .Q (signal_5333) ) ;
    buf_clk cell_3798 ( .C (clk), .D (signal_5340), .Q (signal_5341) ) ;
    buf_clk cell_3806 ( .C (clk), .D (signal_5348), .Q (signal_5349) ) ;
    buf_clk cell_3814 ( .C (clk), .D (signal_5356), .Q (signal_5357) ) ;
    buf_clk cell_3822 ( .C (clk), .D (signal_5364), .Q (signal_5365) ) ;
    buf_clk cell_3830 ( .C (clk), .D (signal_5372), .Q (signal_5373) ) ;
    buf_clk cell_3838 ( .C (clk), .D (signal_5380), .Q (signal_5381) ) ;
    buf_clk cell_3846 ( .C (clk), .D (signal_5388), .Q (signal_5389) ) ;
    buf_clk cell_3854 ( .C (clk), .D (signal_5396), .Q (signal_5397) ) ;
    buf_clk cell_3862 ( .C (clk), .D (signal_5404), .Q (signal_5405) ) ;
    buf_clk cell_3870 ( .C (clk), .D (signal_5412), .Q (signal_5413) ) ;
    buf_clk cell_3878 ( .C (clk), .D (signal_5420), .Q (signal_5421) ) ;
    buf_clk cell_3886 ( .C (clk), .D (signal_5428), .Q (signal_5429) ) ;
    buf_clk cell_3894 ( .C (clk), .D (signal_5436), .Q (signal_5437) ) ;
    buf_clk cell_3902 ( .C (clk), .D (signal_5444), .Q (signal_5445) ) ;
    buf_clk cell_3910 ( .C (clk), .D (signal_5452), .Q (signal_5453) ) ;
    buf_clk cell_3918 ( .C (clk), .D (signal_5460), .Q (signal_5461) ) ;
    buf_clk cell_3926 ( .C (clk), .D (signal_5468), .Q (signal_5469) ) ;
    buf_clk cell_3934 ( .C (clk), .D (signal_5476), .Q (signal_5477) ) ;
    buf_clk cell_3942 ( .C (clk), .D (signal_5484), .Q (signal_5485) ) ;
    buf_clk cell_3950 ( .C (clk), .D (signal_5492), .Q (signal_5493) ) ;
    buf_clk cell_3958 ( .C (clk), .D (signal_5500), .Q (signal_5501) ) ;
    buf_clk cell_3966 ( .C (clk), .D (signal_5508), .Q (signal_5509) ) ;
    buf_clk cell_3974 ( .C (clk), .D (signal_5516), .Q (signal_5517) ) ;
    buf_clk cell_3982 ( .C (clk), .D (signal_5524), .Q (signal_5525) ) ;
    buf_clk cell_3990 ( .C (clk), .D (signal_5532), .Q (signal_5533) ) ;
    buf_clk cell_3998 ( .C (clk), .D (signal_5540), .Q (signal_5541) ) ;
    buf_clk cell_4006 ( .C (clk), .D (signal_5548), .Q (signal_5549) ) ;
    buf_clk cell_4014 ( .C (clk), .D (signal_5556), .Q (signal_5557) ) ;
    buf_clk cell_4022 ( .C (clk), .D (signal_5564), .Q (signal_5565) ) ;
    buf_clk cell_4030 ( .C (clk), .D (signal_5572), .Q (signal_5573) ) ;
    buf_clk cell_4038 ( .C (clk), .D (signal_5580), .Q (signal_5581) ) ;
    buf_clk cell_4046 ( .C (clk), .D (signal_5588), .Q (signal_5589) ) ;
    buf_clk cell_4054 ( .C (clk), .D (signal_5596), .Q (signal_5597) ) ;
    buf_clk cell_4062 ( .C (clk), .D (signal_5604), .Q (signal_5605) ) ;
    buf_clk cell_4070 ( .C (clk), .D (signal_5612), .Q (signal_5613) ) ;
    buf_clk cell_4078 ( .C (clk), .D (signal_5620), .Q (signal_5621) ) ;
    buf_clk cell_4086 ( .C (clk), .D (signal_5628), .Q (signal_5629) ) ;
    buf_clk cell_4094 ( .C (clk), .D (signal_5636), .Q (signal_5637) ) ;
    buf_clk cell_4102 ( .C (clk), .D (signal_5644), .Q (signal_5645) ) ;
    buf_clk cell_4110 ( .C (clk), .D (signal_5652), .Q (signal_5653) ) ;
    buf_clk cell_4118 ( .C (clk), .D (signal_5660), .Q (signal_5661) ) ;
    buf_clk cell_4126 ( .C (clk), .D (signal_5668), .Q (signal_5669) ) ;
    buf_clk cell_4136 ( .C (clk), .D (signal_5678), .Q (signal_5679) ) ;
    buf_clk cell_4144 ( .C (clk), .D (signal_5686), .Q (signal_5687) ) ;
    buf_clk cell_4152 ( .C (clk), .D (signal_5694), .Q (signal_5695) ) ;
    buf_clk cell_4160 ( .C (clk), .D (signal_5702), .Q (signal_5703) ) ;
    buf_clk cell_4168 ( .C (clk), .D (signal_5710), .Q (signal_5711) ) ;
    buf_clk cell_4176 ( .C (clk), .D (signal_5718), .Q (signal_5719) ) ;
    buf_clk cell_4184 ( .C (clk), .D (signal_5726), .Q (signal_5727) ) ;
    buf_clk cell_4192 ( .C (clk), .D (signal_5734), .Q (signal_5735) ) ;
    buf_clk cell_4200 ( .C (clk), .D (signal_5742), .Q (signal_5743) ) ;
    buf_clk cell_4208 ( .C (clk), .D (signal_5750), .Q (signal_5751) ) ;
    buf_clk cell_4216 ( .C (clk), .D (signal_5758), .Q (signal_5759) ) ;
    buf_clk cell_4224 ( .C (clk), .D (signal_5766), .Q (signal_5767) ) ;
    buf_clk cell_4232 ( .C (clk), .D (signal_5774), .Q (signal_5775) ) ;
    buf_clk cell_4240 ( .C (clk), .D (signal_5782), .Q (signal_5783) ) ;
    buf_clk cell_4248 ( .C (clk), .D (signal_5790), .Q (signal_5791) ) ;
    buf_clk cell_4256 ( .C (clk), .D (signal_5798), .Q (signal_5799) ) ;
    buf_clk cell_4264 ( .C (clk), .D (signal_5806), .Q (signal_5807) ) ;
    buf_clk cell_4272 ( .C (clk), .D (signal_5814), .Q (signal_5815) ) ;
    buf_clk cell_4280 ( .C (clk), .D (signal_5822), .Q (signal_5823) ) ;
    buf_clk cell_4288 ( .C (clk), .D (signal_5830), .Q (signal_5831) ) ;
    buf_clk cell_4296 ( .C (clk), .D (signal_5838), .Q (signal_5839) ) ;
    buf_clk cell_4304 ( .C (clk), .D (signal_5846), .Q (signal_5847) ) ;
    buf_clk cell_4312 ( .C (clk), .D (signal_5854), .Q (signal_5855) ) ;
    buf_clk cell_4320 ( .C (clk), .D (signal_5862), .Q (signal_5863) ) ;
    buf_clk cell_4328 ( .C (clk), .D (signal_5870), .Q (signal_5871) ) ;
    buf_clk cell_4336 ( .C (clk), .D (signal_5878), .Q (signal_5879) ) ;
    buf_clk cell_4344 ( .C (clk), .D (signal_5886), .Q (signal_5887) ) ;
    buf_clk cell_4352 ( .C (clk), .D (signal_5894), .Q (signal_5895) ) ;
    buf_clk cell_4360 ( .C (clk), .D (signal_5902), .Q (signal_5903) ) ;
    buf_clk cell_4368 ( .C (clk), .D (signal_5910), .Q (signal_5911) ) ;
    buf_clk cell_4376 ( .C (clk), .D (signal_5918), .Q (signal_5919) ) ;
    buf_clk cell_4384 ( .C (clk), .D (signal_5926), .Q (signal_5927) ) ;
    buf_clk cell_4392 ( .C (clk), .D (signal_5934), .Q (signal_5935) ) ;
    buf_clk cell_4400 ( .C (clk), .D (signal_5942), .Q (signal_5943) ) ;
    buf_clk cell_4408 ( .C (clk), .D (signal_5950), .Q (signal_5951) ) ;
    buf_clk cell_4416 ( .C (clk), .D (signal_5958), .Q (signal_5959) ) ;
    buf_clk cell_4424 ( .C (clk), .D (signal_5966), .Q (signal_5967) ) ;
    buf_clk cell_4432 ( .C (clk), .D (signal_5974), .Q (signal_5975) ) ;
    buf_clk cell_4440 ( .C (clk), .D (signal_5982), .Q (signal_5983) ) ;
    buf_clk cell_4448 ( .C (clk), .D (signal_5990), .Q (signal_5991) ) ;
    buf_clk cell_4456 ( .C (clk), .D (signal_5998), .Q (signal_5999) ) ;
    buf_clk cell_4464 ( .C (clk), .D (signal_6006), .Q (signal_6007) ) ;
    buf_clk cell_4472 ( .C (clk), .D (signal_6014), .Q (signal_6015) ) ;
    buf_clk cell_4480 ( .C (clk), .D (signal_6022), .Q (signal_6023) ) ;
    buf_clk cell_4488 ( .C (clk), .D (signal_6030), .Q (signal_6031) ) ;
    buf_clk cell_4496 ( .C (clk), .D (signal_6038), .Q (signal_6039) ) ;
    buf_clk cell_4504 ( .C (clk), .D (signal_6046), .Q (signal_6047) ) ;
    buf_clk cell_4512 ( .C (clk), .D (signal_6054), .Q (signal_6055) ) ;
    buf_clk cell_4520 ( .C (clk), .D (signal_6062), .Q (signal_6063) ) ;
    buf_clk cell_4528 ( .C (clk), .D (signal_6070), .Q (signal_6071) ) ;
    buf_clk cell_4536 ( .C (clk), .D (signal_6078), .Q (signal_6079) ) ;
    buf_clk cell_4544 ( .C (clk), .D (signal_6086), .Q (signal_6087) ) ;
    buf_clk cell_4552 ( .C (clk), .D (signal_6094), .Q (signal_6095) ) ;
    buf_clk cell_4560 ( .C (clk), .D (signal_6102), .Q (signal_6103) ) ;
    buf_clk cell_4568 ( .C (clk), .D (signal_6110), .Q (signal_6111) ) ;
    buf_clk cell_4576 ( .C (clk), .D (signal_6118), .Q (signal_6119) ) ;
    buf_clk cell_4584 ( .C (clk), .D (signal_6126), .Q (signal_6127) ) ;
    buf_clk cell_4592 ( .C (clk), .D (signal_6134), .Q (signal_6135) ) ;
    buf_clk cell_4600 ( .C (clk), .D (signal_6142), .Q (signal_6143) ) ;
    buf_clk cell_4608 ( .C (clk), .D (signal_6150), .Q (signal_6151) ) ;
    buf_clk cell_4616 ( .C (clk), .D (signal_6158), .Q (signal_6159) ) ;
    buf_clk cell_4624 ( .C (clk), .D (signal_6166), .Q (signal_6167) ) ;
    buf_clk cell_4632 ( .C (clk), .D (signal_6174), .Q (signal_6175) ) ;
    buf_clk cell_4640 ( .C (clk), .D (signal_6182), .Q (signal_6183) ) ;
    buf_clk cell_4646 ( .C (clk), .D (signal_4508), .Q (signal_6189) ) ;
    buf_clk cell_4648 ( .C (clk), .D (signal_4512), .Q (signal_6191) ) ;
    buf_clk cell_4650 ( .C (clk), .D (signal_1553), .Q (signal_6193) ) ;
    buf_clk cell_4652 ( .C (clk), .D (signal_2095), .Q (signal_6195) ) ;
    buf_clk cell_4654 ( .C (clk), .D (signal_4528), .Q (signal_6197) ) ;
    buf_clk cell_4656 ( .C (clk), .D (signal_4532), .Q (signal_6199) ) ;
    buf_clk cell_4658 ( .C (clk), .D (signal_1535), .Q (signal_6201) ) ;
    buf_clk cell_4660 ( .C (clk), .D (signal_2076), .Q (signal_6203) ) ;
    buf_clk cell_4662 ( .C (clk), .D (signal_4556), .Q (signal_6205) ) ;
    buf_clk cell_4664 ( .C (clk), .D (signal_4560), .Q (signal_6207) ) ;
    buf_clk cell_4666 ( .C (clk), .D (signal_1517), .Q (signal_6209) ) ;
    buf_clk cell_4668 ( .C (clk), .D (signal_2050), .Q (signal_6211) ) ;
    buf_clk cell_4670 ( .C (clk), .D (signal_4536), .Q (signal_6213) ) ;
    buf_clk cell_4672 ( .C (clk), .D (signal_4540), .Q (signal_6215) ) ;
    buf_clk cell_4674 ( .C (clk), .D (signal_1532), .Q (signal_6217) ) ;
    buf_clk cell_4676 ( .C (clk), .D (signal_2071), .Q (signal_6219) ) ;
    buf_clk cell_4678 ( .C (clk), .D (signal_4520), .Q (signal_6221) ) ;
    buf_clk cell_4680 ( .C (clk), .D (signal_4524), .Q (signal_6223) ) ;
    buf_clk cell_4682 ( .C (clk), .D (signal_1545), .Q (signal_6225) ) ;
    buf_clk cell_4684 ( .C (clk), .D (signal_2086), .Q (signal_6227) ) ;
    buf_clk cell_4686 ( .C (clk), .D (signal_4572), .Q (signal_6229) ) ;
    buf_clk cell_4688 ( .C (clk), .D (signal_4576), .Q (signal_6231) ) ;
    buf_clk cell_4690 ( .C (clk), .D (signal_1551), .Q (signal_6233) ) ;
    buf_clk cell_4692 ( .C (clk), .D (signal_2092), .Q (signal_6235) ) ;
    buf_clk cell_4694 ( .C (clk), .D (signal_1525), .Q (signal_6237) ) ;
    buf_clk cell_4696 ( .C (clk), .D (signal_2061), .Q (signal_6239) ) ;
    buf_clk cell_4698 ( .C (clk), .D (signal_1534), .Q (signal_6241) ) ;
    buf_clk cell_4700 ( .C (clk), .D (signal_2074), .Q (signal_6243) ) ;
    buf_clk cell_4702 ( .C (clk), .D (signal_1527), .Q (signal_6245) ) ;
    buf_clk cell_4704 ( .C (clk), .D (signal_2063), .Q (signal_6247) ) ;
    buf_clk cell_4706 ( .C (clk), .D (signal_4564), .Q (signal_6249) ) ;
    buf_clk cell_4708 ( .C (clk), .D (signal_4568), .Q (signal_6251) ) ;
    buf_clk cell_4710 ( .C (clk), .D (signal_1499), .Q (signal_6253) ) ;
    buf_clk cell_4712 ( .C (clk), .D (signal_2025), .Q (signal_6255) ) ;
    buf_clk cell_4714 ( .C (clk), .D (signal_4500), .Q (signal_6257) ) ;
    buf_clk cell_4716 ( .C (clk), .D (signal_4504), .Q (signal_6259) ) ;
    buf_clk cell_4718 ( .C (clk), .D (signal_1539), .Q (signal_6261) ) ;
    buf_clk cell_4720 ( .C (clk), .D (signal_2080), .Q (signal_6263) ) ;
    buf_clk cell_4722 ( .C (clk), .D (signal_1522), .Q (signal_6265) ) ;
    buf_clk cell_4724 ( .C (clk), .D (signal_2057), .Q (signal_6267) ) ;
    buf_clk cell_4726 ( .C (clk), .D (signal_1512), .Q (signal_6269) ) ;
    buf_clk cell_4728 ( .C (clk), .D (signal_2044), .Q (signal_6271) ) ;
    buf_clk cell_4730 ( .C (clk), .D (signal_1533), .Q (signal_6273) ) ;
    buf_clk cell_4732 ( .C (clk), .D (signal_2073), .Q (signal_6275) ) ;
    buf_clk cell_4734 ( .C (clk), .D (signal_4464), .Q (signal_6277) ) ;
    buf_clk cell_4736 ( .C (clk), .D (signal_4468), .Q (signal_6279) ) ;
    buf_clk cell_4738 ( .C (clk), .D (signal_1518), .Q (signal_6281) ) ;
    buf_clk cell_4740 ( .C (clk), .D (signal_2051), .Q (signal_6283) ) ;
    buf_clk cell_4742 ( .C (clk), .D (signal_1528), .Q (signal_6285) ) ;
    buf_clk cell_4744 ( .C (clk), .D (signal_2065), .Q (signal_6287) ) ;
    buf_clk cell_4746 ( .C (clk), .D (signal_1513), .Q (signal_6289) ) ;
    buf_clk cell_4748 ( .C (clk), .D (signal_2046), .Q (signal_6291) ) ;
    buf_clk cell_4750 ( .C (clk), .D (signal_4644), .Q (signal_6293) ) ;
    buf_clk cell_4752 ( .C (clk), .D (signal_4648), .Q (signal_6295) ) ;
    buf_clk cell_4754 ( .C (clk), .D (signal_1523), .Q (signal_6297) ) ;
    buf_clk cell_4756 ( .C (clk), .D (signal_2058), .Q (signal_6299) ) ;
    buf_clk cell_4758 ( .C (clk), .D (signal_1538), .Q (signal_6301) ) ;
    buf_clk cell_4760 ( .C (clk), .D (signal_2079), .Q (signal_6303) ) ;
    buf_clk cell_4762 ( .C (clk), .D (signal_4580), .Q (signal_6305) ) ;
    buf_clk cell_4764 ( .C (clk), .D (signal_4584), .Q (signal_6307) ) ;
    buf_clk cell_4766 ( .C (clk), .D (signal_1530), .Q (signal_6309) ) ;
    buf_clk cell_4768 ( .C (clk), .D (signal_2068), .Q (signal_6311) ) ;
    buf_clk cell_4770 ( .C (clk), .D (signal_4548), .Q (signal_6313) ) ;
    buf_clk cell_4772 ( .C (clk), .D (signal_4552), .Q (signal_6315) ) ;
    buf_clk cell_4774 ( .C (clk), .D (signal_1519), .Q (signal_6317) ) ;
    buf_clk cell_4776 ( .C (clk), .D (signal_2053), .Q (signal_6319) ) ;
    buf_clk cell_4778 ( .C (clk), .D (signal_1556), .Q (signal_6321) ) ;
    buf_clk cell_4780 ( .C (clk), .D (signal_2099), .Q (signal_6323) ) ;
    buf_clk cell_4782 ( .C (clk), .D (signal_4596), .Q (signal_6325) ) ;
    buf_clk cell_4784 ( .C (clk), .D (signal_4600), .Q (signal_6327) ) ;
    buf_clk cell_4786 ( .C (clk), .D (signal_1563), .Q (signal_6329) ) ;
    buf_clk cell_4788 ( .C (clk), .D (signal_2107), .Q (signal_6331) ) ;
    buf_clk cell_4790 ( .C (clk), .D (signal_1564), .Q (signal_6333) ) ;
    buf_clk cell_4792 ( .C (clk), .D (signal_2108), .Q (signal_6335) ) ;
    buf_clk cell_4794 ( .C (clk), .D (signal_4608), .Q (signal_6337) ) ;
    buf_clk cell_4796 ( .C (clk), .D (signal_4612), .Q (signal_6339) ) ;
    buf_clk cell_4798 ( .C (clk), .D (signal_1569), .Q (signal_6341) ) ;
    buf_clk cell_4800 ( .C (clk), .D (signal_2114), .Q (signal_6343) ) ;
    buf_clk cell_4802 ( .C (clk), .D (signal_1570), .Q (signal_6345) ) ;
    buf_clk cell_4804 ( .C (clk), .D (signal_2115), .Q (signal_6347) ) ;
    buf_clk cell_4806 ( .C (clk), .D (signal_4620), .Q (signal_6349) ) ;
    buf_clk cell_4808 ( .C (clk), .D (signal_4624), .Q (signal_6351) ) ;
    buf_clk cell_4810 ( .C (clk), .D (signal_1576), .Q (signal_6353) ) ;
    buf_clk cell_4812 ( .C (clk), .D (signal_2122), .Q (signal_6355) ) ;
    buf_clk cell_4814 ( .C (clk), .D (signal_1577), .Q (signal_6357) ) ;
    buf_clk cell_4816 ( .C (clk), .D (signal_2123), .Q (signal_6359) ) ;
    buf_clk cell_4818 ( .C (clk), .D (signal_4632), .Q (signal_6361) ) ;
    buf_clk cell_4820 ( .C (clk), .D (signal_4636), .Q (signal_6363) ) ;
    buf_clk cell_4822 ( .C (clk), .D (signal_1582), .Q (signal_6365) ) ;
    buf_clk cell_4824 ( .C (clk), .D (signal_2129), .Q (signal_6367) ) ;
    buf_clk cell_4826 ( .C (clk), .D (signal_1583), .Q (signal_6369) ) ;
    buf_clk cell_4828 ( .C (clk), .D (signal_2130), .Q (signal_6371) ) ;
    buf_clk cell_4830 ( .C (clk), .D (signal_1588), .Q (signal_6373) ) ;
    buf_clk cell_4832 ( .C (clk), .D (signal_2136), .Q (signal_6375) ) ;
    buf_clk cell_4834 ( .C (clk), .D (signal_1496), .Q (signal_6377) ) ;
    buf_clk cell_4836 ( .C (clk), .D (signal_2020), .Q (signal_6379) ) ;
    buf_clk cell_4842 ( .C (clk), .D (signal_6384), .Q (signal_6385) ) ;
    buf_clk cell_4850 ( .C (clk), .D (signal_6392), .Q (signal_6393) ) ;
    buf_clk cell_4858 ( .C (clk), .D (signal_6400), .Q (signal_6401) ) ;
    buf_clk cell_4866 ( .C (clk), .D (signal_6408), .Q (signal_6409) ) ;

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_89 ( .a ({signal_3304, signal_3298}), .b ({signal_2236, signal_1302}), .c ({signal_2270, signal_255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_91 ( .a ({signal_3316, signal_3310}), .b ({signal_2234, signal_1264}), .c ({signal_2271, signal_257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_93 ( .a ({signal_3328, signal_3322}), .b ({signal_2218, signal_1248}), .c ({signal_2272, signal_201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_95 ( .a ({signal_3340, signal_3334}), .b ({signal_2207, signal_1250}), .c ({signal_2273, signal_203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_97 ( .a ({signal_3352, signal_3346}), .b ({signal_2209, signal_1266}), .c ({signal_2274, signal_259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_98 ( .a ({signal_3364, signal_3358}), .b ({signal_2227, signal_1276}), .c ({signal_2275, signal_205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_100 ( .a ({signal_3376, signal_3370}), .b ({signal_2208, signal_1278}), .c ({signal_2276, signal_207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_102 ( .a ({signal_3388, signal_3382}), .b ({signal_2231, signal_1304}), .c ({signal_2277, signal_209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_104 ( .a ({signal_3400, signal_3394}), .b ({signal_2194, signal_1306}), .c ({signal_2278, signal_211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_106 ( .a ({signal_3412, signal_3406}), .b ({signal_2206, signal_1284}), .c ({signal_2279, signal_213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_109 ( .a ({signal_3424, signal_3418}), .b ({signal_2190, signal_1286}), .c ({signal_2280, signal_215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_111 ( .a ({signal_3436, signal_3430}), .b ({signal_2203, signal_1268}), .c ({signal_2281, signal_217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_113 ( .a ({signal_3448, signal_3442}), .b ({signal_2223, signal_1270}), .c ({signal_2282, signal_219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_115 ( .a ({signal_3460, signal_3454}), .b ({signal_2192, signal_1256}), .c ({signal_2283, signal_221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_117 ( .a ({signal_3472, signal_3466}), .b ({signal_2199, signal_1258}), .c ({signal_2284, signal_223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_119 ( .a ({signal_3484, signal_3478}), .b ({signal_2225, signal_1260}), .c ({signal_2285, signal_261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_120 ( .a ({signal_3496, signal_3490}), .b ({signal_2212, signal_1292}), .c ({signal_2286, signal_225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_122 ( .a ({signal_3508, signal_3502}), .b ({signal_2238, signal_1294}), .c ({signal_2287, signal_227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_124 ( .a ({signal_3520, signal_3514}), .b ({signal_2220, signal_1296}), .c ({signal_2288, signal_229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_126 ( .a ({signal_3532, signal_3526}), .b ({signal_2235, signal_1298}), .c ({signal_2289, signal_231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_128 ( .a ({signal_3544, signal_3538}), .b ({signal_2240, signal_1308}), .c ({signal_2290, signal_233}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_131 ( .a ({signal_3556, signal_3550}), .b ({signal_2243, signal_1310}), .c ({signal_2291, signal_235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_133 ( .a ({signal_3568, signal_3562}), .b ({signal_2246, signal_1280}), .c ({signal_2292, signal_237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_135 ( .a ({signal_3580, signal_3574}), .b ({signal_2248, signal_1282}), .c ({signal_2293, signal_239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_137 ( .a ({signal_3592, signal_3586}), .b ({signal_2251, signal_1252}), .c ({signal_2294, signal_241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_139 ( .a ({signal_3604, signal_3598}), .b ({signal_2253, signal_1254}), .c ({signal_2295, signal_243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_141 ( .a ({signal_3616, signal_3610}), .b ({signal_2255, signal_1262}), .c ({signal_2296, signal_263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_142 ( .a ({signal_3628, signal_3622}), .b ({signal_2257, signal_1272}), .c ({signal_2297, signal_245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_144 ( .a ({signal_3640, signal_3634}), .b ({signal_2259, signal_1274}), .c ({signal_2298, signal_247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_146 ( .a ({signal_3652, signal_3646}), .b ({signal_2262, signal_1288}), .c ({signal_2299, signal_249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_148 ( .a ({signal_3664, signal_3658}), .b ({signal_2264, signal_1290}), .c ({signal_2300, signal_251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_150 ( .a ({signal_3676, signal_3670}), .b ({signal_2267, signal_1300}), .c ({signal_2301, signal_253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .a ({signal_3688, signal_3682}), .b ({signal_2236, signal_1302}), .c ({signal_2302, signal_1238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .a ({signal_3700, signal_3694}), .b ({signal_2234, signal_1264}), .c ({signal_2303, signal_1240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_221 ( .a ({signal_3712, signal_3706}), .b ({signal_2218, signal_1248}), .c ({signal_2304, signal_1184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_223 ( .a ({signal_3724, signal_3718}), .b ({signal_2207, signal_1250}), .c ({signal_2305, signal_1186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_225 ( .a ({signal_3736, signal_3730}), .b ({signal_2209, signal_1266}), .c ({signal_2306, signal_1242}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_226 ( .a ({signal_3748, signal_3742}), .b ({signal_2227, signal_1276}), .c ({signal_2307, signal_1188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .a ({signal_3760, signal_3754}), .b ({signal_2208, signal_1278}), .c ({signal_2308, signal_1190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .a ({signal_3772, signal_3766}), .b ({signal_2231, signal_1304}), .c ({signal_2309, signal_1192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_232 ( .a ({signal_3784, signal_3778}), .b ({signal_2194, signal_1306}), .c ({signal_2310, signal_1194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_234 ( .a ({signal_3796, signal_3790}), .b ({signal_2206, signal_1284}), .c ({signal_2311, signal_1196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({signal_3808, signal_3802}), .b ({signal_2190, signal_1286}), .c ({signal_2312, signal_1198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({signal_3820, signal_3814}), .b ({signal_2203, signal_1268}), .c ({signal_2313, signal_1200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({signal_3832, signal_3826}), .b ({signal_2223, signal_1270}), .c ({signal_2314, signal_1202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({signal_3844, signal_3838}), .b ({signal_2192, signal_1256}), .c ({signal_2315, signal_1204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({signal_3856, signal_3850}), .b ({signal_2199, signal_1258}), .c ({signal_2316, signal_1206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({signal_3868, signal_3862}), .b ({signal_2225, signal_1260}), .c ({signal_2317, signal_1244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({signal_3880, signal_3874}), .b ({signal_2212, signal_1292}), .c ({signal_2318, signal_1208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({signal_3892, signal_3886}), .b ({signal_2238, signal_1294}), .c ({signal_2319, signal_1210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({signal_3904, signal_3898}), .b ({signal_2220, signal_1296}), .c ({signal_2320, signal_1212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({signal_3916, signal_3910}), .b ({signal_2235, signal_1298}), .c ({signal_2321, signal_1214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({signal_3928, signal_3922}), .b ({signal_2240, signal_1308}), .c ({signal_2322, signal_1216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .a ({signal_3940, signal_3934}), .b ({signal_2243, signal_1310}), .c ({signal_2323, signal_1218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .a ({signal_3952, signal_3946}), .b ({signal_2246, signal_1280}), .c ({signal_2324, signal_1220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({signal_3964, signal_3958}), .b ({signal_2248, signal_1282}), .c ({signal_2325, signal_1222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .a ({signal_3976, signal_3970}), .b ({signal_2251, signal_1252}), .c ({signal_2326, signal_1224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .a ({signal_3988, signal_3982}), .b ({signal_2253, signal_1254}), .c ({signal_2327, signal_1226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .a ({signal_4000, signal_3994}), .b ({signal_2255, signal_1262}), .c ({signal_2328, signal_1246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({signal_4012, signal_4006}), .b ({signal_2257, signal_1272}), .c ({signal_2329, signal_1228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .a ({signal_4024, signal_4018}), .b ({signal_2259, signal_1274}), .c ({signal_2330, signal_1230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({signal_4036, signal_4030}), .b ({signal_2262, signal_1288}), .c ({signal_2331, signal_1232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({signal_4048, signal_4042}), .b ({signal_2264, signal_1290}), .c ({signal_2332, signal_1234}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({signal_4060, signal_4054}), .b ({signal_2267, signal_1300}), .c ({signal_2333, signal_1236}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .a ({signal_3688, signal_3682}), .b ({signal_2508, signal_1110}), .c ({signal_2518, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .a ({signal_3700, signal_3694}), .b ({signal_2509, signal_1064}), .c ({signal_2519, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_286 ( .a ({signal_3712, signal_3706}), .b ({signal_2484, signal_1056}), .c ({signal_2520, signal_992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .a ({signal_3724, signal_3718}), .b ({signal_2485, signal_1058}), .c ({signal_2521, signal_994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_291 ( .a ({signal_3736, signal_3730}), .b ({signal_2510, signal_1066}), .c ({signal_2522, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_292 ( .a ({signal_3748, signal_3742}), .b ({signal_2486, signal_1096}), .c ({signal_2523, signal_996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .a ({signal_3760, signal_3754}), .b ({signal_2478, signal_1098}), .c ({signal_2524, signal_998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_297 ( .a ({signal_3772, signal_3766}), .b ({signal_2479, signal_1076}), .c ({signal_2525, signal_1000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_299 ( .a ({signal_3784, signal_3778}), .b ({signal_2480, signal_1078}), .c ({signal_2526, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_302 ( .a ({signal_3796, signal_3790}), .b ({signal_2481, signal_1116}), .c ({signal_2527, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_306 ( .a ({signal_3808, signal_3802}), .b ({signal_2483, signal_1118}), .c ({signal_2528, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_309 ( .a ({signal_3820, signal_3814}), .b ({signal_2494, signal_1112}), .c ({signal_2529, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_311 ( .a ({signal_3832, signal_3826}), .b ({signal_2495, signal_1114}), .c ({signal_2530, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_314 ( .a ({signal_3844, signal_3838}), .b ({signal_2496, signal_1072}), .c ({signal_2531, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_316 ( .a ({signal_3856, signal_3850}), .b ({signal_2488, signal_1074}), .c ({signal_2532, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_319 ( .a ({signal_3868, signal_3862}), .b ({signal_2511, signal_1088}), .c ({signal_2533, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_320 ( .a ({signal_3880, signal_3874}), .b ({signal_2489, signal_1100}), .c ({signal_2534, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_322 ( .a ({signal_3892, signal_3886}), .b ({signal_2490, signal_1102}), .c ({signal_2535, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_325 ( .a ({signal_3904, signal_3898}), .b ({signal_2491, signal_1060}), .c ({signal_2536, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_327 ( .a ({signal_3916, signal_3910}), .b ({signal_2493, signal_1062}), .c ({signal_2537, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_330 ( .a ({signal_3928, signal_3922}), .b ({signal_2504, signal_1092}), .c ({signal_2538, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_333 ( .a ({signal_3940, signal_3934}), .b ({signal_2505, signal_1094}), .c ({signal_2539, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_336 ( .a ({signal_3952, signal_3946}), .b ({signal_2506, signal_1068}), .c ({signal_2540, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_338 ( .a ({signal_3964, signal_3958}), .b ({signal_2498, signal_1070}), .c ({signal_2541, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_341 ( .a ({signal_3976, signal_3970}), .b ({signal_2499, signal_1104}), .c ({signal_2542, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_343 ( .a ({signal_3988, signal_3982}), .b ({signal_2500, signal_1106}), .c ({signal_2543, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_346 ( .a ({signal_4000, signal_3994}), .b ({signal_2513, signal_1090}), .c ({signal_2544, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_347 ( .a ({signal_4012, signal_4006}), .b ({signal_2501, signal_1080}), .c ({signal_2545, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_349 ( .a ({signal_4024, signal_4018}), .b ({signal_2503, signal_1082}), .c ({signal_2546, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_352 ( .a ({signal_4036, signal_4030}), .b ({signal_2514, signal_1084}), .c ({signal_2547, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_354 ( .a ({signal_4048, signal_4042}), .b ({signal_2515, signal_1086}), .c ({signal_2548, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_357 ( .a ({signal_4060, signal_4054}), .b ({signal_2516, signal_1108}), .c ({signal_2549, signal_1044}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_538 ( .s (signal_4066), .b ({signal_2586, signal_1438}), .a ({signal_4078, signal_4072}), .c ({signal_2632, signal_462}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_544 ( .s (signal_4066), .b ({signal_2587, signal_1436}), .a ({signal_4090, signal_4084}), .c ({signal_2633, signal_466}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_550 ( .s (signal_4066), .b ({signal_2588, signal_1434}), .a ({signal_4102, signal_4096}), .c ({signal_2634, signal_470}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_556 ( .s (signal_4066), .b ({signal_2589, signal_1432}), .a ({signal_4114, signal_4108}), .c ({signal_2635, signal_474}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_562 ( .s (signal_4066), .b ({signal_2590, signal_1430}), .a ({signal_4126, signal_4120}), .c ({signal_2636, signal_478}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_568 ( .s (signal_4066), .b ({signal_2591, signal_1428}), .a ({signal_4138, signal_4132}), .c ({signal_2637, signal_482}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_574 ( .s (signal_4066), .b ({signal_2592, signal_1426}), .a ({signal_4150, signal_4144}), .c ({signal_2638, signal_486}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_580 ( .s (signal_4066), .b ({signal_2593, signal_1424}), .a ({signal_4162, signal_4156}), .c ({signal_2639, signal_490}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_586 ( .s (signal_4066), .b ({signal_2594, signal_1422}), .a ({signal_4174, signal_4168}), .c ({signal_2640, signal_494}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_592 ( .s (signal_4066), .b ({signal_2595, signal_1420}), .a ({signal_4186, signal_4180}), .c ({signal_2641, signal_498}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_598 ( .s (signal_4066), .b ({signal_2596, signal_1418}), .a ({signal_4198, signal_4192}), .c ({signal_2642, signal_502}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_604 ( .s (signal_4066), .b ({signal_2597, signal_1416}), .a ({signal_4210, signal_4204}), .c ({signal_2643, signal_506}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_610 ( .s (signal_4066), .b ({signal_2598, signal_1414}), .a ({signal_4222, signal_4216}), .c ({signal_2644, signal_510}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_616 ( .s (signal_4066), .b ({signal_2599, signal_1412}), .a ({signal_4234, signal_4228}), .c ({signal_2645, signal_514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_622 ( .s (signal_4066), .b ({signal_2600, signal_1410}), .a ({signal_4246, signal_4240}), .c ({signal_2646, signal_518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_628 ( .s (signal_4066), .b ({signal_2601, signal_1408}), .a ({signal_4258, signal_4252}), .c ({signal_2647, signal_522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_634 ( .s (signal_4066), .b ({signal_2602, signal_1406}), .a ({signal_4270, signal_4264}), .c ({signal_2648, signal_526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_640 ( .s (signal_4066), .b ({signal_2603, signal_1404}), .a ({signal_4282, signal_4276}), .c ({signal_2649, signal_530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_646 ( .s (signal_4066), .b ({signal_2604, signal_1402}), .a ({signal_4294, signal_4288}), .c ({signal_2650, signal_534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_652 ( .s (signal_4066), .b ({signal_2605, signal_1400}), .a ({signal_4306, signal_4300}), .c ({signal_2651, signal_538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_658 ( .s (signal_4066), .b ({signal_2606, signal_1398}), .a ({signal_4318, signal_4312}), .c ({signal_2652, signal_542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_664 ( .s (signal_4066), .b ({signal_2607, signal_1396}), .a ({signal_4330, signal_4324}), .c ({signal_2653, signal_546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_670 ( .s (signal_4066), .b ({signal_2608, signal_1394}), .a ({signal_4342, signal_4336}), .c ({signal_2654, signal_550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_676 ( .s (signal_4066), .b ({signal_2609, signal_1392}), .a ({signal_4354, signal_4348}), .c ({signal_2655, signal_554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_682 ( .s (signal_4066), .b ({signal_2610, signal_1390}), .a ({signal_4366, signal_4360}), .c ({signal_2656, signal_558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_688 ( .s (signal_4066), .b ({signal_2611, signal_1388}), .a ({signal_4378, signal_4372}), .c ({signal_2657, signal_562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_694 ( .s (signal_4066), .b ({signal_2612, signal_1386}), .a ({signal_4390, signal_4384}), .c ({signal_2658, signal_566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_700 ( .s (signal_4066), .b ({signal_2613, signal_1384}), .a ({signal_4402, signal_4396}), .c ({signal_2659, signal_570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_706 ( .s (signal_4066), .b ({signal_2614, signal_1382}), .a ({signal_4414, signal_4408}), .c ({signal_2660, signal_574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_712 ( .s (signal_4066), .b ({signal_2615, signal_1380}), .a ({signal_4426, signal_4420}), .c ({signal_2661, signal_578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_718 ( .s (signal_4066), .b ({signal_2616, signal_1378}), .a ({signal_4438, signal_4432}), .c ({signal_2662, signal_582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_724 ( .s (signal_4066), .b ({signal_2617, signal_1376}), .a ({signal_4450, signal_4444}), .c ({signal_2663, signal_586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1032 ( .s (signal_4456), .b ({signal_2243, signal_1310}), .a ({signal_2328, signal_1246}), .c ({signal_2414, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1034 ( .s (signal_4456), .b ({signal_2240, signal_1308}), .a ({signal_2317, signal_1244}), .c ({signal_2415, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1036 ( .s (signal_4456), .b ({signal_2194, signal_1306}), .a ({signal_2306, signal_1242}), .c ({signal_2416, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1038 ( .s (signal_4456), .b ({signal_2231, signal_1304}), .a ({signal_2303, signal_1240}), .c ({signal_2417, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1040 ( .s (signal_4456), .b ({signal_2236, signal_1302}), .a ({signal_2302, signal_1238}), .c ({signal_2418, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1042 ( .s (signal_4456), .b ({signal_2267, signal_1300}), .a ({signal_2333, signal_1236}), .c ({signal_2419, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1044 ( .s (signal_4456), .b ({signal_2235, signal_1298}), .a ({signal_2332, signal_1234}), .c ({signal_2420, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1046 ( .s (signal_4456), .b ({signal_2220, signal_1296}), .a ({signal_2331, signal_1232}), .c ({signal_2421, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1048 ( .s (signal_4456), .b ({signal_2238, signal_1294}), .a ({signal_2330, signal_1230}), .c ({signal_2422, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1050 ( .s (signal_4456), .b ({signal_2212, signal_1292}), .a ({signal_2329, signal_1228}), .c ({signal_2423, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1052 ( .s (signal_4456), .b ({signal_2264, signal_1290}), .a ({signal_2327, signal_1226}), .c ({signal_2424, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1054 ( .s (signal_4456), .b ({signal_2262, signal_1288}), .a ({signal_2326, signal_1224}), .c ({signal_2425, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1056 ( .s (signal_4456), .b ({signal_2190, signal_1286}), .a ({signal_2325, signal_1222}), .c ({signal_2426, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1058 ( .s (signal_4456), .b ({signal_2206, signal_1284}), .a ({signal_2324, signal_1220}), .c ({signal_2427, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1060 ( .s (signal_4456), .b ({signal_2248, signal_1282}), .a ({signal_2323, signal_1218}), .c ({signal_2428, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1062 ( .s (signal_4456), .b ({signal_2246, signal_1280}), .a ({signal_2322, signal_1216}), .c ({signal_2429, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1064 ( .s (signal_4456), .b ({signal_2208, signal_1278}), .a ({signal_2321, signal_1214}), .c ({signal_2430, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1066 ( .s (signal_4456), .b ({signal_2227, signal_1276}), .a ({signal_2320, signal_1212}), .c ({signal_2431, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1068 ( .s (signal_4456), .b ({signal_2259, signal_1274}), .a ({signal_2319, signal_1210}), .c ({signal_2432, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1070 ( .s (signal_4456), .b ({signal_2257, signal_1272}), .a ({signal_2318, signal_1208}), .c ({signal_2433, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1072 ( .s (signal_4456), .b ({signal_2223, signal_1270}), .a ({signal_2316, signal_1206}), .c ({signal_2434, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1074 ( .s (signal_4456), .b ({signal_2203, signal_1268}), .a ({signal_2315, signal_1204}), .c ({signal_2435, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1076 ( .s (signal_4456), .b ({signal_2209, signal_1266}), .a ({signal_2314, signal_1202}), .c ({signal_2436, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1078 ( .s (signal_4456), .b ({signal_2234, signal_1264}), .a ({signal_2313, signal_1200}), .c ({signal_2437, signal_1136}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1080 ( .s (signal_4456), .b ({signal_2255, signal_1262}), .a ({signal_2312, signal_1198}), .c ({signal_2438, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1082 ( .s (signal_4456), .b ({signal_2225, signal_1260}), .a ({signal_2311, signal_1196}), .c ({signal_2439, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1084 ( .s (signal_4456), .b ({signal_2199, signal_1258}), .a ({signal_2310, signal_1194}), .c ({signal_2440, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1086 ( .s (signal_4456), .b ({signal_2192, signal_1256}), .a ({signal_2309, signal_1192}), .c ({signal_2441, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1088 ( .s (signal_4456), .b ({signal_2253, signal_1254}), .a ({signal_2308, signal_1190}), .c ({signal_2442, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1090 ( .s (signal_4456), .b ({signal_2251, signal_1252}), .a ({signal_2307, signal_1188}), .c ({signal_2443, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1092 ( .s (signal_4456), .b ({signal_2207, signal_1250}), .a ({signal_2305, signal_1186}), .c ({signal_2444, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1094 ( .s (signal_4456), .b ({signal_2218, signal_1248}), .a ({signal_2304, signal_1184}), .c ({signal_2445, signal_1120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1095 ( .a ({signal_2444, signal_1122}), .b ({signal_2464, signal_828}), .c ({signal_2478, signal_1098}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1097 ( .a ({signal_2439, signal_1132}), .b ({signal_2462, signal_830}), .c ({signal_2479, signal_1076}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1099 ( .a ({signal_2438, signal_1134}), .b ({signal_2463, signal_832}), .c ({signal_2480, signal_1078}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1101 ( .a ({signal_2441, signal_1128}), .b ({signal_2462, signal_830}), .c ({signal_2481, signal_1116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1102 ( .a ({signal_2445, signal_1120}), .b ({signal_2443, signal_1124}), .c ({signal_2462, signal_830}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1105 ( .a ({signal_2440, signal_1130}), .b ({signal_2463, signal_832}), .c ({signal_2483, signal_1118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1106 ( .a ({signal_2442, signal_1126}), .b ({signal_2444, signal_1122}), .c ({signal_2463, signal_832}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1107 ( .a ({signal_2443, signal_1124}), .b ({signal_2465, signal_834}), .c ({signal_2484, signal_1056}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1109 ( .a ({signal_2442, signal_1126}), .b ({signal_2464, signal_828}), .c ({signal_2485, signal_1058}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1110 ( .a ({signal_2438, signal_1134}), .b ({signal_2440, signal_1130}), .c ({signal_2464, signal_828}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1113 ( .a ({signal_2445, signal_1120}), .b ({signal_2465, signal_834}), .c ({signal_2486, signal_1096}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1114 ( .a ({signal_2439, signal_1132}), .b ({signal_2441, signal_1128}), .c ({signal_2465, signal_834}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1119 ( .a ({signal_2436, signal_1138}), .b ({signal_2468, signal_836}), .c ({signal_2488, signal_1074}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1121 ( .a ({signal_2431, signal_1148}), .b ({signal_2466, signal_838}), .c ({signal_2489, signal_1100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1123 ( .a ({signal_2430, signal_1150}), .b ({signal_2467, signal_840}), .c ({signal_2490, signal_1102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1125 ( .a ({signal_2433, signal_1144}), .b ({signal_2466, signal_838}), .c ({signal_2491, signal_1060}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1126 ( .a ({signal_2437, signal_1136}), .b ({signal_2435, signal_1140}), .c ({signal_2466, signal_838}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1129 ( .a ({signal_2432, signal_1146}), .b ({signal_2467, signal_840}), .c ({signal_2493, signal_1062}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1130 ( .a ({signal_2434, signal_1142}), .b ({signal_2436, signal_1138}), .c ({signal_2467, signal_840}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1131 ( .a ({signal_2435, signal_1140}), .b ({signal_2469, signal_842}), .c ({signal_2494, signal_1112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1133 ( .a ({signal_2434, signal_1142}), .b ({signal_2468, signal_836}), .c ({signal_2495, signal_1114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1134 ( .a ({signal_2430, signal_1150}), .b ({signal_2432, signal_1146}), .c ({signal_2468, signal_836}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1137 ( .a ({signal_2437, signal_1136}), .b ({signal_2469, signal_842}), .c ({signal_2496, signal_1072}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1138 ( .a ({signal_2431, signal_1148}), .b ({signal_2433, signal_1144}), .c ({signal_2469, signal_842}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1143 ( .a ({signal_2428, signal_1154}), .b ({signal_2472, signal_844}), .c ({signal_2498, signal_1070}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1145 ( .a ({signal_2423, signal_1164}), .b ({signal_2470, signal_846}), .c ({signal_2499, signal_1104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1147 ( .a ({signal_2422, signal_1166}), .b ({signal_2471, signal_848}), .c ({signal_2500, signal_1106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1149 ( .a ({signal_2425, signal_1160}), .b ({signal_2470, signal_846}), .c ({signal_2501, signal_1080}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1150 ( .a ({signal_2429, signal_1152}), .b ({signal_2427, signal_1156}), .c ({signal_2470, signal_846}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1153 ( .a ({signal_2424, signal_1162}), .b ({signal_2471, signal_848}), .c ({signal_2503, signal_1082}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1154 ( .a ({signal_2426, signal_1158}), .b ({signal_2428, signal_1154}), .c ({signal_2471, signal_848}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1155 ( .a ({signal_2427, signal_1156}), .b ({signal_2473, signal_850}), .c ({signal_2504, signal_1092}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1157 ( .a ({signal_2426, signal_1158}), .b ({signal_2472, signal_844}), .c ({signal_2505, signal_1094}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1158 ( .a ({signal_2422, signal_1166}), .b ({signal_2424, signal_1162}), .c ({signal_2472, signal_844}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1161 ( .a ({signal_2429, signal_1152}), .b ({signal_2473, signal_850}), .c ({signal_2506, signal_1068}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1162 ( .a ({signal_2423, signal_1164}), .b ({signal_2425, signal_1160}), .c ({signal_2473, signal_850}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1167 ( .a ({signal_2420, signal_1170}), .b ({signal_2476, signal_852}), .c ({signal_2508, signal_1110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1169 ( .a ({signal_2415, signal_1180}), .b ({signal_2474, signal_854}), .c ({signal_2509, signal_1064}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1171 ( .a ({signal_2414, signal_1182}), .b ({signal_2475, signal_856}), .c ({signal_2510, signal_1066}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1173 ( .a ({signal_2417, signal_1176}), .b ({signal_2474, signal_854}), .c ({signal_2511, signal_1088}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1174 ( .a ({signal_2421, signal_1168}), .b ({signal_2419, signal_1172}), .c ({signal_2474, signal_854}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1177 ( .a ({signal_2416, signal_1178}), .b ({signal_2475, signal_856}), .c ({signal_2513, signal_1090}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1178 ( .a ({signal_2418, signal_1174}), .b ({signal_2420, signal_1170}), .c ({signal_2475, signal_856}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1179 ( .a ({signal_2419, signal_1172}), .b ({signal_2477, signal_858}), .c ({signal_2514, signal_1084}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1181 ( .a ({signal_2418, signal_1174}), .b ({signal_2476, signal_852}), .c ({signal_2515, signal_1086}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1182 ( .a ({signal_2414, signal_1182}), .b ({signal_2416, signal_1178}), .c ({signal_2476, signal_852}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1185 ( .a ({signal_2421, signal_1168}), .b ({signal_2477, signal_858}), .c ({signal_2516, signal_1108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1186 ( .a ({signal_2415, signal_1180}), .b ({signal_2417, signal_1176}), .c ({signal_2477, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1192 ( .s (signal_4456), .b ({signal_2544, signal_1054}), .a ({signal_2483, signal_1118}), .c ({signal_2586, signal_1438}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1194 ( .s (signal_4456), .b ({signal_2533, signal_1052}), .a ({signal_2481, signal_1116}), .c ({signal_2587, signal_1436}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1196 ( .s (signal_4456), .b ({signal_2522, signal_1050}), .a ({signal_2495, signal_1114}), .c ({signal_2588, signal_1434}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1198 ( .s (signal_4456), .b ({signal_2519, signal_1048}), .a ({signal_2494, signal_1112}), .c ({signal_2589, signal_1432}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1200 ( .s (signal_4456), .b ({signal_2518, signal_1046}), .a ({signal_2508, signal_1110}), .c ({signal_2590, signal_1430}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1202 ( .s (signal_4456), .b ({signal_2549, signal_1044}), .a ({signal_2516, signal_1108}), .c ({signal_2591, signal_1428}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1204 ( .s (signal_4456), .b ({signal_2548, signal_1042}), .a ({signal_2500, signal_1106}), .c ({signal_2592, signal_1426}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1206 ( .s (signal_4456), .b ({signal_2547, signal_1040}), .a ({signal_2499, signal_1104}), .c ({signal_2593, signal_1424}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1208 ( .s (signal_4456), .b ({signal_2546, signal_1038}), .a ({signal_2490, signal_1102}), .c ({signal_2594, signal_1422}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1210 ( .s (signal_4456), .b ({signal_2545, signal_1036}), .a ({signal_2489, signal_1100}), .c ({signal_2595, signal_1420}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1212 ( .s (signal_4456), .b ({signal_2543, signal_1034}), .a ({signal_2478, signal_1098}), .c ({signal_2596, signal_1418}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1214 ( .s (signal_4456), .b ({signal_2542, signal_1032}), .a ({signal_2486, signal_1096}), .c ({signal_2597, signal_1416}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1216 ( .s (signal_4456), .b ({signal_2541, signal_1030}), .a ({signal_2505, signal_1094}), .c ({signal_2598, signal_1414}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1218 ( .s (signal_4456), .b ({signal_2540, signal_1028}), .a ({signal_2504, signal_1092}), .c ({signal_2599, signal_1412}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1220 ( .s (signal_4456), .b ({signal_2539, signal_1026}), .a ({signal_2513, signal_1090}), .c ({signal_2600, signal_1410}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1222 ( .s (signal_4456), .b ({signal_2538, signal_1024}), .a ({signal_2511, signal_1088}), .c ({signal_2601, signal_1408}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1224 ( .s (signal_4456), .b ({signal_2537, signal_1022}), .a ({signal_2515, signal_1086}), .c ({signal_2602, signal_1406}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1226 ( .s (signal_4456), .b ({signal_2536, signal_1020}), .a ({signal_2514, signal_1084}), .c ({signal_2603, signal_1404}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1228 ( .s (signal_4456), .b ({signal_2535, signal_1018}), .a ({signal_2503, signal_1082}), .c ({signal_2604, signal_1402}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1230 ( .s (signal_4456), .b ({signal_2534, signal_1016}), .a ({signal_2501, signal_1080}), .c ({signal_2605, signal_1400}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1232 ( .s (signal_4456), .b ({signal_2532, signal_1014}), .a ({signal_2480, signal_1078}), .c ({signal_2606, signal_1398}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1234 ( .s (signal_4456), .b ({signal_2531, signal_1012}), .a ({signal_2479, signal_1076}), .c ({signal_2607, signal_1396}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1236 ( .s (signal_4456), .b ({signal_2530, signal_1010}), .a ({signal_2488, signal_1074}), .c ({signal_2608, signal_1394}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1238 ( .s (signal_4456), .b ({signal_2529, signal_1008}), .a ({signal_2496, signal_1072}), .c ({signal_2609, signal_1392}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1240 ( .s (signal_4456), .b ({signal_2528, signal_1006}), .a ({signal_2498, signal_1070}), .c ({signal_2610, signal_1390}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1242 ( .s (signal_4456), .b ({signal_2527, signal_1004}), .a ({signal_2506, signal_1068}), .c ({signal_2611, signal_1388}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1244 ( .s (signal_4456), .b ({signal_2526, signal_1002}), .a ({signal_2510, signal_1066}), .c ({signal_2612, signal_1386}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1246 ( .s (signal_4456), .b ({signal_2525, signal_1000}), .a ({signal_2509, signal_1064}), .c ({signal_2613, signal_1384}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1248 ( .s (signal_4456), .b ({signal_2524, signal_998}), .a ({signal_2493, signal_1062}), .c ({signal_2614, signal_1382}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1250 ( .s (signal_4456), .b ({signal_2523, signal_996}), .a ({signal_2491, signal_1060}), .c ({signal_2615, signal_1380}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1252 ( .s (signal_4456), .b ({signal_2521, signal_994}), .a ({signal_2485, signal_1058}), .c ({signal_2616, signal_1378}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1254 ( .s (signal_4456), .b ({signal_2520, signal_992}), .a ({signal_2484, signal_1056}), .c ({signal_2617, signal_1376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .s ({signal_4460, signal_4458}), .b ({signal_2023, signal_1498}), .a ({signal_2037, signal_1507}), .clk (clk), .r (Fresh[135]), .c ({signal_2190, signal_1286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .s ({signal_4468, signal_4464}), .b ({signal_2051, signal_1518}), .a ({signal_2065, signal_1528}), .clk (clk), .r (Fresh[136]), .c ({signal_2192, signal_1256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .s ({signal_4472, signal_4470}), .b ({1'b0, 1'b0}), .a ({signal_2047, signal_1514}), .clk (clk), .r (Fresh[137]), .c ({signal_2193, signal_1591}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .s ({signal_4476, signal_4474}), .b ({signal_2055, signal_1521}), .a ({signal_2077, signal_1536}), .clk (clk), .r (Fresh[138]), .c ({signal_2194, signal_1306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .s ({signal_4476, signal_4474}), .b ({1'b0, 1'b0}), .a ({signal_2031, signal_1503}), .clk (clk), .r (Fresh[139]), .c ({signal_2195, signal_1592}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .s ({signal_4480, signal_4478}), .b ({1'b0, 1'b0}), .a ({signal_2087, signal_1546}), .clk (clk), .r (Fresh[140]), .c ({signal_2196, signal_1593}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .s ({signal_4484, signal_4482}), .b ({signal_2040, signal_1509}), .a ({signal_2096, signal_1554}), .clk (clk), .r (Fresh[141]), .c ({signal_2197, signal_1594}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .s ({signal_4488, signal_4486}), .b ({1'b0, 1'b0}), .a ({signal_2093, signal_1552}), .clk (clk), .r (Fresh[142]), .c ({signal_2198, signal_1595}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .s ({signal_4492, signal_4490}), .b ({signal_2091, signal_1550}), .a ({signal_2062, signal_1526}), .clk (clk), .r (Fresh[143]), .c ({signal_2199, signal_1258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .s ({signal_4496, signal_4494}), .b ({1'b0, 1'b0}), .a ({signal_2042, signal_1511}), .clk (clk), .r (Fresh[144]), .c ({signal_2200, signal_1596}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1400 ( .s ({signal_4476, signal_4474}), .b ({signal_2077, signal_1536}), .a ({signal_2090, signal_1549}), .clk (clk), .r (Fresh[145]), .c ({signal_2201, signal_1597}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1401 ( .s ({signal_4504, signal_4500}), .b ({signal_2080, signal_1539}), .a ({signal_2044, signal_1512}), .clk (clk), .r (Fresh[146]), .c ({signal_2203, signal_1268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1402 ( .s ({signal_4496, signal_4494}), .b ({signal_2089, signal_1548}), .a ({signal_2019, signal_1495}), .clk (clk), .r (Fresh[147]), .c ({signal_2204, signal_1598}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1403 ( .s ({signal_4512, signal_4508}), .b ({signal_2063, signal_1527}), .a ({signal_2095, signal_1553}), .clk (clk), .r (Fresh[148]), .c ({signal_2206, signal_1284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1404 ( .s ({signal_4488, signal_4486}), .b ({signal_2027, signal_1500}), .a ({signal_2081, signal_1540}), .clk (clk), .r (Fresh[149]), .c ({signal_2207, signal_1250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1405 ( .s ({signal_4484, signal_4482}), .b ({signal_2083, signal_1542}), .a ({signal_2040, signal_1509}), .clk (clk), .r (Fresh[150]), .c ({signal_2208, signal_1278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1406 ( .s ({signal_4516, signal_4514}), .b ({signal_2048, signal_1515}), .a ({signal_2021, signal_1497}), .clk (clk), .r (Fresh[151]), .c ({signal_2209, signal_1266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1407 ( .s ({signal_4480, signal_4478}), .b ({signal_2041, signal_1510}), .a ({signal_2066, signal_1529}), .clk (clk), .r (Fresh[152]), .c ({signal_2210, signal_1599}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1408 ( .s ({signal_4524, signal_4520}), .b ({signal_2086, signal_1545}), .a ({signal_2057, signal_1522}), .clk (clk), .r (Fresh[153]), .c ({signal_2212, signal_1292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1409 ( .s ({signal_4516, signal_4514}), .b ({1'b0, 1'b0}), .a ({signal_2049, signal_1516}), .clk (clk), .r (Fresh[154]), .c ({signal_2213, signal_1600}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1410 ( .s ({signal_4516, signal_4514}), .b ({signal_2021, signal_1497}), .a ({signal_2084, signal_1543}), .clk (clk), .r (Fresh[155]), .c ({signal_2214, signal_1601}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1411 ( .s ({signal_4460, signal_4458}), .b ({signal_2037, signal_1507}), .a ({signal_2054, signal_1520}), .clk (clk), .r (Fresh[156]), .c ({signal_2215, signal_1602}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1412 ( .s ({signal_4484, signal_4482}), .b ({1'b0, 1'b0}), .a ({signal_2039, signal_1508}), .clk (clk), .r (Fresh[157]), .c ({signal_2216, signal_1603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1413 ( .s ({signal_4532, signal_4528}), .b ({signal_2074, signal_1534}), .a ({signal_2076, signal_1535}), .clk (clk), .r (Fresh[158]), .c ({signal_2218, signal_1248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1414 ( .s ({signal_4540, signal_4536}), .b ({signal_2061, signal_1525}), .a ({signal_2071, signal_1532}), .clk (clk), .r (Fresh[159]), .c ({signal_2220, signal_1296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1415 ( .s ({signal_4460, signal_4458}), .b ({1'b0, 1'b0}), .a ({signal_2028, signal_1501}), .clk (clk), .r (Fresh[160]), .c ({signal_2221, signal_1604}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .s ({signal_4544, signal_4542}), .b ({signal_2069, signal_1531}), .a ({signal_2082, signal_1541}), .clk (clk), .r (Fresh[161]), .c ({signal_2222, signal_1605}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .s ({signal_4544, signal_4542}), .b ({signal_2060, signal_1524}), .a ({signal_2069, signal_1531}), .clk (clk), .r (Fresh[162]), .c ({signal_2223, signal_1270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .s ({signal_4552, signal_4548}), .b ({signal_2020, signal_1496}), .a ({signal_2053, signal_1519}), .clk (clk), .r (Fresh[163]), .c ({signal_2225, signal_1260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .s ({signal_4560, signal_4556}), .b ({signal_2050, signal_1517}), .a ({signal_2046, signal_1513}), .clk (clk), .r (Fresh[164]), .c ({signal_2227, signal_1276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .s ({signal_4488, signal_4486}), .b ({signal_2081, signal_1540}), .a ({signal_2097, signal_1555}), .clk (clk), .r (Fresh[165]), .c ({signal_2228, signal_1606}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .s ({signal_4544, signal_4542}), .b ({1'b0, 1'b0}), .a ({signal_2078, signal_1537}), .clk (clk), .r (Fresh[166]), .c ({signal_2229, signal_1607}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .s ({signal_4568, signal_4564}), .b ({signal_2079, signal_1538}), .a ({signal_2025, signal_1499}), .clk (clk), .r (Fresh[167]), .c ({signal_2231, signal_1304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .s ({signal_4492, signal_4490}), .b ({1'b0, 1'b0}), .a ({signal_2085, signal_1544}), .clk (clk), .r (Fresh[168]), .c ({signal_2232, signal_1608}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .s ({signal_4576, signal_4572}), .b ({signal_2092, signal_1551}), .a ({signal_2073, signal_1533}), .clk (clk), .r (Fresh[169]), .c ({signal_2234, signal_1264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .s ({signal_4496, signal_4494}), .b ({signal_2029, signal_1502}), .a ({signal_2089, signal_1548}), .clk (clk), .r (Fresh[170]), .c ({signal_2235, signal_1298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .s ({signal_4472, signal_4470}), .b ({signal_2088, signal_1547}), .a ({signal_2032, signal_1504}), .clk (clk), .r (Fresh[171]), .c ({signal_2236, signal_1302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .s ({signal_4492, signal_4490}), .b ({signal_2062, signal_1526}), .a ({signal_2034, signal_1505}), .clk (clk), .r (Fresh[172]), .c ({signal_2237, signal_1609}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .s ({signal_4480, signal_4478}), .b ({signal_2036, signal_1506}), .a ({signal_2041, signal_1510}), .clk (clk), .r (Fresh[173]), .c ({signal_2238, signal_1294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .s ({signal_4584, signal_4580}), .b ({signal_2099, signal_1556}), .a ({signal_2068, signal_1530}), .clk (clk), .r (Fresh[174]), .c ({signal_2240, signal_1308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .s ({signal_4588, signal_4586}), .b ({signal_2101, signal_1558}), .a ({signal_2100, signal_1557}), .clk (clk), .r (Fresh[175]), .c ({signal_2241, signal_1610}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .s ({signal_4592, signal_4590}), .b ({signal_2103, signal_1560}), .a ({signal_2102, signal_1559}), .clk (clk), .r (Fresh[176]), .c ({signal_2242, signal_1611}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .s ({signal_4588, signal_4586}), .b ({signal_2104, signal_1561}), .a ({signal_2101, signal_1558}), .clk (clk), .r (Fresh[177]), .c ({signal_2243, signal_1310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .s ({signal_4588, signal_4586}), .b ({1'b0, 1'b0}), .a ({signal_2105, signal_1562}), .clk (clk), .r (Fresh[178]), .c ({signal_2244, signal_1612}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .s ({signal_4600, signal_4596}), .b ({signal_2108, signal_1564}), .a ({signal_2107, signal_1563}), .clk (clk), .r (Fresh[179]), .c ({signal_2246, signal_1280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .s ({signal_4604, signal_4602}), .b ({signal_2110, signal_1566}), .a ({signal_2109, signal_1565}), .clk (clk), .r (Fresh[180]), .c ({signal_2247, signal_1613}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .s ({signal_4604, signal_4602}), .b ({signal_2111, signal_1567}), .a ({signal_2110, signal_1566}), .clk (clk), .r (Fresh[181]), .c ({signal_2248, signal_1282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .s ({signal_4604, signal_4602}), .b ({1'b0, 1'b0}), .a ({signal_2112, signal_1568}), .clk (clk), .r (Fresh[182]), .c ({signal_2249, signal_1614}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .s ({signal_4612, signal_4608}), .b ({signal_2115, signal_1570}), .a ({signal_2114, signal_1569}), .clk (clk), .r (Fresh[183]), .c ({signal_2251, signal_1252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .s ({signal_4616, signal_4614}), .b ({signal_2117, signal_1572}), .a ({signal_2116, signal_1571}), .clk (clk), .r (Fresh[184]), .c ({signal_2252, signal_1615}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .s ({signal_4616, signal_4614}), .b ({signal_2118, signal_1573}), .a ({signal_2117, signal_1572}), .clk (clk), .r (Fresh[185]), .c ({signal_2253, signal_1254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .s ({signal_4616, signal_4614}), .b ({1'b0, 1'b0}), .a ({signal_2119, signal_1574}), .clk (clk), .r (Fresh[186]), .c ({signal_2254, signal_1616}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .s ({signal_4592, signal_4590}), .b ({signal_2120, signal_1575}), .a ({signal_2103, signal_1560}), .clk (clk), .r (Fresh[187]), .c ({signal_2255, signal_1262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .s ({signal_4624, signal_4620}), .b ({signal_2123, signal_1577}), .a ({signal_2122, signal_1576}), .clk (clk), .r (Fresh[188]), .c ({signal_2257, signal_1272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .s ({signal_4628, signal_4626}), .b ({signal_2125, signal_1579}), .a ({signal_2124, signal_1578}), .clk (clk), .r (Fresh[189]), .c ({signal_2258, signal_1617}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .s ({signal_4628, signal_4626}), .b ({signal_2126, signal_1580}), .a ({signal_2125, signal_1579}), .clk (clk), .r (Fresh[190]), .c ({signal_2259, signal_1274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .s ({signal_4628, signal_4626}), .b ({1'b0, 1'b0}), .a ({signal_2127, signal_1581}), .clk (clk), .r (Fresh[191]), .c ({signal_2260, signal_1618}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .s ({signal_4636, signal_4632}), .b ({signal_2130, signal_1583}), .a ({signal_2129, signal_1582}), .clk (clk), .r (Fresh[192]), .c ({signal_2262, signal_1288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .s ({signal_4640, signal_4638}), .b ({signal_2132, signal_1585}), .a ({signal_2131, signal_1584}), .clk (clk), .r (Fresh[193]), .c ({signal_2263, signal_1619}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .s ({signal_4640, signal_4638}), .b ({signal_2133, signal_1586}), .a ({signal_2132, signal_1585}), .clk (clk), .r (Fresh[194]), .c ({signal_2264, signal_1290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .s ({signal_4640, signal_4638}), .b ({1'b0, 1'b0}), .a ({signal_2134, signal_1587}), .clk (clk), .r (Fresh[195]), .c ({signal_2265, signal_1620}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .s ({signal_4648, signal_4644}), .b ({signal_2058, signal_1523}), .a ({signal_2136, signal_1588}), .clk (clk), .r (Fresh[196]), .c ({signal_2267, signal_1300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .s ({signal_4472, signal_4470}), .b ({signal_2032, signal_1504}), .a ({signal_2137, signal_1589}), .clk (clk), .r (Fresh[197]), .c ({signal_2268, signal_1621}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .s ({signal_4592, signal_4590}), .b ({1'b0, 1'b0}), .a ({signal_2138, signal_1590}), .clk (clk), .r (Fresh[198]), .c ({signal_2269, signal_1622}) ) ;
    buf_clk cell_1555 ( .C (clk), .D (signal_3097), .Q (signal_3098) ) ;
    buf_clk cell_1755 ( .C (clk), .D (signal_3297), .Q (signal_3298) ) ;
    buf_clk cell_1761 ( .C (clk), .D (signal_3303), .Q (signal_3304) ) ;
    buf_clk cell_1767 ( .C (clk), .D (signal_3309), .Q (signal_3310) ) ;
    buf_clk cell_1773 ( .C (clk), .D (signal_3315), .Q (signal_3316) ) ;
    buf_clk cell_1779 ( .C (clk), .D (signal_3321), .Q (signal_3322) ) ;
    buf_clk cell_1785 ( .C (clk), .D (signal_3327), .Q (signal_3328) ) ;
    buf_clk cell_1791 ( .C (clk), .D (signal_3333), .Q (signal_3334) ) ;
    buf_clk cell_1797 ( .C (clk), .D (signal_3339), .Q (signal_3340) ) ;
    buf_clk cell_1803 ( .C (clk), .D (signal_3345), .Q (signal_3346) ) ;
    buf_clk cell_1809 ( .C (clk), .D (signal_3351), .Q (signal_3352) ) ;
    buf_clk cell_1815 ( .C (clk), .D (signal_3357), .Q (signal_3358) ) ;
    buf_clk cell_1821 ( .C (clk), .D (signal_3363), .Q (signal_3364) ) ;
    buf_clk cell_1827 ( .C (clk), .D (signal_3369), .Q (signal_3370) ) ;
    buf_clk cell_1833 ( .C (clk), .D (signal_3375), .Q (signal_3376) ) ;
    buf_clk cell_1839 ( .C (clk), .D (signal_3381), .Q (signal_3382) ) ;
    buf_clk cell_1845 ( .C (clk), .D (signal_3387), .Q (signal_3388) ) ;
    buf_clk cell_1851 ( .C (clk), .D (signal_3393), .Q (signal_3394) ) ;
    buf_clk cell_1857 ( .C (clk), .D (signal_3399), .Q (signal_3400) ) ;
    buf_clk cell_1863 ( .C (clk), .D (signal_3405), .Q (signal_3406) ) ;
    buf_clk cell_1869 ( .C (clk), .D (signal_3411), .Q (signal_3412) ) ;
    buf_clk cell_1875 ( .C (clk), .D (signal_3417), .Q (signal_3418) ) ;
    buf_clk cell_1881 ( .C (clk), .D (signal_3423), .Q (signal_3424) ) ;
    buf_clk cell_1887 ( .C (clk), .D (signal_3429), .Q (signal_3430) ) ;
    buf_clk cell_1893 ( .C (clk), .D (signal_3435), .Q (signal_3436) ) ;
    buf_clk cell_1899 ( .C (clk), .D (signal_3441), .Q (signal_3442) ) ;
    buf_clk cell_1905 ( .C (clk), .D (signal_3447), .Q (signal_3448) ) ;
    buf_clk cell_1911 ( .C (clk), .D (signal_3453), .Q (signal_3454) ) ;
    buf_clk cell_1917 ( .C (clk), .D (signal_3459), .Q (signal_3460) ) ;
    buf_clk cell_1923 ( .C (clk), .D (signal_3465), .Q (signal_3466) ) ;
    buf_clk cell_1929 ( .C (clk), .D (signal_3471), .Q (signal_3472) ) ;
    buf_clk cell_1935 ( .C (clk), .D (signal_3477), .Q (signal_3478) ) ;
    buf_clk cell_1941 ( .C (clk), .D (signal_3483), .Q (signal_3484) ) ;
    buf_clk cell_1947 ( .C (clk), .D (signal_3489), .Q (signal_3490) ) ;
    buf_clk cell_1953 ( .C (clk), .D (signal_3495), .Q (signal_3496) ) ;
    buf_clk cell_1959 ( .C (clk), .D (signal_3501), .Q (signal_3502) ) ;
    buf_clk cell_1965 ( .C (clk), .D (signal_3507), .Q (signal_3508) ) ;
    buf_clk cell_1971 ( .C (clk), .D (signal_3513), .Q (signal_3514) ) ;
    buf_clk cell_1977 ( .C (clk), .D (signal_3519), .Q (signal_3520) ) ;
    buf_clk cell_1983 ( .C (clk), .D (signal_3525), .Q (signal_3526) ) ;
    buf_clk cell_1989 ( .C (clk), .D (signal_3531), .Q (signal_3532) ) ;
    buf_clk cell_1995 ( .C (clk), .D (signal_3537), .Q (signal_3538) ) ;
    buf_clk cell_2001 ( .C (clk), .D (signal_3543), .Q (signal_3544) ) ;
    buf_clk cell_2007 ( .C (clk), .D (signal_3549), .Q (signal_3550) ) ;
    buf_clk cell_2013 ( .C (clk), .D (signal_3555), .Q (signal_3556) ) ;
    buf_clk cell_2019 ( .C (clk), .D (signal_3561), .Q (signal_3562) ) ;
    buf_clk cell_2025 ( .C (clk), .D (signal_3567), .Q (signal_3568) ) ;
    buf_clk cell_2031 ( .C (clk), .D (signal_3573), .Q (signal_3574) ) ;
    buf_clk cell_2037 ( .C (clk), .D (signal_3579), .Q (signal_3580) ) ;
    buf_clk cell_2043 ( .C (clk), .D (signal_3585), .Q (signal_3586) ) ;
    buf_clk cell_2049 ( .C (clk), .D (signal_3591), .Q (signal_3592) ) ;
    buf_clk cell_2055 ( .C (clk), .D (signal_3597), .Q (signal_3598) ) ;
    buf_clk cell_2061 ( .C (clk), .D (signal_3603), .Q (signal_3604) ) ;
    buf_clk cell_2067 ( .C (clk), .D (signal_3609), .Q (signal_3610) ) ;
    buf_clk cell_2073 ( .C (clk), .D (signal_3615), .Q (signal_3616) ) ;
    buf_clk cell_2079 ( .C (clk), .D (signal_3621), .Q (signal_3622) ) ;
    buf_clk cell_2085 ( .C (clk), .D (signal_3627), .Q (signal_3628) ) ;
    buf_clk cell_2091 ( .C (clk), .D (signal_3633), .Q (signal_3634) ) ;
    buf_clk cell_2097 ( .C (clk), .D (signal_3639), .Q (signal_3640) ) ;
    buf_clk cell_2103 ( .C (clk), .D (signal_3645), .Q (signal_3646) ) ;
    buf_clk cell_2109 ( .C (clk), .D (signal_3651), .Q (signal_3652) ) ;
    buf_clk cell_2115 ( .C (clk), .D (signal_3657), .Q (signal_3658) ) ;
    buf_clk cell_2121 ( .C (clk), .D (signal_3663), .Q (signal_3664) ) ;
    buf_clk cell_2127 ( .C (clk), .D (signal_3669), .Q (signal_3670) ) ;
    buf_clk cell_2133 ( .C (clk), .D (signal_3675), .Q (signal_3676) ) ;
    buf_clk cell_2139 ( .C (clk), .D (signal_3681), .Q (signal_3682) ) ;
    buf_clk cell_2145 ( .C (clk), .D (signal_3687), .Q (signal_3688) ) ;
    buf_clk cell_2151 ( .C (clk), .D (signal_3693), .Q (signal_3694) ) ;
    buf_clk cell_2157 ( .C (clk), .D (signal_3699), .Q (signal_3700) ) ;
    buf_clk cell_2163 ( .C (clk), .D (signal_3705), .Q (signal_3706) ) ;
    buf_clk cell_2169 ( .C (clk), .D (signal_3711), .Q (signal_3712) ) ;
    buf_clk cell_2175 ( .C (clk), .D (signal_3717), .Q (signal_3718) ) ;
    buf_clk cell_2181 ( .C (clk), .D (signal_3723), .Q (signal_3724) ) ;
    buf_clk cell_2187 ( .C (clk), .D (signal_3729), .Q (signal_3730) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_3735), .Q (signal_3736) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_3741), .Q (signal_3742) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_3747), .Q (signal_3748) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_3753), .Q (signal_3754) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_3759), .Q (signal_3760) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_3765), .Q (signal_3766) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_3771), .Q (signal_3772) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_3777), .Q (signal_3778) ) ;
    buf_clk cell_2241 ( .C (clk), .D (signal_3783), .Q (signal_3784) ) ;
    buf_clk cell_2247 ( .C (clk), .D (signal_3789), .Q (signal_3790) ) ;
    buf_clk cell_2253 ( .C (clk), .D (signal_3795), .Q (signal_3796) ) ;
    buf_clk cell_2259 ( .C (clk), .D (signal_3801), .Q (signal_3802) ) ;
    buf_clk cell_2265 ( .C (clk), .D (signal_3807), .Q (signal_3808) ) ;
    buf_clk cell_2271 ( .C (clk), .D (signal_3813), .Q (signal_3814) ) ;
    buf_clk cell_2277 ( .C (clk), .D (signal_3819), .Q (signal_3820) ) ;
    buf_clk cell_2283 ( .C (clk), .D (signal_3825), .Q (signal_3826) ) ;
    buf_clk cell_2289 ( .C (clk), .D (signal_3831), .Q (signal_3832) ) ;
    buf_clk cell_2295 ( .C (clk), .D (signal_3837), .Q (signal_3838) ) ;
    buf_clk cell_2301 ( .C (clk), .D (signal_3843), .Q (signal_3844) ) ;
    buf_clk cell_2307 ( .C (clk), .D (signal_3849), .Q (signal_3850) ) ;
    buf_clk cell_2313 ( .C (clk), .D (signal_3855), .Q (signal_3856) ) ;
    buf_clk cell_2319 ( .C (clk), .D (signal_3861), .Q (signal_3862) ) ;
    buf_clk cell_2325 ( .C (clk), .D (signal_3867), .Q (signal_3868) ) ;
    buf_clk cell_2331 ( .C (clk), .D (signal_3873), .Q (signal_3874) ) ;
    buf_clk cell_2337 ( .C (clk), .D (signal_3879), .Q (signal_3880) ) ;
    buf_clk cell_2343 ( .C (clk), .D (signal_3885), .Q (signal_3886) ) ;
    buf_clk cell_2349 ( .C (clk), .D (signal_3891), .Q (signal_3892) ) ;
    buf_clk cell_2355 ( .C (clk), .D (signal_3897), .Q (signal_3898) ) ;
    buf_clk cell_2361 ( .C (clk), .D (signal_3903), .Q (signal_3904) ) ;
    buf_clk cell_2367 ( .C (clk), .D (signal_3909), .Q (signal_3910) ) ;
    buf_clk cell_2373 ( .C (clk), .D (signal_3915), .Q (signal_3916) ) ;
    buf_clk cell_2379 ( .C (clk), .D (signal_3921), .Q (signal_3922) ) ;
    buf_clk cell_2385 ( .C (clk), .D (signal_3927), .Q (signal_3928) ) ;
    buf_clk cell_2391 ( .C (clk), .D (signal_3933), .Q (signal_3934) ) ;
    buf_clk cell_2397 ( .C (clk), .D (signal_3939), .Q (signal_3940) ) ;
    buf_clk cell_2403 ( .C (clk), .D (signal_3945), .Q (signal_3946) ) ;
    buf_clk cell_2409 ( .C (clk), .D (signal_3951), .Q (signal_3952) ) ;
    buf_clk cell_2415 ( .C (clk), .D (signal_3957), .Q (signal_3958) ) ;
    buf_clk cell_2421 ( .C (clk), .D (signal_3963), .Q (signal_3964) ) ;
    buf_clk cell_2427 ( .C (clk), .D (signal_3969), .Q (signal_3970) ) ;
    buf_clk cell_2433 ( .C (clk), .D (signal_3975), .Q (signal_3976) ) ;
    buf_clk cell_2439 ( .C (clk), .D (signal_3981), .Q (signal_3982) ) ;
    buf_clk cell_2445 ( .C (clk), .D (signal_3987), .Q (signal_3988) ) ;
    buf_clk cell_2451 ( .C (clk), .D (signal_3993), .Q (signal_3994) ) ;
    buf_clk cell_2457 ( .C (clk), .D (signal_3999), .Q (signal_4000) ) ;
    buf_clk cell_2463 ( .C (clk), .D (signal_4005), .Q (signal_4006) ) ;
    buf_clk cell_2469 ( .C (clk), .D (signal_4011), .Q (signal_4012) ) ;
    buf_clk cell_2475 ( .C (clk), .D (signal_4017), .Q (signal_4018) ) ;
    buf_clk cell_2481 ( .C (clk), .D (signal_4023), .Q (signal_4024) ) ;
    buf_clk cell_2487 ( .C (clk), .D (signal_4029), .Q (signal_4030) ) ;
    buf_clk cell_2493 ( .C (clk), .D (signal_4035), .Q (signal_4036) ) ;
    buf_clk cell_2499 ( .C (clk), .D (signal_4041), .Q (signal_4042) ) ;
    buf_clk cell_2505 ( .C (clk), .D (signal_4047), .Q (signal_4048) ) ;
    buf_clk cell_2511 ( .C (clk), .D (signal_4053), .Q (signal_4054) ) ;
    buf_clk cell_2517 ( .C (clk), .D (signal_4059), .Q (signal_4060) ) ;
    buf_clk cell_2523 ( .C (clk), .D (signal_4065), .Q (signal_4066) ) ;
    buf_clk cell_2529 ( .C (clk), .D (signal_4071), .Q (signal_4072) ) ;
    buf_clk cell_2535 ( .C (clk), .D (signal_4077), .Q (signal_4078) ) ;
    buf_clk cell_2541 ( .C (clk), .D (signal_4083), .Q (signal_4084) ) ;
    buf_clk cell_2547 ( .C (clk), .D (signal_4089), .Q (signal_4090) ) ;
    buf_clk cell_2553 ( .C (clk), .D (signal_4095), .Q (signal_4096) ) ;
    buf_clk cell_2559 ( .C (clk), .D (signal_4101), .Q (signal_4102) ) ;
    buf_clk cell_2565 ( .C (clk), .D (signal_4107), .Q (signal_4108) ) ;
    buf_clk cell_2571 ( .C (clk), .D (signal_4113), .Q (signal_4114) ) ;
    buf_clk cell_2577 ( .C (clk), .D (signal_4119), .Q (signal_4120) ) ;
    buf_clk cell_2583 ( .C (clk), .D (signal_4125), .Q (signal_4126) ) ;
    buf_clk cell_2589 ( .C (clk), .D (signal_4131), .Q (signal_4132) ) ;
    buf_clk cell_2595 ( .C (clk), .D (signal_4137), .Q (signal_4138) ) ;
    buf_clk cell_2601 ( .C (clk), .D (signal_4143), .Q (signal_4144) ) ;
    buf_clk cell_2607 ( .C (clk), .D (signal_4149), .Q (signal_4150) ) ;
    buf_clk cell_2613 ( .C (clk), .D (signal_4155), .Q (signal_4156) ) ;
    buf_clk cell_2619 ( .C (clk), .D (signal_4161), .Q (signal_4162) ) ;
    buf_clk cell_2625 ( .C (clk), .D (signal_4167), .Q (signal_4168) ) ;
    buf_clk cell_2631 ( .C (clk), .D (signal_4173), .Q (signal_4174) ) ;
    buf_clk cell_2637 ( .C (clk), .D (signal_4179), .Q (signal_4180) ) ;
    buf_clk cell_2643 ( .C (clk), .D (signal_4185), .Q (signal_4186) ) ;
    buf_clk cell_2649 ( .C (clk), .D (signal_4191), .Q (signal_4192) ) ;
    buf_clk cell_2655 ( .C (clk), .D (signal_4197), .Q (signal_4198) ) ;
    buf_clk cell_2661 ( .C (clk), .D (signal_4203), .Q (signal_4204) ) ;
    buf_clk cell_2667 ( .C (clk), .D (signal_4209), .Q (signal_4210) ) ;
    buf_clk cell_2673 ( .C (clk), .D (signal_4215), .Q (signal_4216) ) ;
    buf_clk cell_2679 ( .C (clk), .D (signal_4221), .Q (signal_4222) ) ;
    buf_clk cell_2685 ( .C (clk), .D (signal_4227), .Q (signal_4228) ) ;
    buf_clk cell_2691 ( .C (clk), .D (signal_4233), .Q (signal_4234) ) ;
    buf_clk cell_2697 ( .C (clk), .D (signal_4239), .Q (signal_4240) ) ;
    buf_clk cell_2703 ( .C (clk), .D (signal_4245), .Q (signal_4246) ) ;
    buf_clk cell_2709 ( .C (clk), .D (signal_4251), .Q (signal_4252) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_4257), .Q (signal_4258) ) ;
    buf_clk cell_2721 ( .C (clk), .D (signal_4263), .Q (signal_4264) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_4269), .Q (signal_4270) ) ;
    buf_clk cell_2733 ( .C (clk), .D (signal_4275), .Q (signal_4276) ) ;
    buf_clk cell_2739 ( .C (clk), .D (signal_4281), .Q (signal_4282) ) ;
    buf_clk cell_2745 ( .C (clk), .D (signal_4287), .Q (signal_4288) ) ;
    buf_clk cell_2751 ( .C (clk), .D (signal_4293), .Q (signal_4294) ) ;
    buf_clk cell_2757 ( .C (clk), .D (signal_4299), .Q (signal_4300) ) ;
    buf_clk cell_2763 ( .C (clk), .D (signal_4305), .Q (signal_4306) ) ;
    buf_clk cell_2769 ( .C (clk), .D (signal_4311), .Q (signal_4312) ) ;
    buf_clk cell_2775 ( .C (clk), .D (signal_4317), .Q (signal_4318) ) ;
    buf_clk cell_2781 ( .C (clk), .D (signal_4323), .Q (signal_4324) ) ;
    buf_clk cell_2787 ( .C (clk), .D (signal_4329), .Q (signal_4330) ) ;
    buf_clk cell_2793 ( .C (clk), .D (signal_4335), .Q (signal_4336) ) ;
    buf_clk cell_2799 ( .C (clk), .D (signal_4341), .Q (signal_4342) ) ;
    buf_clk cell_2805 ( .C (clk), .D (signal_4347), .Q (signal_4348) ) ;
    buf_clk cell_2811 ( .C (clk), .D (signal_4353), .Q (signal_4354) ) ;
    buf_clk cell_2817 ( .C (clk), .D (signal_4359), .Q (signal_4360) ) ;
    buf_clk cell_2823 ( .C (clk), .D (signal_4365), .Q (signal_4366) ) ;
    buf_clk cell_2829 ( .C (clk), .D (signal_4371), .Q (signal_4372) ) ;
    buf_clk cell_2835 ( .C (clk), .D (signal_4377), .Q (signal_4378) ) ;
    buf_clk cell_2841 ( .C (clk), .D (signal_4383), .Q (signal_4384) ) ;
    buf_clk cell_2847 ( .C (clk), .D (signal_4389), .Q (signal_4390) ) ;
    buf_clk cell_2853 ( .C (clk), .D (signal_4395), .Q (signal_4396) ) ;
    buf_clk cell_2859 ( .C (clk), .D (signal_4401), .Q (signal_4402) ) ;
    buf_clk cell_2865 ( .C (clk), .D (signal_4407), .Q (signal_4408) ) ;
    buf_clk cell_2871 ( .C (clk), .D (signal_4413), .Q (signal_4414) ) ;
    buf_clk cell_2877 ( .C (clk), .D (signal_4419), .Q (signal_4420) ) ;
    buf_clk cell_2883 ( .C (clk), .D (signal_4425), .Q (signal_4426) ) ;
    buf_clk cell_2889 ( .C (clk), .D (signal_4431), .Q (signal_4432) ) ;
    buf_clk cell_2895 ( .C (clk), .D (signal_4437), .Q (signal_4438) ) ;
    buf_clk cell_2901 ( .C (clk), .D (signal_4443), .Q (signal_4444) ) ;
    buf_clk cell_2907 ( .C (clk), .D (signal_4449), .Q (signal_4450) ) ;
    buf_clk cell_2913 ( .C (clk), .D (signal_4455), .Q (signal_4456) ) ;
    buf_clk cell_3111 ( .C (clk), .D (signal_4653), .Q (signal_4654) ) ;
    buf_clk cell_3119 ( .C (clk), .D (signal_4661), .Q (signal_4662) ) ;
    buf_clk cell_3127 ( .C (clk), .D (signal_4669), .Q (signal_4670) ) ;
    buf_clk cell_3135 ( .C (clk), .D (signal_4677), .Q (signal_4678) ) ;
    buf_clk cell_3143 ( .C (clk), .D (signal_4685), .Q (signal_4686) ) ;
    buf_clk cell_3151 ( .C (clk), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_3159 ( .C (clk), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_3167 ( .C (clk), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_3175 ( .C (clk), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_3183 ( .C (clk), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_3191 ( .C (clk), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_3199 ( .C (clk), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_3207 ( .C (clk), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_3215 ( .C (clk), .D (signal_4757), .Q (signal_4758) ) ;
    buf_clk cell_3223 ( .C (clk), .D (signal_4765), .Q (signal_4766) ) ;
    buf_clk cell_3231 ( .C (clk), .D (signal_4773), .Q (signal_4774) ) ;
    buf_clk cell_3239 ( .C (clk), .D (signal_4781), .Q (signal_4782) ) ;
    buf_clk cell_3247 ( .C (clk), .D (signal_4789), .Q (signal_4790) ) ;
    buf_clk cell_3255 ( .C (clk), .D (signal_4797), .Q (signal_4798) ) ;
    buf_clk cell_3263 ( .C (clk), .D (signal_4805), .Q (signal_4806) ) ;
    buf_clk cell_3271 ( .C (clk), .D (signal_4813), .Q (signal_4814) ) ;
    buf_clk cell_3279 ( .C (clk), .D (signal_4821), .Q (signal_4822) ) ;
    buf_clk cell_3287 ( .C (clk), .D (signal_4829), .Q (signal_4830) ) ;
    buf_clk cell_3295 ( .C (clk), .D (signal_4837), .Q (signal_4838) ) ;
    buf_clk cell_3303 ( .C (clk), .D (signal_4845), .Q (signal_4846) ) ;
    buf_clk cell_3311 ( .C (clk), .D (signal_4853), .Q (signal_4854) ) ;
    buf_clk cell_3319 ( .C (clk), .D (signal_4861), .Q (signal_4862) ) ;
    buf_clk cell_3327 ( .C (clk), .D (signal_4869), .Q (signal_4870) ) ;
    buf_clk cell_3335 ( .C (clk), .D (signal_4877), .Q (signal_4878) ) ;
    buf_clk cell_3343 ( .C (clk), .D (signal_4885), .Q (signal_4886) ) ;
    buf_clk cell_3351 ( .C (clk), .D (signal_4893), .Q (signal_4894) ) ;
    buf_clk cell_3359 ( .C (clk), .D (signal_4901), .Q (signal_4902) ) ;
    buf_clk cell_3367 ( .C (clk), .D (signal_4909), .Q (signal_4910) ) ;
    buf_clk cell_3375 ( .C (clk), .D (signal_4917), .Q (signal_4918) ) ;
    buf_clk cell_3383 ( .C (clk), .D (signal_4925), .Q (signal_4926) ) ;
    buf_clk cell_3391 ( .C (clk), .D (signal_4933), .Q (signal_4934) ) ;
    buf_clk cell_3399 ( .C (clk), .D (signal_4941), .Q (signal_4942) ) ;
    buf_clk cell_3407 ( .C (clk), .D (signal_4949), .Q (signal_4950) ) ;
    buf_clk cell_3415 ( .C (clk), .D (signal_4957), .Q (signal_4958) ) ;
    buf_clk cell_3423 ( .C (clk), .D (signal_4965), .Q (signal_4966) ) ;
    buf_clk cell_3431 ( .C (clk), .D (signal_4973), .Q (signal_4974) ) ;
    buf_clk cell_3439 ( .C (clk), .D (signal_4981), .Q (signal_4982) ) ;
    buf_clk cell_3447 ( .C (clk), .D (signal_4989), .Q (signal_4990) ) ;
    buf_clk cell_3455 ( .C (clk), .D (signal_4997), .Q (signal_4998) ) ;
    buf_clk cell_3463 ( .C (clk), .D (signal_5005), .Q (signal_5006) ) ;
    buf_clk cell_3471 ( .C (clk), .D (signal_5013), .Q (signal_5014) ) ;
    buf_clk cell_3479 ( .C (clk), .D (signal_5021), .Q (signal_5022) ) ;
    buf_clk cell_3487 ( .C (clk), .D (signal_5029), .Q (signal_5030) ) ;
    buf_clk cell_3495 ( .C (clk), .D (signal_5037), .Q (signal_5038) ) ;
    buf_clk cell_3503 ( .C (clk), .D (signal_5045), .Q (signal_5046) ) ;
    buf_clk cell_3511 ( .C (clk), .D (signal_5053), .Q (signal_5054) ) ;
    buf_clk cell_3519 ( .C (clk), .D (signal_5061), .Q (signal_5062) ) ;
    buf_clk cell_3527 ( .C (clk), .D (signal_5069), .Q (signal_5070) ) ;
    buf_clk cell_3535 ( .C (clk), .D (signal_5077), .Q (signal_5078) ) ;
    buf_clk cell_3543 ( .C (clk), .D (signal_5085), .Q (signal_5086) ) ;
    buf_clk cell_3551 ( .C (clk), .D (signal_5093), .Q (signal_5094) ) ;
    buf_clk cell_3559 ( .C (clk), .D (signal_5101), .Q (signal_5102) ) ;
    buf_clk cell_3567 ( .C (clk), .D (signal_5109), .Q (signal_5110) ) ;
    buf_clk cell_3575 ( .C (clk), .D (signal_5117), .Q (signal_5118) ) ;
    buf_clk cell_3583 ( .C (clk), .D (signal_5125), .Q (signal_5126) ) ;
    buf_clk cell_3591 ( .C (clk), .D (signal_5133), .Q (signal_5134) ) ;
    buf_clk cell_3599 ( .C (clk), .D (signal_5141), .Q (signal_5142) ) ;
    buf_clk cell_3607 ( .C (clk), .D (signal_5149), .Q (signal_5150) ) ;
    buf_clk cell_3615 ( .C (clk), .D (signal_5157), .Q (signal_5158) ) ;
    buf_clk cell_3623 ( .C (clk), .D (signal_5165), .Q (signal_5166) ) ;
    buf_clk cell_3631 ( .C (clk), .D (signal_5173), .Q (signal_5174) ) ;
    buf_clk cell_3639 ( .C (clk), .D (signal_5181), .Q (signal_5182) ) ;
    buf_clk cell_3647 ( .C (clk), .D (signal_5189), .Q (signal_5190) ) ;
    buf_clk cell_3655 ( .C (clk), .D (signal_5197), .Q (signal_5198) ) ;
    buf_clk cell_3663 ( .C (clk), .D (signal_5205), .Q (signal_5206) ) ;
    buf_clk cell_3671 ( .C (clk), .D (signal_5213), .Q (signal_5214) ) ;
    buf_clk cell_3679 ( .C (clk), .D (signal_5221), .Q (signal_5222) ) ;
    buf_clk cell_3687 ( .C (clk), .D (signal_5229), .Q (signal_5230) ) ;
    buf_clk cell_3695 ( .C (clk), .D (signal_5237), .Q (signal_5238) ) ;
    buf_clk cell_3703 ( .C (clk), .D (signal_5245), .Q (signal_5246) ) ;
    buf_clk cell_3711 ( .C (clk), .D (signal_5253), .Q (signal_5254) ) ;
    buf_clk cell_3719 ( .C (clk), .D (signal_5261), .Q (signal_5262) ) ;
    buf_clk cell_3727 ( .C (clk), .D (signal_5269), .Q (signal_5270) ) ;
    buf_clk cell_3735 ( .C (clk), .D (signal_5277), .Q (signal_5278) ) ;
    buf_clk cell_3743 ( .C (clk), .D (signal_5285), .Q (signal_5286) ) ;
    buf_clk cell_3751 ( .C (clk), .D (signal_5293), .Q (signal_5294) ) ;
    buf_clk cell_3759 ( .C (clk), .D (signal_5301), .Q (signal_5302) ) ;
    buf_clk cell_3767 ( .C (clk), .D (signal_5309), .Q (signal_5310) ) ;
    buf_clk cell_3775 ( .C (clk), .D (signal_5317), .Q (signal_5318) ) ;
    buf_clk cell_3783 ( .C (clk), .D (signal_5325), .Q (signal_5326) ) ;
    buf_clk cell_3791 ( .C (clk), .D (signal_5333), .Q (signal_5334) ) ;
    buf_clk cell_3799 ( .C (clk), .D (signal_5341), .Q (signal_5342) ) ;
    buf_clk cell_3807 ( .C (clk), .D (signal_5349), .Q (signal_5350) ) ;
    buf_clk cell_3815 ( .C (clk), .D (signal_5357), .Q (signal_5358) ) ;
    buf_clk cell_3823 ( .C (clk), .D (signal_5365), .Q (signal_5366) ) ;
    buf_clk cell_3831 ( .C (clk), .D (signal_5373), .Q (signal_5374) ) ;
    buf_clk cell_3839 ( .C (clk), .D (signal_5381), .Q (signal_5382) ) ;
    buf_clk cell_3847 ( .C (clk), .D (signal_5389), .Q (signal_5390) ) ;
    buf_clk cell_3855 ( .C (clk), .D (signal_5397), .Q (signal_5398) ) ;
    buf_clk cell_3863 ( .C (clk), .D (signal_5405), .Q (signal_5406) ) ;
    buf_clk cell_3871 ( .C (clk), .D (signal_5413), .Q (signal_5414) ) ;
    buf_clk cell_3879 ( .C (clk), .D (signal_5421), .Q (signal_5422) ) ;
    buf_clk cell_3887 ( .C (clk), .D (signal_5429), .Q (signal_5430) ) ;
    buf_clk cell_3895 ( .C (clk), .D (signal_5437), .Q (signal_5438) ) ;
    buf_clk cell_3903 ( .C (clk), .D (signal_5445), .Q (signal_5446) ) ;
    buf_clk cell_3911 ( .C (clk), .D (signal_5453), .Q (signal_5454) ) ;
    buf_clk cell_3919 ( .C (clk), .D (signal_5461), .Q (signal_5462) ) ;
    buf_clk cell_3927 ( .C (clk), .D (signal_5469), .Q (signal_5470) ) ;
    buf_clk cell_3935 ( .C (clk), .D (signal_5477), .Q (signal_5478) ) ;
    buf_clk cell_3943 ( .C (clk), .D (signal_5485), .Q (signal_5486) ) ;
    buf_clk cell_3951 ( .C (clk), .D (signal_5493), .Q (signal_5494) ) ;
    buf_clk cell_3959 ( .C (clk), .D (signal_5501), .Q (signal_5502) ) ;
    buf_clk cell_3967 ( .C (clk), .D (signal_5509), .Q (signal_5510) ) ;
    buf_clk cell_3975 ( .C (clk), .D (signal_5517), .Q (signal_5518) ) ;
    buf_clk cell_3983 ( .C (clk), .D (signal_5525), .Q (signal_5526) ) ;
    buf_clk cell_3991 ( .C (clk), .D (signal_5533), .Q (signal_5534) ) ;
    buf_clk cell_3999 ( .C (clk), .D (signal_5541), .Q (signal_5542) ) ;
    buf_clk cell_4007 ( .C (clk), .D (signal_5549), .Q (signal_5550) ) ;
    buf_clk cell_4015 ( .C (clk), .D (signal_5557), .Q (signal_5558) ) ;
    buf_clk cell_4023 ( .C (clk), .D (signal_5565), .Q (signal_5566) ) ;
    buf_clk cell_4031 ( .C (clk), .D (signal_5573), .Q (signal_5574) ) ;
    buf_clk cell_4039 ( .C (clk), .D (signal_5581), .Q (signal_5582) ) ;
    buf_clk cell_4047 ( .C (clk), .D (signal_5589), .Q (signal_5590) ) ;
    buf_clk cell_4055 ( .C (clk), .D (signal_5597), .Q (signal_5598) ) ;
    buf_clk cell_4063 ( .C (clk), .D (signal_5605), .Q (signal_5606) ) ;
    buf_clk cell_4071 ( .C (clk), .D (signal_5613), .Q (signal_5614) ) ;
    buf_clk cell_4079 ( .C (clk), .D (signal_5621), .Q (signal_5622) ) ;
    buf_clk cell_4087 ( .C (clk), .D (signal_5629), .Q (signal_5630) ) ;
    buf_clk cell_4095 ( .C (clk), .D (signal_5637), .Q (signal_5638) ) ;
    buf_clk cell_4103 ( .C (clk), .D (signal_5645), .Q (signal_5646) ) ;
    buf_clk cell_4111 ( .C (clk), .D (signal_5653), .Q (signal_5654) ) ;
    buf_clk cell_4119 ( .C (clk), .D (signal_5661), .Q (signal_5662) ) ;
    buf_clk cell_4127 ( .C (clk), .D (signal_5669), .Q (signal_5670) ) ;
    buf_clk cell_4137 ( .C (clk), .D (signal_5679), .Q (signal_5680) ) ;
    buf_clk cell_4145 ( .C (clk), .D (signal_5687), .Q (signal_5688) ) ;
    buf_clk cell_4153 ( .C (clk), .D (signal_5695), .Q (signal_5696) ) ;
    buf_clk cell_4161 ( .C (clk), .D (signal_5703), .Q (signal_5704) ) ;
    buf_clk cell_4169 ( .C (clk), .D (signal_5711), .Q (signal_5712) ) ;
    buf_clk cell_4177 ( .C (clk), .D (signal_5719), .Q (signal_5720) ) ;
    buf_clk cell_4185 ( .C (clk), .D (signal_5727), .Q (signal_5728) ) ;
    buf_clk cell_4193 ( .C (clk), .D (signal_5735), .Q (signal_5736) ) ;
    buf_clk cell_4201 ( .C (clk), .D (signal_5743), .Q (signal_5744) ) ;
    buf_clk cell_4209 ( .C (clk), .D (signal_5751), .Q (signal_5752) ) ;
    buf_clk cell_4217 ( .C (clk), .D (signal_5759), .Q (signal_5760) ) ;
    buf_clk cell_4225 ( .C (clk), .D (signal_5767), .Q (signal_5768) ) ;
    buf_clk cell_4233 ( .C (clk), .D (signal_5775), .Q (signal_5776) ) ;
    buf_clk cell_4241 ( .C (clk), .D (signal_5783), .Q (signal_5784) ) ;
    buf_clk cell_4249 ( .C (clk), .D (signal_5791), .Q (signal_5792) ) ;
    buf_clk cell_4257 ( .C (clk), .D (signal_5799), .Q (signal_5800) ) ;
    buf_clk cell_4265 ( .C (clk), .D (signal_5807), .Q (signal_5808) ) ;
    buf_clk cell_4273 ( .C (clk), .D (signal_5815), .Q (signal_5816) ) ;
    buf_clk cell_4281 ( .C (clk), .D (signal_5823), .Q (signal_5824) ) ;
    buf_clk cell_4289 ( .C (clk), .D (signal_5831), .Q (signal_5832) ) ;
    buf_clk cell_4297 ( .C (clk), .D (signal_5839), .Q (signal_5840) ) ;
    buf_clk cell_4305 ( .C (clk), .D (signal_5847), .Q (signal_5848) ) ;
    buf_clk cell_4313 ( .C (clk), .D (signal_5855), .Q (signal_5856) ) ;
    buf_clk cell_4321 ( .C (clk), .D (signal_5863), .Q (signal_5864) ) ;
    buf_clk cell_4329 ( .C (clk), .D (signal_5871), .Q (signal_5872) ) ;
    buf_clk cell_4337 ( .C (clk), .D (signal_5879), .Q (signal_5880) ) ;
    buf_clk cell_4345 ( .C (clk), .D (signal_5887), .Q (signal_5888) ) ;
    buf_clk cell_4353 ( .C (clk), .D (signal_5895), .Q (signal_5896) ) ;
    buf_clk cell_4361 ( .C (clk), .D (signal_5903), .Q (signal_5904) ) ;
    buf_clk cell_4369 ( .C (clk), .D (signal_5911), .Q (signal_5912) ) ;
    buf_clk cell_4377 ( .C (clk), .D (signal_5919), .Q (signal_5920) ) ;
    buf_clk cell_4385 ( .C (clk), .D (signal_5927), .Q (signal_5928) ) ;
    buf_clk cell_4393 ( .C (clk), .D (signal_5935), .Q (signal_5936) ) ;
    buf_clk cell_4401 ( .C (clk), .D (signal_5943), .Q (signal_5944) ) ;
    buf_clk cell_4409 ( .C (clk), .D (signal_5951), .Q (signal_5952) ) ;
    buf_clk cell_4417 ( .C (clk), .D (signal_5959), .Q (signal_5960) ) ;
    buf_clk cell_4425 ( .C (clk), .D (signal_5967), .Q (signal_5968) ) ;
    buf_clk cell_4433 ( .C (clk), .D (signal_5975), .Q (signal_5976) ) ;
    buf_clk cell_4441 ( .C (clk), .D (signal_5983), .Q (signal_5984) ) ;
    buf_clk cell_4449 ( .C (clk), .D (signal_5991), .Q (signal_5992) ) ;
    buf_clk cell_4457 ( .C (clk), .D (signal_5999), .Q (signal_6000) ) ;
    buf_clk cell_4465 ( .C (clk), .D (signal_6007), .Q (signal_6008) ) ;
    buf_clk cell_4473 ( .C (clk), .D (signal_6015), .Q (signal_6016) ) ;
    buf_clk cell_4481 ( .C (clk), .D (signal_6023), .Q (signal_6024) ) ;
    buf_clk cell_4489 ( .C (clk), .D (signal_6031), .Q (signal_6032) ) ;
    buf_clk cell_4497 ( .C (clk), .D (signal_6039), .Q (signal_6040) ) ;
    buf_clk cell_4505 ( .C (clk), .D (signal_6047), .Q (signal_6048) ) ;
    buf_clk cell_4513 ( .C (clk), .D (signal_6055), .Q (signal_6056) ) ;
    buf_clk cell_4521 ( .C (clk), .D (signal_6063), .Q (signal_6064) ) ;
    buf_clk cell_4529 ( .C (clk), .D (signal_6071), .Q (signal_6072) ) ;
    buf_clk cell_4537 ( .C (clk), .D (signal_6079), .Q (signal_6080) ) ;
    buf_clk cell_4545 ( .C (clk), .D (signal_6087), .Q (signal_6088) ) ;
    buf_clk cell_4553 ( .C (clk), .D (signal_6095), .Q (signal_6096) ) ;
    buf_clk cell_4561 ( .C (clk), .D (signal_6103), .Q (signal_6104) ) ;
    buf_clk cell_4569 ( .C (clk), .D (signal_6111), .Q (signal_6112) ) ;
    buf_clk cell_4577 ( .C (clk), .D (signal_6119), .Q (signal_6120) ) ;
    buf_clk cell_4585 ( .C (clk), .D (signal_6127), .Q (signal_6128) ) ;
    buf_clk cell_4593 ( .C (clk), .D (signal_6135), .Q (signal_6136) ) ;
    buf_clk cell_4601 ( .C (clk), .D (signal_6143), .Q (signal_6144) ) ;
    buf_clk cell_4609 ( .C (clk), .D (signal_6151), .Q (signal_6152) ) ;
    buf_clk cell_4617 ( .C (clk), .D (signal_6159), .Q (signal_6160) ) ;
    buf_clk cell_4625 ( .C (clk), .D (signal_6167), .Q (signal_6168) ) ;
    buf_clk cell_4633 ( .C (clk), .D (signal_6175), .Q (signal_6176) ) ;
    buf_clk cell_4641 ( .C (clk), .D (signal_6183), .Q (signal_6184) ) ;
    buf_clk cell_4647 ( .C (clk), .D (signal_6189), .Q (signal_6190) ) ;
    buf_clk cell_4649 ( .C (clk), .D (signal_6191), .Q (signal_6192) ) ;
    buf_clk cell_4651 ( .C (clk), .D (signal_6193), .Q (signal_6194) ) ;
    buf_clk cell_4653 ( .C (clk), .D (signal_6195), .Q (signal_6196) ) ;
    buf_clk cell_4655 ( .C (clk), .D (signal_6197), .Q (signal_6198) ) ;
    buf_clk cell_4657 ( .C (clk), .D (signal_6199), .Q (signal_6200) ) ;
    buf_clk cell_4659 ( .C (clk), .D (signal_6201), .Q (signal_6202) ) ;
    buf_clk cell_4661 ( .C (clk), .D (signal_6203), .Q (signal_6204) ) ;
    buf_clk cell_4663 ( .C (clk), .D (signal_6205), .Q (signal_6206) ) ;
    buf_clk cell_4665 ( .C (clk), .D (signal_6207), .Q (signal_6208) ) ;
    buf_clk cell_4667 ( .C (clk), .D (signal_6209), .Q (signal_6210) ) ;
    buf_clk cell_4669 ( .C (clk), .D (signal_6211), .Q (signal_6212) ) ;
    buf_clk cell_4671 ( .C (clk), .D (signal_6213), .Q (signal_6214) ) ;
    buf_clk cell_4673 ( .C (clk), .D (signal_6215), .Q (signal_6216) ) ;
    buf_clk cell_4675 ( .C (clk), .D (signal_6217), .Q (signal_6218) ) ;
    buf_clk cell_4677 ( .C (clk), .D (signal_6219), .Q (signal_6220) ) ;
    buf_clk cell_4679 ( .C (clk), .D (signal_6221), .Q (signal_6222) ) ;
    buf_clk cell_4681 ( .C (clk), .D (signal_6223), .Q (signal_6224) ) ;
    buf_clk cell_4683 ( .C (clk), .D (signal_6225), .Q (signal_6226) ) ;
    buf_clk cell_4685 ( .C (clk), .D (signal_6227), .Q (signal_6228) ) ;
    buf_clk cell_4687 ( .C (clk), .D (signal_6229), .Q (signal_6230) ) ;
    buf_clk cell_4689 ( .C (clk), .D (signal_6231), .Q (signal_6232) ) ;
    buf_clk cell_4691 ( .C (clk), .D (signal_6233), .Q (signal_6234) ) ;
    buf_clk cell_4693 ( .C (clk), .D (signal_6235), .Q (signal_6236) ) ;
    buf_clk cell_4695 ( .C (clk), .D (signal_6237), .Q (signal_6238) ) ;
    buf_clk cell_4697 ( .C (clk), .D (signal_6239), .Q (signal_6240) ) ;
    buf_clk cell_4699 ( .C (clk), .D (signal_6241), .Q (signal_6242) ) ;
    buf_clk cell_4701 ( .C (clk), .D (signal_6243), .Q (signal_6244) ) ;
    buf_clk cell_4703 ( .C (clk), .D (signal_6245), .Q (signal_6246) ) ;
    buf_clk cell_4705 ( .C (clk), .D (signal_6247), .Q (signal_6248) ) ;
    buf_clk cell_4707 ( .C (clk), .D (signal_6249), .Q (signal_6250) ) ;
    buf_clk cell_4709 ( .C (clk), .D (signal_6251), .Q (signal_6252) ) ;
    buf_clk cell_4711 ( .C (clk), .D (signal_6253), .Q (signal_6254) ) ;
    buf_clk cell_4713 ( .C (clk), .D (signal_6255), .Q (signal_6256) ) ;
    buf_clk cell_4715 ( .C (clk), .D (signal_6257), .Q (signal_6258) ) ;
    buf_clk cell_4717 ( .C (clk), .D (signal_6259), .Q (signal_6260) ) ;
    buf_clk cell_4719 ( .C (clk), .D (signal_6261), .Q (signal_6262) ) ;
    buf_clk cell_4721 ( .C (clk), .D (signal_6263), .Q (signal_6264) ) ;
    buf_clk cell_4723 ( .C (clk), .D (signal_6265), .Q (signal_6266) ) ;
    buf_clk cell_4725 ( .C (clk), .D (signal_6267), .Q (signal_6268) ) ;
    buf_clk cell_4727 ( .C (clk), .D (signal_6269), .Q (signal_6270) ) ;
    buf_clk cell_4729 ( .C (clk), .D (signal_6271), .Q (signal_6272) ) ;
    buf_clk cell_4731 ( .C (clk), .D (signal_6273), .Q (signal_6274) ) ;
    buf_clk cell_4733 ( .C (clk), .D (signal_6275), .Q (signal_6276) ) ;
    buf_clk cell_4735 ( .C (clk), .D (signal_6277), .Q (signal_6278) ) ;
    buf_clk cell_4737 ( .C (clk), .D (signal_6279), .Q (signal_6280) ) ;
    buf_clk cell_4739 ( .C (clk), .D (signal_6281), .Q (signal_6282) ) ;
    buf_clk cell_4741 ( .C (clk), .D (signal_6283), .Q (signal_6284) ) ;
    buf_clk cell_4743 ( .C (clk), .D (signal_6285), .Q (signal_6286) ) ;
    buf_clk cell_4745 ( .C (clk), .D (signal_6287), .Q (signal_6288) ) ;
    buf_clk cell_4747 ( .C (clk), .D (signal_6289), .Q (signal_6290) ) ;
    buf_clk cell_4749 ( .C (clk), .D (signal_6291), .Q (signal_6292) ) ;
    buf_clk cell_4751 ( .C (clk), .D (signal_6293), .Q (signal_6294) ) ;
    buf_clk cell_4753 ( .C (clk), .D (signal_6295), .Q (signal_6296) ) ;
    buf_clk cell_4755 ( .C (clk), .D (signal_6297), .Q (signal_6298) ) ;
    buf_clk cell_4757 ( .C (clk), .D (signal_6299), .Q (signal_6300) ) ;
    buf_clk cell_4759 ( .C (clk), .D (signal_6301), .Q (signal_6302) ) ;
    buf_clk cell_4761 ( .C (clk), .D (signal_6303), .Q (signal_6304) ) ;
    buf_clk cell_4763 ( .C (clk), .D (signal_6305), .Q (signal_6306) ) ;
    buf_clk cell_4765 ( .C (clk), .D (signal_6307), .Q (signal_6308) ) ;
    buf_clk cell_4767 ( .C (clk), .D (signal_6309), .Q (signal_6310) ) ;
    buf_clk cell_4769 ( .C (clk), .D (signal_6311), .Q (signal_6312) ) ;
    buf_clk cell_4771 ( .C (clk), .D (signal_6313), .Q (signal_6314) ) ;
    buf_clk cell_4773 ( .C (clk), .D (signal_6315), .Q (signal_6316) ) ;
    buf_clk cell_4775 ( .C (clk), .D (signal_6317), .Q (signal_6318) ) ;
    buf_clk cell_4777 ( .C (clk), .D (signal_6319), .Q (signal_6320) ) ;
    buf_clk cell_4779 ( .C (clk), .D (signal_6321), .Q (signal_6322) ) ;
    buf_clk cell_4781 ( .C (clk), .D (signal_6323), .Q (signal_6324) ) ;
    buf_clk cell_4783 ( .C (clk), .D (signal_6325), .Q (signal_6326) ) ;
    buf_clk cell_4785 ( .C (clk), .D (signal_6327), .Q (signal_6328) ) ;
    buf_clk cell_4787 ( .C (clk), .D (signal_6329), .Q (signal_6330) ) ;
    buf_clk cell_4789 ( .C (clk), .D (signal_6331), .Q (signal_6332) ) ;
    buf_clk cell_4791 ( .C (clk), .D (signal_6333), .Q (signal_6334) ) ;
    buf_clk cell_4793 ( .C (clk), .D (signal_6335), .Q (signal_6336) ) ;
    buf_clk cell_4795 ( .C (clk), .D (signal_6337), .Q (signal_6338) ) ;
    buf_clk cell_4797 ( .C (clk), .D (signal_6339), .Q (signal_6340) ) ;
    buf_clk cell_4799 ( .C (clk), .D (signal_6341), .Q (signal_6342) ) ;
    buf_clk cell_4801 ( .C (clk), .D (signal_6343), .Q (signal_6344) ) ;
    buf_clk cell_4803 ( .C (clk), .D (signal_6345), .Q (signal_6346) ) ;
    buf_clk cell_4805 ( .C (clk), .D (signal_6347), .Q (signal_6348) ) ;
    buf_clk cell_4807 ( .C (clk), .D (signal_6349), .Q (signal_6350) ) ;
    buf_clk cell_4809 ( .C (clk), .D (signal_6351), .Q (signal_6352) ) ;
    buf_clk cell_4811 ( .C (clk), .D (signal_6353), .Q (signal_6354) ) ;
    buf_clk cell_4813 ( .C (clk), .D (signal_6355), .Q (signal_6356) ) ;
    buf_clk cell_4815 ( .C (clk), .D (signal_6357), .Q (signal_6358) ) ;
    buf_clk cell_4817 ( .C (clk), .D (signal_6359), .Q (signal_6360) ) ;
    buf_clk cell_4819 ( .C (clk), .D (signal_6361), .Q (signal_6362) ) ;
    buf_clk cell_4821 ( .C (clk), .D (signal_6363), .Q (signal_6364) ) ;
    buf_clk cell_4823 ( .C (clk), .D (signal_6365), .Q (signal_6366) ) ;
    buf_clk cell_4825 ( .C (clk), .D (signal_6367), .Q (signal_6368) ) ;
    buf_clk cell_4827 ( .C (clk), .D (signal_6369), .Q (signal_6370) ) ;
    buf_clk cell_4829 ( .C (clk), .D (signal_6371), .Q (signal_6372) ) ;
    buf_clk cell_4831 ( .C (clk), .D (signal_6373), .Q (signal_6374) ) ;
    buf_clk cell_4833 ( .C (clk), .D (signal_6375), .Q (signal_6376) ) ;
    buf_clk cell_4835 ( .C (clk), .D (signal_6377), .Q (signal_6378) ) ;
    buf_clk cell_4837 ( .C (clk), .D (signal_6379), .Q (signal_6380) ) ;
    buf_clk cell_4843 ( .C (clk), .D (signal_6385), .Q (signal_6386) ) ;
    buf_clk cell_4851 ( .C (clk), .D (signal_6393), .Q (signal_6394) ) ;
    buf_clk cell_4859 ( .C (clk), .D (signal_6401), .Q (signal_6402) ) ;
    buf_clk cell_4867 ( .C (clk), .D (signal_6409), .Q (signal_6410) ) ;

    /* cells in depth 7 */
    buf_clk cell_1486 ( .C (clk), .D (signal_201), .Q (signal_3029) ) ;
    buf_clk cell_1488 ( .C (clk), .D (signal_203), .Q (signal_3031) ) ;
    buf_clk cell_1490 ( .C (clk), .D (signal_205), .Q (signal_3033) ) ;
    buf_clk cell_1492 ( .C (clk), .D (signal_207), .Q (signal_3035) ) ;
    buf_clk cell_1494 ( .C (clk), .D (signal_209), .Q (signal_3037) ) ;
    buf_clk cell_1496 ( .C (clk), .D (signal_211), .Q (signal_3039) ) ;
    buf_clk cell_1498 ( .C (clk), .D (signal_213), .Q (signal_3041) ) ;
    buf_clk cell_1500 ( .C (clk), .D (signal_215), .Q (signal_3043) ) ;
    buf_clk cell_1502 ( .C (clk), .D (signal_217), .Q (signal_3045) ) ;
    buf_clk cell_1504 ( .C (clk), .D (signal_219), .Q (signal_3047) ) ;
    buf_clk cell_1506 ( .C (clk), .D (signal_221), .Q (signal_3049) ) ;
    buf_clk cell_1508 ( .C (clk), .D (signal_223), .Q (signal_3051) ) ;
    buf_clk cell_1510 ( .C (clk), .D (signal_225), .Q (signal_3053) ) ;
    buf_clk cell_1512 ( .C (clk), .D (signal_227), .Q (signal_3055) ) ;
    buf_clk cell_1514 ( .C (clk), .D (signal_229), .Q (signal_3057) ) ;
    buf_clk cell_1516 ( .C (clk), .D (signal_231), .Q (signal_3059) ) ;
    buf_clk cell_1518 ( .C (clk), .D (signal_233), .Q (signal_3061) ) ;
    buf_clk cell_1520 ( .C (clk), .D (signal_235), .Q (signal_3063) ) ;
    buf_clk cell_1522 ( .C (clk), .D (signal_237), .Q (signal_3065) ) ;
    buf_clk cell_1524 ( .C (clk), .D (signal_239), .Q (signal_3067) ) ;
    buf_clk cell_1526 ( .C (clk), .D (signal_241), .Q (signal_3069) ) ;
    buf_clk cell_1528 ( .C (clk), .D (signal_243), .Q (signal_3071) ) ;
    buf_clk cell_1530 ( .C (clk), .D (signal_245), .Q (signal_3073) ) ;
    buf_clk cell_1532 ( .C (clk), .D (signal_247), .Q (signal_3075) ) ;
    buf_clk cell_1534 ( .C (clk), .D (signal_249), .Q (signal_3077) ) ;
    buf_clk cell_1536 ( .C (clk), .D (signal_251), .Q (signal_3079) ) ;
    buf_clk cell_1538 ( .C (clk), .D (signal_253), .Q (signal_3081) ) ;
    buf_clk cell_1540 ( .C (clk), .D (signal_255), .Q (signal_3083) ) ;
    buf_clk cell_1542 ( .C (clk), .D (signal_257), .Q (signal_3085) ) ;
    buf_clk cell_1544 ( .C (clk), .D (signal_259), .Q (signal_3087) ) ;
    buf_clk cell_1546 ( .C (clk), .D (signal_261), .Q (signal_3089) ) ;
    buf_clk cell_1548 ( .C (clk), .D (signal_263), .Q (signal_3091) ) ;
    buf_clk cell_1556 ( .C (clk), .D (signal_3098), .Q (signal_3099) ) ;
    buf_clk cell_1558 ( .C (clk), .D (signal_2270), .Q (signal_3101) ) ;
    buf_clk cell_1560 ( .C (clk), .D (signal_2271), .Q (signal_3103) ) ;
    buf_clk cell_1562 ( .C (clk), .D (signal_2272), .Q (signal_3105) ) ;
    buf_clk cell_1564 ( .C (clk), .D (signal_2273), .Q (signal_3107) ) ;
    buf_clk cell_1566 ( .C (clk), .D (signal_2274), .Q (signal_3109) ) ;
    buf_clk cell_1568 ( .C (clk), .D (signal_2275), .Q (signal_3111) ) ;
    buf_clk cell_1570 ( .C (clk), .D (signal_2276), .Q (signal_3113) ) ;
    buf_clk cell_1572 ( .C (clk), .D (signal_2277), .Q (signal_3115) ) ;
    buf_clk cell_1574 ( .C (clk), .D (signal_2278), .Q (signal_3117) ) ;
    buf_clk cell_1576 ( .C (clk), .D (signal_2279), .Q (signal_3119) ) ;
    buf_clk cell_1578 ( .C (clk), .D (signal_2280), .Q (signal_3121) ) ;
    buf_clk cell_1580 ( .C (clk), .D (signal_2281), .Q (signal_3123) ) ;
    buf_clk cell_1582 ( .C (clk), .D (signal_2282), .Q (signal_3125) ) ;
    buf_clk cell_1584 ( .C (clk), .D (signal_2283), .Q (signal_3127) ) ;
    buf_clk cell_1586 ( .C (clk), .D (signal_2284), .Q (signal_3129) ) ;
    buf_clk cell_1588 ( .C (clk), .D (signal_2285), .Q (signal_3131) ) ;
    buf_clk cell_1590 ( .C (clk), .D (signal_2286), .Q (signal_3133) ) ;
    buf_clk cell_1592 ( .C (clk), .D (signal_2287), .Q (signal_3135) ) ;
    buf_clk cell_1594 ( .C (clk), .D (signal_2288), .Q (signal_3137) ) ;
    buf_clk cell_1596 ( .C (clk), .D (signal_2289), .Q (signal_3139) ) ;
    buf_clk cell_1598 ( .C (clk), .D (signal_2290), .Q (signal_3141) ) ;
    buf_clk cell_1600 ( .C (clk), .D (signal_2291), .Q (signal_3143) ) ;
    buf_clk cell_1602 ( .C (clk), .D (signal_2292), .Q (signal_3145) ) ;
    buf_clk cell_1604 ( .C (clk), .D (signal_2293), .Q (signal_3147) ) ;
    buf_clk cell_1606 ( .C (clk), .D (signal_2294), .Q (signal_3149) ) ;
    buf_clk cell_1608 ( .C (clk), .D (signal_2295), .Q (signal_3151) ) ;
    buf_clk cell_1610 ( .C (clk), .D (signal_2296), .Q (signal_3153) ) ;
    buf_clk cell_1612 ( .C (clk), .D (signal_2297), .Q (signal_3155) ) ;
    buf_clk cell_1614 ( .C (clk), .D (signal_2298), .Q (signal_3157) ) ;
    buf_clk cell_1616 ( .C (clk), .D (signal_2299), .Q (signal_3159) ) ;
    buf_clk cell_1618 ( .C (clk), .D (signal_2300), .Q (signal_3161) ) ;
    buf_clk cell_1620 ( .C (clk), .D (signal_2301), .Q (signal_3163) ) ;
    buf_clk cell_3112 ( .C (clk), .D (signal_4654), .Q (signal_4655) ) ;
    buf_clk cell_3120 ( .C (clk), .D (signal_4662), .Q (signal_4663) ) ;
    buf_clk cell_3128 ( .C (clk), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_3136 ( .C (clk), .D (signal_4678), .Q (signal_4679) ) ;
    buf_clk cell_3144 ( .C (clk), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_3152 ( .C (clk), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_3160 ( .C (clk), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_3168 ( .C (clk), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_3176 ( .C (clk), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_3184 ( .C (clk), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_3192 ( .C (clk), .D (signal_4734), .Q (signal_4735) ) ;
    buf_clk cell_3200 ( .C (clk), .D (signal_4742), .Q (signal_4743) ) ;
    buf_clk cell_3208 ( .C (clk), .D (signal_4750), .Q (signal_4751) ) ;
    buf_clk cell_3216 ( .C (clk), .D (signal_4758), .Q (signal_4759) ) ;
    buf_clk cell_3224 ( .C (clk), .D (signal_4766), .Q (signal_4767) ) ;
    buf_clk cell_3232 ( .C (clk), .D (signal_4774), .Q (signal_4775) ) ;
    buf_clk cell_3240 ( .C (clk), .D (signal_4782), .Q (signal_4783) ) ;
    buf_clk cell_3248 ( .C (clk), .D (signal_4790), .Q (signal_4791) ) ;
    buf_clk cell_3256 ( .C (clk), .D (signal_4798), .Q (signal_4799) ) ;
    buf_clk cell_3264 ( .C (clk), .D (signal_4806), .Q (signal_4807) ) ;
    buf_clk cell_3272 ( .C (clk), .D (signal_4814), .Q (signal_4815) ) ;
    buf_clk cell_3280 ( .C (clk), .D (signal_4822), .Q (signal_4823) ) ;
    buf_clk cell_3288 ( .C (clk), .D (signal_4830), .Q (signal_4831) ) ;
    buf_clk cell_3296 ( .C (clk), .D (signal_4838), .Q (signal_4839) ) ;
    buf_clk cell_3304 ( .C (clk), .D (signal_4846), .Q (signal_4847) ) ;
    buf_clk cell_3312 ( .C (clk), .D (signal_4854), .Q (signal_4855) ) ;
    buf_clk cell_3320 ( .C (clk), .D (signal_4862), .Q (signal_4863) ) ;
    buf_clk cell_3328 ( .C (clk), .D (signal_4870), .Q (signal_4871) ) ;
    buf_clk cell_3336 ( .C (clk), .D (signal_4878), .Q (signal_4879) ) ;
    buf_clk cell_3344 ( .C (clk), .D (signal_4886), .Q (signal_4887) ) ;
    buf_clk cell_3352 ( .C (clk), .D (signal_4894), .Q (signal_4895) ) ;
    buf_clk cell_3360 ( .C (clk), .D (signal_4902), .Q (signal_4903) ) ;
    buf_clk cell_3368 ( .C (clk), .D (signal_4910), .Q (signal_4911) ) ;
    buf_clk cell_3376 ( .C (clk), .D (signal_4918), .Q (signal_4919) ) ;
    buf_clk cell_3384 ( .C (clk), .D (signal_4926), .Q (signal_4927) ) ;
    buf_clk cell_3392 ( .C (clk), .D (signal_4934), .Q (signal_4935) ) ;
    buf_clk cell_3400 ( .C (clk), .D (signal_4942), .Q (signal_4943) ) ;
    buf_clk cell_3408 ( .C (clk), .D (signal_4950), .Q (signal_4951) ) ;
    buf_clk cell_3416 ( .C (clk), .D (signal_4958), .Q (signal_4959) ) ;
    buf_clk cell_3424 ( .C (clk), .D (signal_4966), .Q (signal_4967) ) ;
    buf_clk cell_3432 ( .C (clk), .D (signal_4974), .Q (signal_4975) ) ;
    buf_clk cell_3440 ( .C (clk), .D (signal_4982), .Q (signal_4983) ) ;
    buf_clk cell_3448 ( .C (clk), .D (signal_4990), .Q (signal_4991) ) ;
    buf_clk cell_3456 ( .C (clk), .D (signal_4998), .Q (signal_4999) ) ;
    buf_clk cell_3464 ( .C (clk), .D (signal_5006), .Q (signal_5007) ) ;
    buf_clk cell_3472 ( .C (clk), .D (signal_5014), .Q (signal_5015) ) ;
    buf_clk cell_3480 ( .C (clk), .D (signal_5022), .Q (signal_5023) ) ;
    buf_clk cell_3488 ( .C (clk), .D (signal_5030), .Q (signal_5031) ) ;
    buf_clk cell_3496 ( .C (clk), .D (signal_5038), .Q (signal_5039) ) ;
    buf_clk cell_3504 ( .C (clk), .D (signal_5046), .Q (signal_5047) ) ;
    buf_clk cell_3512 ( .C (clk), .D (signal_5054), .Q (signal_5055) ) ;
    buf_clk cell_3520 ( .C (clk), .D (signal_5062), .Q (signal_5063) ) ;
    buf_clk cell_3528 ( .C (clk), .D (signal_5070), .Q (signal_5071) ) ;
    buf_clk cell_3536 ( .C (clk), .D (signal_5078), .Q (signal_5079) ) ;
    buf_clk cell_3544 ( .C (clk), .D (signal_5086), .Q (signal_5087) ) ;
    buf_clk cell_3552 ( .C (clk), .D (signal_5094), .Q (signal_5095) ) ;
    buf_clk cell_3560 ( .C (clk), .D (signal_5102), .Q (signal_5103) ) ;
    buf_clk cell_3568 ( .C (clk), .D (signal_5110), .Q (signal_5111) ) ;
    buf_clk cell_3576 ( .C (clk), .D (signal_5118), .Q (signal_5119) ) ;
    buf_clk cell_3584 ( .C (clk), .D (signal_5126), .Q (signal_5127) ) ;
    buf_clk cell_3592 ( .C (clk), .D (signal_5134), .Q (signal_5135) ) ;
    buf_clk cell_3600 ( .C (clk), .D (signal_5142), .Q (signal_5143) ) ;
    buf_clk cell_3608 ( .C (clk), .D (signal_5150), .Q (signal_5151) ) ;
    buf_clk cell_3616 ( .C (clk), .D (signal_5158), .Q (signal_5159) ) ;
    buf_clk cell_3624 ( .C (clk), .D (signal_5166), .Q (signal_5167) ) ;
    buf_clk cell_3632 ( .C (clk), .D (signal_5174), .Q (signal_5175) ) ;
    buf_clk cell_3640 ( .C (clk), .D (signal_5182), .Q (signal_5183) ) ;
    buf_clk cell_3648 ( .C (clk), .D (signal_5190), .Q (signal_5191) ) ;
    buf_clk cell_3656 ( .C (clk), .D (signal_5198), .Q (signal_5199) ) ;
    buf_clk cell_3664 ( .C (clk), .D (signal_5206), .Q (signal_5207) ) ;
    buf_clk cell_3672 ( .C (clk), .D (signal_5214), .Q (signal_5215) ) ;
    buf_clk cell_3680 ( .C (clk), .D (signal_5222), .Q (signal_5223) ) ;
    buf_clk cell_3688 ( .C (clk), .D (signal_5230), .Q (signal_5231) ) ;
    buf_clk cell_3696 ( .C (clk), .D (signal_5238), .Q (signal_5239) ) ;
    buf_clk cell_3704 ( .C (clk), .D (signal_5246), .Q (signal_5247) ) ;
    buf_clk cell_3712 ( .C (clk), .D (signal_5254), .Q (signal_5255) ) ;
    buf_clk cell_3720 ( .C (clk), .D (signal_5262), .Q (signal_5263) ) ;
    buf_clk cell_3728 ( .C (clk), .D (signal_5270), .Q (signal_5271) ) ;
    buf_clk cell_3736 ( .C (clk), .D (signal_5278), .Q (signal_5279) ) ;
    buf_clk cell_3744 ( .C (clk), .D (signal_5286), .Q (signal_5287) ) ;
    buf_clk cell_3752 ( .C (clk), .D (signal_5294), .Q (signal_5295) ) ;
    buf_clk cell_3760 ( .C (clk), .D (signal_5302), .Q (signal_5303) ) ;
    buf_clk cell_3768 ( .C (clk), .D (signal_5310), .Q (signal_5311) ) ;
    buf_clk cell_3776 ( .C (clk), .D (signal_5318), .Q (signal_5319) ) ;
    buf_clk cell_3784 ( .C (clk), .D (signal_5326), .Q (signal_5327) ) ;
    buf_clk cell_3792 ( .C (clk), .D (signal_5334), .Q (signal_5335) ) ;
    buf_clk cell_3800 ( .C (clk), .D (signal_5342), .Q (signal_5343) ) ;
    buf_clk cell_3808 ( .C (clk), .D (signal_5350), .Q (signal_5351) ) ;
    buf_clk cell_3816 ( .C (clk), .D (signal_5358), .Q (signal_5359) ) ;
    buf_clk cell_3824 ( .C (clk), .D (signal_5366), .Q (signal_5367) ) ;
    buf_clk cell_3832 ( .C (clk), .D (signal_5374), .Q (signal_5375) ) ;
    buf_clk cell_3840 ( .C (clk), .D (signal_5382), .Q (signal_5383) ) ;
    buf_clk cell_3848 ( .C (clk), .D (signal_5390), .Q (signal_5391) ) ;
    buf_clk cell_3856 ( .C (clk), .D (signal_5398), .Q (signal_5399) ) ;
    buf_clk cell_3864 ( .C (clk), .D (signal_5406), .Q (signal_5407) ) ;
    buf_clk cell_3872 ( .C (clk), .D (signal_5414), .Q (signal_5415) ) ;
    buf_clk cell_3880 ( .C (clk), .D (signal_5422), .Q (signal_5423) ) ;
    buf_clk cell_3888 ( .C (clk), .D (signal_5430), .Q (signal_5431) ) ;
    buf_clk cell_3896 ( .C (clk), .D (signal_5438), .Q (signal_5439) ) ;
    buf_clk cell_3904 ( .C (clk), .D (signal_5446), .Q (signal_5447) ) ;
    buf_clk cell_3912 ( .C (clk), .D (signal_5454), .Q (signal_5455) ) ;
    buf_clk cell_3920 ( .C (clk), .D (signal_5462), .Q (signal_5463) ) ;
    buf_clk cell_3928 ( .C (clk), .D (signal_5470), .Q (signal_5471) ) ;
    buf_clk cell_3936 ( .C (clk), .D (signal_5478), .Q (signal_5479) ) ;
    buf_clk cell_3944 ( .C (clk), .D (signal_5486), .Q (signal_5487) ) ;
    buf_clk cell_3952 ( .C (clk), .D (signal_5494), .Q (signal_5495) ) ;
    buf_clk cell_3960 ( .C (clk), .D (signal_5502), .Q (signal_5503) ) ;
    buf_clk cell_3968 ( .C (clk), .D (signal_5510), .Q (signal_5511) ) ;
    buf_clk cell_3976 ( .C (clk), .D (signal_5518), .Q (signal_5519) ) ;
    buf_clk cell_3984 ( .C (clk), .D (signal_5526), .Q (signal_5527) ) ;
    buf_clk cell_3992 ( .C (clk), .D (signal_5534), .Q (signal_5535) ) ;
    buf_clk cell_4000 ( .C (clk), .D (signal_5542), .Q (signal_5543) ) ;
    buf_clk cell_4008 ( .C (clk), .D (signal_5550), .Q (signal_5551) ) ;
    buf_clk cell_4016 ( .C (clk), .D (signal_5558), .Q (signal_5559) ) ;
    buf_clk cell_4024 ( .C (clk), .D (signal_5566), .Q (signal_5567) ) ;
    buf_clk cell_4032 ( .C (clk), .D (signal_5574), .Q (signal_5575) ) ;
    buf_clk cell_4040 ( .C (clk), .D (signal_5582), .Q (signal_5583) ) ;
    buf_clk cell_4048 ( .C (clk), .D (signal_5590), .Q (signal_5591) ) ;
    buf_clk cell_4056 ( .C (clk), .D (signal_5598), .Q (signal_5599) ) ;
    buf_clk cell_4064 ( .C (clk), .D (signal_5606), .Q (signal_5607) ) ;
    buf_clk cell_4072 ( .C (clk), .D (signal_5614), .Q (signal_5615) ) ;
    buf_clk cell_4080 ( .C (clk), .D (signal_5622), .Q (signal_5623) ) ;
    buf_clk cell_4088 ( .C (clk), .D (signal_5630), .Q (signal_5631) ) ;
    buf_clk cell_4096 ( .C (clk), .D (signal_5638), .Q (signal_5639) ) ;
    buf_clk cell_4104 ( .C (clk), .D (signal_5646), .Q (signal_5647) ) ;
    buf_clk cell_4112 ( .C (clk), .D (signal_5654), .Q (signal_5655) ) ;
    buf_clk cell_4120 ( .C (clk), .D (signal_5662), .Q (signal_5663) ) ;
    buf_clk cell_4128 ( .C (clk), .D (signal_5670), .Q (signal_5671) ) ;
    buf_clk cell_4130 ( .C (clk), .D (signal_4066), .Q (signal_5673) ) ;
    buf_clk cell_4138 ( .C (clk), .D (signal_5680), .Q (signal_5681) ) ;
    buf_clk cell_4146 ( .C (clk), .D (signal_5688), .Q (signal_5689) ) ;
    buf_clk cell_4154 ( .C (clk), .D (signal_5696), .Q (signal_5697) ) ;
    buf_clk cell_4162 ( .C (clk), .D (signal_5704), .Q (signal_5705) ) ;
    buf_clk cell_4170 ( .C (clk), .D (signal_5712), .Q (signal_5713) ) ;
    buf_clk cell_4178 ( .C (clk), .D (signal_5720), .Q (signal_5721) ) ;
    buf_clk cell_4186 ( .C (clk), .D (signal_5728), .Q (signal_5729) ) ;
    buf_clk cell_4194 ( .C (clk), .D (signal_5736), .Q (signal_5737) ) ;
    buf_clk cell_4202 ( .C (clk), .D (signal_5744), .Q (signal_5745) ) ;
    buf_clk cell_4210 ( .C (clk), .D (signal_5752), .Q (signal_5753) ) ;
    buf_clk cell_4218 ( .C (clk), .D (signal_5760), .Q (signal_5761) ) ;
    buf_clk cell_4226 ( .C (clk), .D (signal_5768), .Q (signal_5769) ) ;
    buf_clk cell_4234 ( .C (clk), .D (signal_5776), .Q (signal_5777) ) ;
    buf_clk cell_4242 ( .C (clk), .D (signal_5784), .Q (signal_5785) ) ;
    buf_clk cell_4250 ( .C (clk), .D (signal_5792), .Q (signal_5793) ) ;
    buf_clk cell_4258 ( .C (clk), .D (signal_5800), .Q (signal_5801) ) ;
    buf_clk cell_4266 ( .C (clk), .D (signal_5808), .Q (signal_5809) ) ;
    buf_clk cell_4274 ( .C (clk), .D (signal_5816), .Q (signal_5817) ) ;
    buf_clk cell_4282 ( .C (clk), .D (signal_5824), .Q (signal_5825) ) ;
    buf_clk cell_4290 ( .C (clk), .D (signal_5832), .Q (signal_5833) ) ;
    buf_clk cell_4298 ( .C (clk), .D (signal_5840), .Q (signal_5841) ) ;
    buf_clk cell_4306 ( .C (clk), .D (signal_5848), .Q (signal_5849) ) ;
    buf_clk cell_4314 ( .C (clk), .D (signal_5856), .Q (signal_5857) ) ;
    buf_clk cell_4322 ( .C (clk), .D (signal_5864), .Q (signal_5865) ) ;
    buf_clk cell_4330 ( .C (clk), .D (signal_5872), .Q (signal_5873) ) ;
    buf_clk cell_4338 ( .C (clk), .D (signal_5880), .Q (signal_5881) ) ;
    buf_clk cell_4346 ( .C (clk), .D (signal_5888), .Q (signal_5889) ) ;
    buf_clk cell_4354 ( .C (clk), .D (signal_5896), .Q (signal_5897) ) ;
    buf_clk cell_4362 ( .C (clk), .D (signal_5904), .Q (signal_5905) ) ;
    buf_clk cell_4370 ( .C (clk), .D (signal_5912), .Q (signal_5913) ) ;
    buf_clk cell_4378 ( .C (clk), .D (signal_5920), .Q (signal_5921) ) ;
    buf_clk cell_4386 ( .C (clk), .D (signal_5928), .Q (signal_5929) ) ;
    buf_clk cell_4394 ( .C (clk), .D (signal_5936), .Q (signal_5937) ) ;
    buf_clk cell_4402 ( .C (clk), .D (signal_5944), .Q (signal_5945) ) ;
    buf_clk cell_4410 ( .C (clk), .D (signal_5952), .Q (signal_5953) ) ;
    buf_clk cell_4418 ( .C (clk), .D (signal_5960), .Q (signal_5961) ) ;
    buf_clk cell_4426 ( .C (clk), .D (signal_5968), .Q (signal_5969) ) ;
    buf_clk cell_4434 ( .C (clk), .D (signal_5976), .Q (signal_5977) ) ;
    buf_clk cell_4442 ( .C (clk), .D (signal_5984), .Q (signal_5985) ) ;
    buf_clk cell_4450 ( .C (clk), .D (signal_5992), .Q (signal_5993) ) ;
    buf_clk cell_4458 ( .C (clk), .D (signal_6000), .Q (signal_6001) ) ;
    buf_clk cell_4466 ( .C (clk), .D (signal_6008), .Q (signal_6009) ) ;
    buf_clk cell_4474 ( .C (clk), .D (signal_6016), .Q (signal_6017) ) ;
    buf_clk cell_4482 ( .C (clk), .D (signal_6024), .Q (signal_6025) ) ;
    buf_clk cell_4490 ( .C (clk), .D (signal_6032), .Q (signal_6033) ) ;
    buf_clk cell_4498 ( .C (clk), .D (signal_6040), .Q (signal_6041) ) ;
    buf_clk cell_4506 ( .C (clk), .D (signal_6048), .Q (signal_6049) ) ;
    buf_clk cell_4514 ( .C (clk), .D (signal_6056), .Q (signal_6057) ) ;
    buf_clk cell_4522 ( .C (clk), .D (signal_6064), .Q (signal_6065) ) ;
    buf_clk cell_4530 ( .C (clk), .D (signal_6072), .Q (signal_6073) ) ;
    buf_clk cell_4538 ( .C (clk), .D (signal_6080), .Q (signal_6081) ) ;
    buf_clk cell_4546 ( .C (clk), .D (signal_6088), .Q (signal_6089) ) ;
    buf_clk cell_4554 ( .C (clk), .D (signal_6096), .Q (signal_6097) ) ;
    buf_clk cell_4562 ( .C (clk), .D (signal_6104), .Q (signal_6105) ) ;
    buf_clk cell_4570 ( .C (clk), .D (signal_6112), .Q (signal_6113) ) ;
    buf_clk cell_4578 ( .C (clk), .D (signal_6120), .Q (signal_6121) ) ;
    buf_clk cell_4586 ( .C (clk), .D (signal_6128), .Q (signal_6129) ) ;
    buf_clk cell_4594 ( .C (clk), .D (signal_6136), .Q (signal_6137) ) ;
    buf_clk cell_4602 ( .C (clk), .D (signal_6144), .Q (signal_6145) ) ;
    buf_clk cell_4610 ( .C (clk), .D (signal_6152), .Q (signal_6153) ) ;
    buf_clk cell_4618 ( .C (clk), .D (signal_6160), .Q (signal_6161) ) ;
    buf_clk cell_4626 ( .C (clk), .D (signal_6168), .Q (signal_6169) ) ;
    buf_clk cell_4634 ( .C (clk), .D (signal_6176), .Q (signal_6177) ) ;
    buf_clk cell_4642 ( .C (clk), .D (signal_6184), .Q (signal_6185) ) ;
    buf_clk cell_4644 ( .C (clk), .D (signal_4456), .Q (signal_6187) ) ;
    buf_clk cell_4844 ( .C (clk), .D (signal_6386), .Q (signal_6387) ) ;
    buf_clk cell_4852 ( .C (clk), .D (signal_6394), .Q (signal_6395) ) ;
    buf_clk cell_4860 ( .C (clk), .D (signal_6402), .Q (signal_6403) ) ;
    buf_clk cell_4868 ( .C (clk), .D (signal_6410), .Q (signal_6411) ) ;
    buf_clk cell_4870 ( .C (clk), .D (signal_462), .Q (signal_6413) ) ;
    buf_clk cell_4872 ( .C (clk), .D (signal_2632), .Q (signal_6415) ) ;
    buf_clk cell_4874 ( .C (clk), .D (signal_466), .Q (signal_6417) ) ;
    buf_clk cell_4876 ( .C (clk), .D (signal_2633), .Q (signal_6419) ) ;
    buf_clk cell_4878 ( .C (clk), .D (signal_470), .Q (signal_6421) ) ;
    buf_clk cell_4880 ( .C (clk), .D (signal_2634), .Q (signal_6423) ) ;
    buf_clk cell_4882 ( .C (clk), .D (signal_474), .Q (signal_6425) ) ;
    buf_clk cell_4884 ( .C (clk), .D (signal_2635), .Q (signal_6427) ) ;
    buf_clk cell_4886 ( .C (clk), .D (signal_478), .Q (signal_6429) ) ;
    buf_clk cell_4888 ( .C (clk), .D (signal_2636), .Q (signal_6431) ) ;
    buf_clk cell_4890 ( .C (clk), .D (signal_482), .Q (signal_6433) ) ;
    buf_clk cell_4892 ( .C (clk), .D (signal_2637), .Q (signal_6435) ) ;
    buf_clk cell_4894 ( .C (clk), .D (signal_486), .Q (signal_6437) ) ;
    buf_clk cell_4896 ( .C (clk), .D (signal_2638), .Q (signal_6439) ) ;
    buf_clk cell_4898 ( .C (clk), .D (signal_490), .Q (signal_6441) ) ;
    buf_clk cell_4900 ( .C (clk), .D (signal_2639), .Q (signal_6443) ) ;
    buf_clk cell_4902 ( .C (clk), .D (signal_494), .Q (signal_6445) ) ;
    buf_clk cell_4904 ( .C (clk), .D (signal_2640), .Q (signal_6447) ) ;
    buf_clk cell_4906 ( .C (clk), .D (signal_498), .Q (signal_6449) ) ;
    buf_clk cell_4908 ( .C (clk), .D (signal_2641), .Q (signal_6451) ) ;
    buf_clk cell_4910 ( .C (clk), .D (signal_502), .Q (signal_6453) ) ;
    buf_clk cell_4912 ( .C (clk), .D (signal_2642), .Q (signal_6455) ) ;
    buf_clk cell_4914 ( .C (clk), .D (signal_506), .Q (signal_6457) ) ;
    buf_clk cell_4916 ( .C (clk), .D (signal_2643), .Q (signal_6459) ) ;
    buf_clk cell_4918 ( .C (clk), .D (signal_510), .Q (signal_6461) ) ;
    buf_clk cell_4920 ( .C (clk), .D (signal_2644), .Q (signal_6463) ) ;
    buf_clk cell_4922 ( .C (clk), .D (signal_514), .Q (signal_6465) ) ;
    buf_clk cell_4924 ( .C (clk), .D (signal_2645), .Q (signal_6467) ) ;
    buf_clk cell_4926 ( .C (clk), .D (signal_518), .Q (signal_6469) ) ;
    buf_clk cell_4928 ( .C (clk), .D (signal_2646), .Q (signal_6471) ) ;
    buf_clk cell_4930 ( .C (clk), .D (signal_522), .Q (signal_6473) ) ;
    buf_clk cell_4932 ( .C (clk), .D (signal_2647), .Q (signal_6475) ) ;
    buf_clk cell_4934 ( .C (clk), .D (signal_526), .Q (signal_6477) ) ;
    buf_clk cell_4936 ( .C (clk), .D (signal_2648), .Q (signal_6479) ) ;
    buf_clk cell_4938 ( .C (clk), .D (signal_530), .Q (signal_6481) ) ;
    buf_clk cell_4940 ( .C (clk), .D (signal_2649), .Q (signal_6483) ) ;
    buf_clk cell_4942 ( .C (clk), .D (signal_534), .Q (signal_6485) ) ;
    buf_clk cell_4944 ( .C (clk), .D (signal_2650), .Q (signal_6487) ) ;
    buf_clk cell_4946 ( .C (clk), .D (signal_538), .Q (signal_6489) ) ;
    buf_clk cell_4948 ( .C (clk), .D (signal_2651), .Q (signal_6491) ) ;
    buf_clk cell_4950 ( .C (clk), .D (signal_542), .Q (signal_6493) ) ;
    buf_clk cell_4952 ( .C (clk), .D (signal_2652), .Q (signal_6495) ) ;
    buf_clk cell_4954 ( .C (clk), .D (signal_546), .Q (signal_6497) ) ;
    buf_clk cell_4956 ( .C (clk), .D (signal_2653), .Q (signal_6499) ) ;
    buf_clk cell_4958 ( .C (clk), .D (signal_550), .Q (signal_6501) ) ;
    buf_clk cell_4960 ( .C (clk), .D (signal_2654), .Q (signal_6503) ) ;
    buf_clk cell_4962 ( .C (clk), .D (signal_554), .Q (signal_6505) ) ;
    buf_clk cell_4964 ( .C (clk), .D (signal_2655), .Q (signal_6507) ) ;
    buf_clk cell_4966 ( .C (clk), .D (signal_558), .Q (signal_6509) ) ;
    buf_clk cell_4968 ( .C (clk), .D (signal_2656), .Q (signal_6511) ) ;
    buf_clk cell_4970 ( .C (clk), .D (signal_562), .Q (signal_6513) ) ;
    buf_clk cell_4972 ( .C (clk), .D (signal_2657), .Q (signal_6515) ) ;
    buf_clk cell_4974 ( .C (clk), .D (signal_566), .Q (signal_6517) ) ;
    buf_clk cell_4976 ( .C (clk), .D (signal_2658), .Q (signal_6519) ) ;
    buf_clk cell_4978 ( .C (clk), .D (signal_570), .Q (signal_6521) ) ;
    buf_clk cell_4980 ( .C (clk), .D (signal_2659), .Q (signal_6523) ) ;
    buf_clk cell_4982 ( .C (clk), .D (signal_574), .Q (signal_6525) ) ;
    buf_clk cell_4984 ( .C (clk), .D (signal_2660), .Q (signal_6527) ) ;
    buf_clk cell_4986 ( .C (clk), .D (signal_578), .Q (signal_6529) ) ;
    buf_clk cell_4988 ( .C (clk), .D (signal_2661), .Q (signal_6531) ) ;
    buf_clk cell_4990 ( .C (clk), .D (signal_582), .Q (signal_6533) ) ;
    buf_clk cell_4992 ( .C (clk), .D (signal_2662), .Q (signal_6535) ) ;
    buf_clk cell_4994 ( .C (clk), .D (signal_586), .Q (signal_6537) ) ;
    buf_clk cell_4996 ( .C (clk), .D (signal_2663), .Q (signal_6539) ) ;

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_90 ( .a ({signal_4664, signal_4656}), .b ({signal_2351, signal_1303}), .c ({DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_92 ( .a ({signal_4680, signal_4672}), .b ({signal_2347, signal_1265}), .c ({DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_94 ( .a ({signal_4696, signal_4688}), .b ({signal_2335, signal_1249}), .c ({DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_96 ( .a ({signal_4712, signal_4704}), .b ({signal_2341, signal_1251}), .c ({DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_99 ( .a ({signal_4728, signal_4720}), .b ({signal_2350, signal_1277}), .c ({DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_101 ( .a ({signal_4744, signal_4736}), .b ({signal_2336, signal_1279}), .c ({DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_103 ( .a ({signal_4760, signal_4752}), .b ({signal_2343, signal_1305}), .c ({DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_105 ( .a ({signal_4776, signal_4768}), .b ({signal_2352, signal_1307}), .c ({DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_107 ( .a ({signal_4792, signal_4784}), .b ({signal_2334, signal_1285}), .c ({DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_108 ( .a ({signal_4808, signal_4800}), .b ({signal_2339, signal_1267}), .c ({DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_110 ( .a ({signal_4824, signal_4816}), .b ({signal_2342, signal_1287}), .c ({DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_112 ( .a ({signal_4840, signal_4832}), .b ({signal_2346, signal_1269}), .c ({DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_114 ( .a ({signal_4856, signal_4848}), .b ({signal_2344, signal_1271}), .c ({DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_116 ( .a ({signal_4872, signal_4864}), .b ({signal_2349, signal_1257}), .c ({DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_118 ( .a ({signal_4888, signal_4880}), .b ({signal_2348, signal_1259}), .c ({DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_121 ( .a ({signal_4904, signal_4896}), .b ({signal_2345, signal_1293}), .c ({DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_123 ( .a ({signal_4920, signal_4912}), .b ({signal_2338, signal_1295}), .c ({DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_125 ( .a ({signal_4936, signal_4928}), .b ({signal_2337, signal_1297}), .c ({DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_127 ( .a ({signal_4952, signal_4944}), .b ({signal_2340, signal_1299}), .c ({DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_129 ( .a ({signal_4968, signal_4960}), .b ({signal_2353, signal_1309}), .c ({DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_130 ( .a ({signal_4984, signal_4976}), .b ({signal_2354, signal_1261}), .c ({DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_132 ( .a ({signal_5000, signal_4992}), .b ({signal_2355, signal_1311}), .c ({DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_134 ( .a ({signal_5016, signal_5008}), .b ({signal_2356, signal_1281}), .c ({DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_136 ( .a ({signal_5032, signal_5024}), .b ({signal_2357, signal_1283}), .c ({DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_138 ( .a ({signal_5048, signal_5040}), .b ({signal_2358, signal_1253}), .c ({DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_140 ( .a ({signal_5064, signal_5056}), .b ({signal_2359, signal_1255}), .c ({DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_143 ( .a ({signal_5080, signal_5072}), .b ({signal_2360, signal_1273}), .c ({DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_145 ( .a ({signal_5096, signal_5088}), .b ({signal_2361, signal_1275}), .c ({DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_147 ( .a ({signal_5112, signal_5104}), .b ({signal_2362, signal_1289}), .c ({DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_149 ( .a ({signal_5128, signal_5120}), .b ({signal_2363, signal_1291}), .c ({DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_151 ( .a ({signal_5144, signal_5136}), .b ({signal_2364, signal_1301}), .c ({DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_152 ( .a ({signal_5160, signal_5152}), .b ({signal_2365, signal_1263}), .c ({DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .a ({signal_2351, signal_1303}), .b ({signal_5176, signal_5168}), .c ({signal_2618, signal_1239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .a ({signal_5192, signal_5184}), .b ({signal_2347, signal_1265}), .c ({signal_2398, signal_1241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_222 ( .a ({signal_5208, signal_5200}), .b ({signal_2335, signal_1249}), .c ({signal_2399, signal_1185}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_224 ( .a ({signal_2341, signal_1251}), .b ({signal_5224, signal_5216}), .c ({signal_2680, signal_1187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .a ({signal_5240, signal_5232}), .b ({signal_2350, signal_1277}), .c ({signal_2400, signal_1189}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .a ({signal_2336, signal_1279}), .b ({signal_5256, signal_5248}), .c ({signal_2681, signal_1191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .a ({signal_5272, signal_5264}), .b ({signal_2343, signal_1305}), .c ({signal_2401, signal_1193}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_233 ( .a ({signal_2352, signal_1307}), .b ({signal_5288, signal_5280}), .c ({signal_2682, signal_1195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({signal_5304, signal_5296}), .b ({signal_2334, signal_1285}), .c ({signal_2402, signal_1197}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({signal_2339, signal_1267}), .b ({signal_5320, signal_5312}), .c ({signal_2683, signal_1243}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({signal_2342, signal_1287}), .b ({signal_5336, signal_5328}), .c ({signal_2723, signal_1199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({signal_5352, signal_5344}), .b ({signal_2346, signal_1269}), .c ({signal_2403, signal_1201}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({signal_2344, signal_1271}), .b ({signal_5368, signal_5360}), .c ({signal_2619, signal_1203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({signal_5384, signal_5376}), .b ({signal_2349, signal_1257}), .c ({signal_2404, signal_1205}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({signal_2348, signal_1259}), .b ({signal_5400, signal_5392}), .c ({signal_2684, signal_1207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({signal_5416, signal_5408}), .b ({signal_2345, signal_1293}), .c ({signal_2405, signal_1209}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({signal_2338, signal_1295}), .b ({signal_5432, signal_5424}), .c ({signal_2620, signal_1211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({signal_5448, signal_5440}), .b ({signal_2337, signal_1297}), .c ({signal_2406, signal_1213}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({signal_2340, signal_1299}), .b ({signal_5464, signal_5456}), .c ({signal_2685, signal_1215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .a ({signal_5480, signal_5472}), .b ({signal_2353, signal_1309}), .c ({signal_2407, signal_1217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .a ({signal_5496, signal_5488}), .b ({signal_2354, signal_1261}), .c ({signal_2408, signal_1245}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .a ({signal_2355, signal_1311}), .b ({signal_5512, signal_5504}), .c ({signal_2711, signal_1219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({signal_5528, signal_5520}), .b ({signal_2356, signal_1281}), .c ({signal_2409, signal_1221}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({signal_2357, signal_1283}), .b ({signal_5544, signal_5536}), .c ({signal_2686, signal_1223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .a ({signal_5560, signal_5552}), .b ({signal_2358, signal_1253}), .c ({signal_2410, signal_1225}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .a ({signal_2359, signal_1255}), .b ({signal_5576, signal_5568}), .c ({signal_2621, signal_1227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({signal_5592, signal_5584}), .b ({signal_2360, signal_1273}), .c ({signal_2411, signal_1229}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({signal_2361, signal_1275}), .b ({signal_5608, signal_5600}), .c ({signal_2687, signal_1231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({signal_5624, signal_5616}), .b ({signal_2362, signal_1289}), .c ({signal_2412, signal_1233}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({signal_2363, signal_1291}), .b ({signal_5640, signal_5632}), .c ({signal_2688, signal_1235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .a ({signal_5656, signal_5648}), .b ({signal_2364, signal_1301}), .c ({signal_2413, signal_1237}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .a ({signal_2365, signal_1263}), .b ({signal_5672, signal_5664}), .c ({signal_2689, signal_1247}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .a ({signal_2740, signal_1111}), .b ({signal_5176, signal_5168}), .c ({signal_2744, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .a ({signal_5192, signal_5184}), .b ({signal_2562, signal_1065}), .c ({signal_2567, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .a ({signal_5208, signal_5200}), .b ({signal_2552, signal_1057}), .c ({signal_2568, signal_993}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .a ({signal_2763, signal_1059}), .b ({signal_5224, signal_5216}), .c ({signal_2775, signal_995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .a ({signal_5240, signal_5232}), .b ({signal_2553, signal_1097}), .c ({signal_2569, signal_997}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .a ({signal_2762, signal_1099}), .b ({signal_5256, signal_5248}), .c ({signal_2776, signal_999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .a ({signal_5272, signal_5264}), .b ({signal_2550, signal_1077}), .c ({signal_2570, signal_1001}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_300 ( .a ({signal_2755, signal_1079}), .b ({signal_5288, signal_5280}), .c ({signal_2759, signal_1003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_303 ( .a ({signal_5304, signal_5296}), .b ({signal_2551, signal_1117}), .c ({signal_2571, signal_1005}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_304 ( .a ({signal_2741, signal_1067}), .b ({signal_5320, signal_5312}), .c ({signal_2745, signal_1051}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_307 ( .a ({signal_2732, signal_1119}), .b ({signal_5336, signal_5328}), .c ({signal_2746, signal_1007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_310 ( .a ({signal_5352, signal_5344}), .b ({signal_2556, signal_1113}), .c ({signal_2572, signal_1009}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_312 ( .a ({signal_2735, signal_1115}), .b ({signal_5368, signal_5360}), .c ({signal_2747, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_315 ( .a ({signal_5384, signal_5376}), .b ({signal_2557, signal_1073}), .c ({signal_2574, signal_1013}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_317 ( .a ({signal_2733, signal_1075}), .b ({signal_5400, signal_5392}), .c ({signal_2748, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_321 ( .a ({signal_5416, signal_5408}), .b ({signal_2554, signal_1101}), .c ({signal_2575, signal_1017}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_323 ( .a ({signal_2734, signal_1103}), .b ({signal_5432, signal_5424}), .c ({signal_2749, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_326 ( .a ({signal_5448, signal_5440}), .b ({signal_2555, signal_1061}), .c ({signal_2577, signal_1021}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_328 ( .a ({signal_2736, signal_1063}), .b ({signal_5464, signal_5456}), .c ({signal_2750, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_331 ( .a ({signal_5480, signal_5472}), .b ({signal_2560, signal_1093}), .c ({signal_2578, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_332 ( .a ({signal_5496, signal_5488}), .b ({signal_2563, signal_1089}), .c ({signal_2579, signal_1053}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_334 ( .a ({signal_2738, signal_1095}), .b ({signal_5512, signal_5504}), .c ({signal_2751, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_337 ( .a ({signal_5528, signal_5520}), .b ({signal_2561, signal_1069}), .c ({signal_2580, signal_1029}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_339 ( .a ({signal_2737, signal_1071}), .b ({signal_5544, signal_5536}), .c ({signal_2752, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_342 ( .a ({signal_5560, signal_5552}), .b ({signal_2558, signal_1105}), .c ({signal_2581, signal_1033}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_344 ( .a ({signal_2757, signal_1107}), .b ({signal_5576, signal_5568}), .c ({signal_2760, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_348 ( .a ({signal_5592, signal_5584}), .b ({signal_2559, signal_1081}), .c ({signal_2583, signal_1037}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_350 ( .a ({signal_2758, signal_1083}), .b ({signal_5608, signal_5600}), .c ({signal_2761, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_353 ( .a ({signal_5624, signal_5616}), .b ({signal_2564, signal_1085}), .c ({signal_2584, signal_1041}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_355 ( .a ({signal_2742, signal_1087}), .b ({signal_5640, signal_5632}), .c ({signal_2753, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_358 ( .a ({signal_5656, signal_5648}), .b ({signal_2565, signal_1109}), .c ({signal_2585, signal_1045}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_359 ( .a ({signal_2743, signal_1091}), .b ({signal_5672, signal_5664}), .c ({signal_2754, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_535 ( .s (signal_5674), .b ({signal_2764, signal_1439}), .a ({signal_5690, signal_5682}), .c ({signal_2777, signal_460}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_541 ( .s (signal_5674), .b ({signal_2664, signal_1437}), .a ({signal_5706, signal_5698}), .c ({signal_2691, signal_464}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_547 ( .s (signal_5674), .b ({signal_2765, signal_1435}), .a ({signal_5722, signal_5714}), .c ({signal_2778, signal_468}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_553 ( .s (signal_5674), .b ({signal_2665, signal_1433}), .a ({signal_5738, signal_5730}), .c ({signal_2692, signal_472}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_559 ( .s (signal_5674), .b ({signal_2766, signal_1431}), .a ({signal_5754, signal_5746}), .c ({signal_2779, signal_476}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_565 ( .s (signal_5674), .b ({signal_2666, signal_1429}), .a ({signal_5770, signal_5762}), .c ({signal_2693, signal_480}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_571 ( .s (signal_5674), .b ({signal_2767, signal_1427}), .a ({signal_5786, signal_5778}), .c ({signal_2780, signal_484}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_577 ( .s (signal_5674), .b ({signal_2667, signal_1425}), .a ({signal_5802, signal_5794}), .c ({signal_2694, signal_488}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_583 ( .s (signal_5674), .b ({signal_2788, signal_1423}), .a ({signal_5818, signal_5810}), .c ({signal_2791, signal_492}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_589 ( .s (signal_5674), .b ({signal_2668, signal_1421}), .a ({signal_5834, signal_5826}), .c ({signal_2695, signal_496}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_595 ( .s (signal_5674), .b ({signal_2789, signal_1419}), .a ({signal_5850, signal_5842}), .c ({signal_2792, signal_500}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_601 ( .s (signal_5674), .b ({signal_2669, signal_1417}), .a ({signal_5866, signal_5858}), .c ({signal_2696, signal_504}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_607 ( .s (signal_5674), .b ({signal_2768, signal_1415}), .a ({signal_5882, signal_5874}), .c ({signal_2781, signal_508}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_613 ( .s (signal_5674), .b ({signal_2670, signal_1413}), .a ({signal_5898, signal_5890}), .c ({signal_2697, signal_512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_619 ( .s (signal_5674), .b ({signal_2769, signal_1411}), .a ({signal_5914, signal_5906}), .c ({signal_2782, signal_516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_625 ( .s (signal_5674), .b ({signal_2671, signal_1409}), .a ({signal_5930, signal_5922}), .c ({signal_2698, signal_520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_631 ( .s (signal_5674), .b ({signal_2770, signal_1407}), .a ({signal_5946, signal_5938}), .c ({signal_2783, signal_524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_637 ( .s (signal_5674), .b ({signal_2672, signal_1405}), .a ({signal_5962, signal_5954}), .c ({signal_2699, signal_528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_643 ( .s (signal_5674), .b ({signal_2771, signal_1403}), .a ({signal_5978, signal_5970}), .c ({signal_2784, signal_532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_649 ( .s (signal_5674), .b ({signal_2673, signal_1401}), .a ({signal_5994, signal_5986}), .c ({signal_2700, signal_536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_655 ( .s (signal_5674), .b ({signal_2772, signal_1399}), .a ({signal_6010, signal_6002}), .c ({signal_2785, signal_540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_661 ( .s (signal_5674), .b ({signal_2674, signal_1397}), .a ({signal_6026, signal_6018}), .c ({signal_2701, signal_544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_667 ( .s (signal_5674), .b ({signal_2773, signal_1395}), .a ({signal_6042, signal_6034}), .c ({signal_2786, signal_548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_673 ( .s (signal_5674), .b ({signal_2675, signal_1393}), .a ({signal_6058, signal_6050}), .c ({signal_2702, signal_552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_679 ( .s (signal_5674), .b ({signal_2774, signal_1391}), .a ({signal_6074, signal_6066}), .c ({signal_2787, signal_556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_685 ( .s (signal_5674), .b ({signal_2676, signal_1389}), .a ({signal_6090, signal_6082}), .c ({signal_2703, signal_560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_691 ( .s (signal_5674), .b ({signal_2790, signal_1387}), .a ({signal_6106, signal_6098}), .c ({signal_2793, signal_564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_697 ( .s (signal_5674), .b ({signal_2677, signal_1385}), .a ({signal_6122, signal_6114}), .c ({signal_2704, signal_568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_703 ( .s (signal_5674), .b ({signal_2794, signal_1383}), .a ({signal_6138, signal_6130}), .c ({signal_2796, signal_572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_709 ( .s (signal_5674), .b ({signal_2678, signal_1381}), .a ({signal_6154, signal_6146}), .c ({signal_2705, signal_576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_715 ( .s (signal_5674), .b ({signal_2795, signal_1379}), .a ({signal_6170, signal_6162}), .c ({signal_2797, signal_580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_721 ( .s (signal_5674), .b ({signal_2679, signal_1377}), .a ({signal_6186, signal_6178}), .c ({signal_2706, signal_584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .s (signal_6188), .b ({signal_2355, signal_1311}), .a ({signal_2689, signal_1247}), .c ({signal_2713, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .s (signal_6188), .b ({signal_2353, signal_1309}), .a ({signal_2408, signal_1245}), .c ({signal_2446, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .s (signal_6188), .b ({signal_2352, signal_1307}), .a ({signal_2683, signal_1243}), .c ({signal_2714, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .s (signal_6188), .b ({signal_2343, signal_1305}), .a ({signal_2398, signal_1241}), .c ({signal_2447, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .s (signal_6188), .b ({signal_2351, signal_1303}), .a ({signal_2618, signal_1239}), .c ({signal_2707, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .s (signal_6188), .b ({signal_2364, signal_1301}), .a ({signal_2413, signal_1237}), .c ({signal_2448, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .s (signal_6188), .b ({signal_2340, signal_1299}), .a ({signal_2688, signal_1235}), .c ({signal_2715, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .s (signal_6188), .b ({signal_2337, signal_1297}), .a ({signal_2412, signal_1233}), .c ({signal_2449, signal_1169}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .s (signal_6188), .b ({signal_2338, signal_1295}), .a ({signal_2687, signal_1231}), .c ({signal_2716, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .s (signal_6188), .b ({signal_2345, signal_1293}), .a ({signal_2411, signal_1229}), .c ({signal_2450, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .s (signal_6188), .b ({signal_2363, signal_1291}), .a ({signal_2621, signal_1227}), .c ({signal_2708, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1053 ( .s (signal_6188), .b ({signal_2362, signal_1289}), .a ({signal_2410, signal_1225}), .c ({signal_2451, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1055 ( .s (signal_6188), .b ({signal_2342, signal_1287}), .a ({signal_2686, signal_1223}), .c ({signal_2717, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1057 ( .s (signal_6188), .b ({signal_2334, signal_1285}), .a ({signal_2409, signal_1221}), .c ({signal_2452, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1059 ( .s (signal_6188), .b ({signal_2357, signal_1283}), .a ({signal_2711, signal_1219}), .c ({signal_2724, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1061 ( .s (signal_6188), .b ({signal_2356, signal_1281}), .a ({signal_2407, signal_1217}), .c ({signal_2453, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1063 ( .s (signal_6188), .b ({signal_2336, signal_1279}), .a ({signal_2685, signal_1215}), .c ({signal_2718, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1065 ( .s (signal_6188), .b ({signal_2350, signal_1277}), .a ({signal_2406, signal_1213}), .c ({signal_2454, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1067 ( .s (signal_6188), .b ({signal_2361, signal_1275}), .a ({signal_2620, signal_1211}), .c ({signal_2709, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1069 ( .s (signal_6188), .b ({signal_2360, signal_1273}), .a ({signal_2405, signal_1209}), .c ({signal_2455, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1071 ( .s (signal_6188), .b ({signal_2344, signal_1271}), .a ({signal_2684, signal_1207}), .c ({signal_2719, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1073 ( .s (signal_6188), .b ({signal_2346, signal_1269}), .a ({signal_2404, signal_1205}), .c ({signal_2456, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1075 ( .s (signal_6188), .b ({signal_2339, signal_1267}), .a ({signal_2619, signal_1203}), .c ({signal_2710, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1077 ( .s (signal_6188), .b ({signal_2347, signal_1265}), .a ({signal_2403, signal_1201}), .c ({signal_2457, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1079 ( .s (signal_6188), .b ({signal_2365, signal_1263}), .a ({signal_2723, signal_1199}), .c ({signal_2731, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1081 ( .s (signal_6188), .b ({signal_2354, signal_1261}), .a ({signal_2402, signal_1197}), .c ({signal_2458, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1083 ( .s (signal_6188), .b ({signal_2348, signal_1259}), .a ({signal_2682, signal_1195}), .c ({signal_2720, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1085 ( .s (signal_6188), .b ({signal_2349, signal_1257}), .a ({signal_2401, signal_1193}), .c ({signal_2459, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1087 ( .s (signal_6188), .b ({signal_2359, signal_1255}), .a ({signal_2681, signal_1191}), .c ({signal_2721, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1089 ( .s (signal_6188), .b ({signal_2358, signal_1253}), .a ({signal_2400, signal_1189}), .c ({signal_2460, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1091 ( .s (signal_6188), .b ({signal_2341, signal_1251}), .a ({signal_2680, signal_1187}), .c ({signal_2722, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1093 ( .s (signal_6188), .b ({signal_2335, signal_1249}), .a ({signal_2399, signal_1185}), .c ({signal_2461, signal_1121}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1096 ( .a ({signal_2722, signal_1123}), .b ({signal_2756, signal_829}), .c ({signal_2762, signal_1099}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1098 ( .a ({signal_2458, signal_1133}), .b ({signal_2482, signal_831}), .c ({signal_2550, signal_1077}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1100 ( .a ({signal_2731, signal_1135}), .b ({signal_2725, signal_833}), .c ({signal_2755, signal_1079}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1103 ( .a ({signal_2459, signal_1129}), .b ({signal_2482, signal_831}), .c ({signal_2551, signal_1117}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1104 ( .a ({signal_2461, signal_1121}), .b ({signal_2460, signal_1125}), .c ({signal_2482, signal_831}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1108 ( .a ({signal_2460, signal_1125}), .b ({signal_2487, signal_835}), .c ({signal_2552, signal_1057}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1111 ( .a ({signal_2721, signal_1127}), .b ({signal_2756, signal_829}), .c ({signal_2763, signal_1059}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1112 ( .a ({signal_2720, signal_1131}), .b ({signal_2731, signal_1135}), .c ({signal_2756, signal_829}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1115 ( .a ({signal_2461, signal_1121}), .b ({signal_2487, signal_835}), .c ({signal_2553, signal_1097}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1116 ( .a ({signal_2458, signal_1133}), .b ({signal_2459, signal_1129}), .c ({signal_2487, signal_835}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1117 ( .a ({signal_2720, signal_1131}), .b ({signal_2725, signal_833}), .c ({signal_2732, signal_1119}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1118 ( .a ({signal_2722, signal_1123}), .b ({signal_2721, signal_1127}), .c ({signal_2725, signal_833}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1120 ( .a ({signal_2710, signal_1139}), .b ({signal_2726, signal_837}), .c ({signal_2733, signal_1075}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1122 ( .a ({signal_2454, signal_1149}), .b ({signal_2492, signal_839}), .c ({signal_2554, signal_1101}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1124 ( .a ({signal_2718, signal_1151}), .b ({signal_2727, signal_841}), .c ({signal_2734, signal_1103}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1127 ( .a ({signal_2455, signal_1145}), .b ({signal_2492, signal_839}), .c ({signal_2555, signal_1061}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1128 ( .a ({signal_2457, signal_1137}), .b ({signal_2456, signal_1141}), .c ({signal_2492, signal_839}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1132 ( .a ({signal_2456, signal_1141}), .b ({signal_2497, signal_843}), .c ({signal_2556, signal_1113}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1135 ( .a ({signal_2719, signal_1143}), .b ({signal_2726, signal_837}), .c ({signal_2735, signal_1115}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1136 ( .a ({signal_2709, signal_1147}), .b ({signal_2718, signal_1151}), .c ({signal_2726, signal_837}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1139 ( .a ({signal_2457, signal_1137}), .b ({signal_2497, signal_843}), .c ({signal_2557, signal_1073}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1140 ( .a ({signal_2454, signal_1149}), .b ({signal_2455, signal_1145}), .c ({signal_2497, signal_843}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1141 ( .a ({signal_2709, signal_1147}), .b ({signal_2727, signal_841}), .c ({signal_2736, signal_1063}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1142 ( .a ({signal_2710, signal_1139}), .b ({signal_2719, signal_1143}), .c ({signal_2727, signal_841}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1144 ( .a ({signal_2724, signal_1155}), .b ({signal_2728, signal_845}), .c ({signal_2737, signal_1071}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1146 ( .a ({signal_2450, signal_1165}), .b ({signal_2502, signal_847}), .c ({signal_2558, signal_1105}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1148 ( .a ({signal_2716, signal_1167}), .b ({signal_2739, signal_849}), .c ({signal_2757, signal_1107}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1151 ( .a ({signal_2451, signal_1161}), .b ({signal_2502, signal_847}), .c ({signal_2559, signal_1081}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1152 ( .a ({signal_2453, signal_1153}), .b ({signal_2452, signal_1157}), .c ({signal_2502, signal_847}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1156 ( .a ({signal_2452, signal_1157}), .b ({signal_2507, signal_851}), .c ({signal_2560, signal_1093}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1159 ( .a ({signal_2717, signal_1159}), .b ({signal_2728, signal_845}), .c ({signal_2738, signal_1095}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1160 ( .a ({signal_2708, signal_1163}), .b ({signal_2716, signal_1167}), .c ({signal_2728, signal_845}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1163 ( .a ({signal_2453, signal_1153}), .b ({signal_2507, signal_851}), .c ({signal_2561, signal_1069}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1164 ( .a ({signal_2450, signal_1165}), .b ({signal_2451, signal_1161}), .c ({signal_2507, signal_851}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1165 ( .a ({signal_2708, signal_1163}), .b ({signal_2739, signal_849}), .c ({signal_2758, signal_1083}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1166 ( .a ({signal_2724, signal_1155}), .b ({signal_2717, signal_1159}), .c ({signal_2739, signal_849}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1168 ( .a ({signal_2715, signal_1171}), .b ({signal_2729, signal_853}), .c ({signal_2740, signal_1111}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1170 ( .a ({signal_2446, signal_1181}), .b ({signal_2512, signal_855}), .c ({signal_2562, signal_1065}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1172 ( .a ({signal_2713, signal_1183}), .b ({signal_2730, signal_857}), .c ({signal_2741, signal_1067}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1175 ( .a ({signal_2447, signal_1177}), .b ({signal_2512, signal_855}), .c ({signal_2563, signal_1089}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1176 ( .a ({signal_2449, signal_1169}), .b ({signal_2448, signal_1173}), .c ({signal_2512, signal_855}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1180 ( .a ({signal_2448, signal_1173}), .b ({signal_2517, signal_859}), .c ({signal_2564, signal_1085}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1183 ( .a ({signal_2707, signal_1175}), .b ({signal_2729, signal_853}), .c ({signal_2742, signal_1087}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1184 ( .a ({signal_2714, signal_1179}), .b ({signal_2713, signal_1183}), .c ({signal_2729, signal_853}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1187 ( .a ({signal_2449, signal_1169}), .b ({signal_2517, signal_859}), .c ({signal_2565, signal_1109}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1188 ( .a ({signal_2446, signal_1181}), .b ({signal_2447, signal_1177}), .c ({signal_2517, signal_859}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1189 ( .a ({signal_2714, signal_1179}), .b ({signal_2730, signal_857}), .c ({signal_2743, signal_1091}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1190 ( .a ({signal_2715, signal_1171}), .b ({signal_2707, signal_1175}), .c ({signal_2730, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1191 ( .s (signal_6188), .b ({signal_2754, signal_1055}), .a ({signal_2732, signal_1119}), .c ({signal_2764, signal_1439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1193 ( .s (signal_6188), .b ({signal_2579, signal_1053}), .a ({signal_2551, signal_1117}), .c ({signal_2664, signal_1437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1195 ( .s (signal_6188), .b ({signal_2745, signal_1051}), .a ({signal_2735, signal_1115}), .c ({signal_2765, signal_1435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1197 ( .s (signal_6188), .b ({signal_2567, signal_1049}), .a ({signal_2556, signal_1113}), .c ({signal_2665, signal_1433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1199 ( .s (signal_6188), .b ({signal_2744, signal_1047}), .a ({signal_2740, signal_1111}), .c ({signal_2766, signal_1431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1201 ( .s (signal_6188), .b ({signal_2585, signal_1045}), .a ({signal_2565, signal_1109}), .c ({signal_2666, signal_1429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1203 ( .s (signal_6188), .b ({signal_2753, signal_1043}), .a ({signal_2757, signal_1107}), .c ({signal_2767, signal_1427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1205 ( .s (signal_6188), .b ({signal_2584, signal_1041}), .a ({signal_2558, signal_1105}), .c ({signal_2667, signal_1425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1207 ( .s (signal_6188), .b ({signal_2761, signal_1039}), .a ({signal_2734, signal_1103}), .c ({signal_2788, signal_1423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1209 ( .s (signal_6188), .b ({signal_2583, signal_1037}), .a ({signal_2554, signal_1101}), .c ({signal_2668, signal_1421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1211 ( .s (signal_6188), .b ({signal_2760, signal_1035}), .a ({signal_2762, signal_1099}), .c ({signal_2789, signal_1419}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1213 ( .s (signal_6188), .b ({signal_2581, signal_1033}), .a ({signal_2553, signal_1097}), .c ({signal_2669, signal_1417}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1215 ( .s (signal_6188), .b ({signal_2752, signal_1031}), .a ({signal_2738, signal_1095}), .c ({signal_2768, signal_1415}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1217 ( .s (signal_6188), .b ({signal_2580, signal_1029}), .a ({signal_2560, signal_1093}), .c ({signal_2670, signal_1413}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1219 ( .s (signal_6188), .b ({signal_2751, signal_1027}), .a ({signal_2743, signal_1091}), .c ({signal_2769, signal_1411}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1221 ( .s (signal_6188), .b ({signal_2578, signal_1025}), .a ({signal_2563, signal_1089}), .c ({signal_2671, signal_1409}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1223 ( .s (signal_6188), .b ({signal_2750, signal_1023}), .a ({signal_2742, signal_1087}), .c ({signal_2770, signal_1407}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1225 ( .s (signal_6188), .b ({signal_2577, signal_1021}), .a ({signal_2564, signal_1085}), .c ({signal_2672, signal_1405}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1227 ( .s (signal_6188), .b ({signal_2749, signal_1019}), .a ({signal_2758, signal_1083}), .c ({signal_2771, signal_1403}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1229 ( .s (signal_6188), .b ({signal_2575, signal_1017}), .a ({signal_2559, signal_1081}), .c ({signal_2673, signal_1401}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1231 ( .s (signal_6188), .b ({signal_2748, signal_1015}), .a ({signal_2755, signal_1079}), .c ({signal_2772, signal_1399}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1233 ( .s (signal_6188), .b ({signal_2574, signal_1013}), .a ({signal_2550, signal_1077}), .c ({signal_2674, signal_1397}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1235 ( .s (signal_6188), .b ({signal_2747, signal_1011}), .a ({signal_2733, signal_1075}), .c ({signal_2773, signal_1395}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1237 ( .s (signal_6188), .b ({signal_2572, signal_1009}), .a ({signal_2557, signal_1073}), .c ({signal_2675, signal_1393}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1239 ( .s (signal_6188), .b ({signal_2746, signal_1007}), .a ({signal_2737, signal_1071}), .c ({signal_2774, signal_1391}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1241 ( .s (signal_6188), .b ({signal_2571, signal_1005}), .a ({signal_2561, signal_1069}), .c ({signal_2676, signal_1389}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1243 ( .s (signal_6188), .b ({signal_2759, signal_1003}), .a ({signal_2741, signal_1067}), .c ({signal_2790, signal_1387}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1245 ( .s (signal_6188), .b ({signal_2570, signal_1001}), .a ({signal_2562, signal_1065}), .c ({signal_2677, signal_1385}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1247 ( .s (signal_6188), .b ({signal_2776, signal_999}), .a ({signal_2736, signal_1063}), .c ({signal_2794, signal_1383}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1249 ( .s (signal_6188), .b ({signal_2569, signal_997}), .a ({signal_2555, signal_1061}), .c ({signal_2678, signal_1381}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1251 ( .s (signal_6188), .b ({signal_2775, signal_995}), .a ({signal_2763, signal_1059}), .c ({signal_2795, signal_1379}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1253 ( .s (signal_6188), .b ({signal_2568, signal_993}), .a ({signal_2552, signal_1057}), .c ({signal_2679, signal_1377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .s ({signal_6192, signal_6190}), .b ({signal_6196, signal_6194}), .a ({signal_2215, signal_1602}), .clk (clk), .r (Fresh[199]), .c ({signal_2334, signal_1285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .s ({signal_6200, signal_6198}), .b ({signal_6204, signal_6202}), .a ({signal_2228, signal_1606}), .clk (clk), .r (Fresh[200]), .c ({signal_2335, signal_1249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .s ({signal_6208, signal_6206}), .b ({signal_2216, signal_1603}), .a ({signal_6212, signal_6210}), .clk (clk), .r (Fresh[201]), .c ({signal_2336, signal_1279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .s ({signal_6216, signal_6214}), .b ({signal_6220, signal_6218}), .a ({signal_2204, signal_1598}), .clk (clk), .r (Fresh[202]), .c ({signal_2337, signal_1297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .s ({signal_6224, signal_6222}), .b ({signal_2196, signal_1593}), .a ({signal_6228, signal_6226}), .clk (clk), .r (Fresh[203]), .c ({signal_2338, signal_1295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .s ({signal_6232, signal_6230}), .b ({signal_2213, signal_1600}), .a ({signal_6236, signal_6234}), .clk (clk), .r (Fresh[204]), .c ({signal_2339, signal_1267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .s ({signal_6216, signal_6214}), .b ({signal_2200, signal_1596}), .a ({signal_6240, signal_6238}), .clk (clk), .r (Fresh[205]), .c ({signal_2340, signal_1299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .s ({signal_6200, signal_6198}), .b ({signal_2198, signal_1595}), .a ({signal_6244, signal_6242}), .clk (clk), .r (Fresh[206]), .c ({signal_2341, signal_1251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .s ({signal_6192, signal_6190}), .b ({signal_2221, signal_1604}), .a ({signal_6248, signal_6246}), .clk (clk), .r (Fresh[207]), .c ({signal_2342, signal_1287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .s ({signal_6252, signal_6250}), .b ({signal_6256, signal_6254}), .a ({signal_2201, signal_1597}), .clk (clk), .r (Fresh[208]), .c ({signal_2343, signal_1305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .s ({signal_6260, signal_6258}), .b ({signal_2229, signal_1607}), .a ({signal_6264, signal_6262}), .clk (clk), .r (Fresh[209]), .c ({signal_2344, signal_1271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .s ({signal_6224, signal_6222}), .b ({signal_6268, signal_6266}), .a ({signal_2210, signal_1599}), .clk (clk), .r (Fresh[210]), .c ({signal_2345, signal_1293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .s ({signal_6260, signal_6258}), .b ({signal_6272, signal_6270}), .a ({signal_2222, signal_1605}), .clk (clk), .r (Fresh[211]), .c ({signal_2346, signal_1269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .s ({signal_6232, signal_6230}), .b ({signal_6276, signal_6274}), .a ({signal_2214, signal_1601}), .clk (clk), .r (Fresh[212]), .c ({signal_2347, signal_1265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .s ({signal_6280, signal_6278}), .b ({signal_2232, signal_1608}), .a ({signal_6284, signal_6282}), .clk (clk), .r (Fresh[213]), .c ({signal_2348, signal_1259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .s ({signal_6280, signal_6278}), .b ({signal_6288, signal_6286}), .a ({signal_2237, signal_1609}), .clk (clk), .r (Fresh[214]), .c ({signal_2349, signal_1257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .s ({signal_6208, signal_6206}), .b ({signal_6292, signal_6290}), .a ({signal_2197, signal_1594}), .clk (clk), .r (Fresh[215]), .c ({signal_2350, signal_1277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .s ({signal_6296, signal_6294}), .b ({signal_2193, signal_1591}), .a ({signal_6300, signal_6298}), .clk (clk), .r (Fresh[216]), .c ({signal_2351, signal_1303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .s ({signal_6252, signal_6250}), .b ({signal_2195, signal_1592}), .a ({signal_6304, signal_6302}), .clk (clk), .r (Fresh[217]), .c ({signal_2352, signal_1307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .s ({signal_6308, signal_6306}), .b ({signal_6312, signal_6310}), .a ({signal_2241, signal_1610}), .clk (clk), .r (Fresh[218]), .c ({signal_2353, signal_1309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .s ({signal_6316, signal_6314}), .b ({signal_6320, signal_6318}), .a ({signal_2242, signal_1611}), .clk (clk), .r (Fresh[219]), .c ({signal_2354, signal_1261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .s ({signal_6308, signal_6306}), .b ({signal_2244, signal_1612}), .a ({signal_6324, signal_6322}), .clk (clk), .r (Fresh[220]), .c ({signal_2355, signal_1311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .s ({signal_6328, signal_6326}), .b ({signal_6332, signal_6330}), .a ({signal_2247, signal_1613}), .clk (clk), .r (Fresh[221]), .c ({signal_2356, signal_1281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .s ({signal_6328, signal_6326}), .b ({signal_2249, signal_1614}), .a ({signal_6336, signal_6334}), .clk (clk), .r (Fresh[222]), .c ({signal_2357, signal_1283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .s ({signal_6340, signal_6338}), .b ({signal_6344, signal_6342}), .a ({signal_2252, signal_1615}), .clk (clk), .r (Fresh[223]), .c ({signal_2358, signal_1253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .s ({signal_6340, signal_6338}), .b ({signal_2254, signal_1616}), .a ({signal_6348, signal_6346}), .clk (clk), .r (Fresh[224]), .c ({signal_2359, signal_1255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .s ({signal_6352, signal_6350}), .b ({signal_6356, signal_6354}), .a ({signal_2258, signal_1617}), .clk (clk), .r (Fresh[225]), .c ({signal_2360, signal_1273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .s ({signal_6352, signal_6350}), .b ({signal_2260, signal_1618}), .a ({signal_6360, signal_6358}), .clk (clk), .r (Fresh[226]), .c ({signal_2361, signal_1275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .s ({signal_6364, signal_6362}), .b ({signal_6368, signal_6366}), .a ({signal_2263, signal_1619}), .clk (clk), .r (Fresh[227]), .c ({signal_2362, signal_1289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .s ({signal_6364, signal_6362}), .b ({signal_2265, signal_1620}), .a ({signal_6372, signal_6370}), .clk (clk), .r (Fresh[228]), .c ({signal_2363, signal_1291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .s ({signal_6296, signal_6294}), .b ({signal_6376, signal_6374}), .a ({signal_2268, signal_1621}), .clk (clk), .r (Fresh[229]), .c ({signal_2364, signal_1301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .s ({signal_6316, signal_6314}), .b ({signal_2269, signal_1622}), .a ({signal_6380, signal_6378}), .clk (clk), .r (Fresh[230]), .c ({signal_2365, signal_1263}) ) ;
    buf_clk cell_1487 ( .C (clk), .D (signal_3029), .Q (DataOut_s0[63]) ) ;
    buf_clk cell_1489 ( .C (clk), .D (signal_3031), .Q (DataOut_s0[61]) ) ;
    buf_clk cell_1491 ( .C (clk), .D (signal_3033), .Q (DataOut_s0[59]) ) ;
    buf_clk cell_1493 ( .C (clk), .D (signal_3035), .Q (DataOut_s0[57]) ) ;
    buf_clk cell_1495 ( .C (clk), .D (signal_3037), .Q (DataOut_s0[55]) ) ;
    buf_clk cell_1497 ( .C (clk), .D (signal_3039), .Q (DataOut_s0[53]) ) ;
    buf_clk cell_1499 ( .C (clk), .D (signal_3041), .Q (DataOut_s0[51]) ) ;
    buf_clk cell_1501 ( .C (clk), .D (signal_3043), .Q (DataOut_s0[49]) ) ;
    buf_clk cell_1503 ( .C (clk), .D (signal_3045), .Q (DataOut_s0[47]) ) ;
    buf_clk cell_1505 ( .C (clk), .D (signal_3047), .Q (DataOut_s0[45]) ) ;
    buf_clk cell_1507 ( .C (clk), .D (signal_3049), .Q (DataOut_s0[43]) ) ;
    buf_clk cell_1509 ( .C (clk), .D (signal_3051), .Q (DataOut_s0[41]) ) ;
    buf_clk cell_1511 ( .C (clk), .D (signal_3053), .Q (DataOut_s0[39]) ) ;
    buf_clk cell_1513 ( .C (clk), .D (signal_3055), .Q (DataOut_s0[37]) ) ;
    buf_clk cell_1515 ( .C (clk), .D (signal_3057), .Q (DataOut_s0[35]) ) ;
    buf_clk cell_1517 ( .C (clk), .D (signal_3059), .Q (DataOut_s0[33]) ) ;
    buf_clk cell_1519 ( .C (clk), .D (signal_3061), .Q (DataOut_s0[31]) ) ;
    buf_clk cell_1521 ( .C (clk), .D (signal_3063), .Q (DataOut_s0[29]) ) ;
    buf_clk cell_1523 ( .C (clk), .D (signal_3065), .Q (DataOut_s0[27]) ) ;
    buf_clk cell_1525 ( .C (clk), .D (signal_3067), .Q (DataOut_s0[25]) ) ;
    buf_clk cell_1527 ( .C (clk), .D (signal_3069), .Q (DataOut_s0[23]) ) ;
    buf_clk cell_1529 ( .C (clk), .D (signal_3071), .Q (DataOut_s0[21]) ) ;
    buf_clk cell_1531 ( .C (clk), .D (signal_3073), .Q (DataOut_s0[19]) ) ;
    buf_clk cell_1533 ( .C (clk), .D (signal_3075), .Q (DataOut_s0[17]) ) ;
    buf_clk cell_1535 ( .C (clk), .D (signal_3077), .Q (DataOut_s0[15]) ) ;
    buf_clk cell_1537 ( .C (clk), .D (signal_3079), .Q (DataOut_s0[13]) ) ;
    buf_clk cell_1539 ( .C (clk), .D (signal_3081), .Q (DataOut_s0[11]) ) ;
    buf_clk cell_1541 ( .C (clk), .D (signal_3083), .Q (DataOut_s0[9]) ) ;
    buf_clk cell_1543 ( .C (clk), .D (signal_3085), .Q (DataOut_s0[7]) ) ;
    buf_clk cell_1545 ( .C (clk), .D (signal_3087), .Q (DataOut_s0[5]) ) ;
    buf_clk cell_1547 ( .C (clk), .D (signal_3089), .Q (DataOut_s0[3]) ) ;
    buf_clk cell_1549 ( .C (clk), .D (signal_3091), .Q (DataOut_s0[1]) ) ;
    buf_clk cell_1557 ( .C (clk), .D (signal_3099), .Q (done) ) ;
    buf_clk cell_1559 ( .C (clk), .D (signal_3101), .Q (DataOut_s1[9]) ) ;
    buf_clk cell_1561 ( .C (clk), .D (signal_3103), .Q (DataOut_s1[7]) ) ;
    buf_clk cell_1563 ( .C (clk), .D (signal_3105), .Q (DataOut_s1[63]) ) ;
    buf_clk cell_1565 ( .C (clk), .D (signal_3107), .Q (DataOut_s1[61]) ) ;
    buf_clk cell_1567 ( .C (clk), .D (signal_3109), .Q (DataOut_s1[5]) ) ;
    buf_clk cell_1569 ( .C (clk), .D (signal_3111), .Q (DataOut_s1[59]) ) ;
    buf_clk cell_1571 ( .C (clk), .D (signal_3113), .Q (DataOut_s1[57]) ) ;
    buf_clk cell_1573 ( .C (clk), .D (signal_3115), .Q (DataOut_s1[55]) ) ;
    buf_clk cell_1575 ( .C (clk), .D (signal_3117), .Q (DataOut_s1[53]) ) ;
    buf_clk cell_1577 ( .C (clk), .D (signal_3119), .Q (DataOut_s1[51]) ) ;
    buf_clk cell_1579 ( .C (clk), .D (signal_3121), .Q (DataOut_s1[49]) ) ;
    buf_clk cell_1581 ( .C (clk), .D (signal_3123), .Q (DataOut_s1[47]) ) ;
    buf_clk cell_1583 ( .C (clk), .D (signal_3125), .Q (DataOut_s1[45]) ) ;
    buf_clk cell_1585 ( .C (clk), .D (signal_3127), .Q (DataOut_s1[43]) ) ;
    buf_clk cell_1587 ( .C (clk), .D (signal_3129), .Q (DataOut_s1[41]) ) ;
    buf_clk cell_1589 ( .C (clk), .D (signal_3131), .Q (DataOut_s1[3]) ) ;
    buf_clk cell_1591 ( .C (clk), .D (signal_3133), .Q (DataOut_s1[39]) ) ;
    buf_clk cell_1593 ( .C (clk), .D (signal_3135), .Q (DataOut_s1[37]) ) ;
    buf_clk cell_1595 ( .C (clk), .D (signal_3137), .Q (DataOut_s1[35]) ) ;
    buf_clk cell_1597 ( .C (clk), .D (signal_3139), .Q (DataOut_s1[33]) ) ;
    buf_clk cell_1599 ( .C (clk), .D (signal_3141), .Q (DataOut_s1[31]) ) ;
    buf_clk cell_1601 ( .C (clk), .D (signal_3143), .Q (DataOut_s1[29]) ) ;
    buf_clk cell_1603 ( .C (clk), .D (signal_3145), .Q (DataOut_s1[27]) ) ;
    buf_clk cell_1605 ( .C (clk), .D (signal_3147), .Q (DataOut_s1[25]) ) ;
    buf_clk cell_1607 ( .C (clk), .D (signal_3149), .Q (DataOut_s1[23]) ) ;
    buf_clk cell_1609 ( .C (clk), .D (signal_3151), .Q (DataOut_s1[21]) ) ;
    buf_clk cell_1611 ( .C (clk), .D (signal_3153), .Q (DataOut_s1[1]) ) ;
    buf_clk cell_1613 ( .C (clk), .D (signal_3155), .Q (DataOut_s1[19]) ) ;
    buf_clk cell_1615 ( .C (clk), .D (signal_3157), .Q (DataOut_s1[17]) ) ;
    buf_clk cell_1617 ( .C (clk), .D (signal_3159), .Q (DataOut_s1[15]) ) ;
    buf_clk cell_1619 ( .C (clk), .D (signal_3161), .Q (DataOut_s1[13]) ) ;
    buf_clk cell_1621 ( .C (clk), .D (signal_3163), .Q (DataOut_s1[11]) ) ;
    buf_clk cell_3113 ( .C (clk), .D (signal_4655), .Q (signal_4656) ) ;
    buf_clk cell_3121 ( .C (clk), .D (signal_4663), .Q (signal_4664) ) ;
    buf_clk cell_3129 ( .C (clk), .D (signal_4671), .Q (signal_4672) ) ;
    buf_clk cell_3137 ( .C (clk), .D (signal_4679), .Q (signal_4680) ) ;
    buf_clk cell_3145 ( .C (clk), .D (signal_4687), .Q (signal_4688) ) ;
    buf_clk cell_3153 ( .C (clk), .D (signal_4695), .Q (signal_4696) ) ;
    buf_clk cell_3161 ( .C (clk), .D (signal_4703), .Q (signal_4704) ) ;
    buf_clk cell_3169 ( .C (clk), .D (signal_4711), .Q (signal_4712) ) ;
    buf_clk cell_3177 ( .C (clk), .D (signal_4719), .Q (signal_4720) ) ;
    buf_clk cell_3185 ( .C (clk), .D (signal_4727), .Q (signal_4728) ) ;
    buf_clk cell_3193 ( .C (clk), .D (signal_4735), .Q (signal_4736) ) ;
    buf_clk cell_3201 ( .C (clk), .D (signal_4743), .Q (signal_4744) ) ;
    buf_clk cell_3209 ( .C (clk), .D (signal_4751), .Q (signal_4752) ) ;
    buf_clk cell_3217 ( .C (clk), .D (signal_4759), .Q (signal_4760) ) ;
    buf_clk cell_3225 ( .C (clk), .D (signal_4767), .Q (signal_4768) ) ;
    buf_clk cell_3233 ( .C (clk), .D (signal_4775), .Q (signal_4776) ) ;
    buf_clk cell_3241 ( .C (clk), .D (signal_4783), .Q (signal_4784) ) ;
    buf_clk cell_3249 ( .C (clk), .D (signal_4791), .Q (signal_4792) ) ;
    buf_clk cell_3257 ( .C (clk), .D (signal_4799), .Q (signal_4800) ) ;
    buf_clk cell_3265 ( .C (clk), .D (signal_4807), .Q (signal_4808) ) ;
    buf_clk cell_3273 ( .C (clk), .D (signal_4815), .Q (signal_4816) ) ;
    buf_clk cell_3281 ( .C (clk), .D (signal_4823), .Q (signal_4824) ) ;
    buf_clk cell_3289 ( .C (clk), .D (signal_4831), .Q (signal_4832) ) ;
    buf_clk cell_3297 ( .C (clk), .D (signal_4839), .Q (signal_4840) ) ;
    buf_clk cell_3305 ( .C (clk), .D (signal_4847), .Q (signal_4848) ) ;
    buf_clk cell_3313 ( .C (clk), .D (signal_4855), .Q (signal_4856) ) ;
    buf_clk cell_3321 ( .C (clk), .D (signal_4863), .Q (signal_4864) ) ;
    buf_clk cell_3329 ( .C (clk), .D (signal_4871), .Q (signal_4872) ) ;
    buf_clk cell_3337 ( .C (clk), .D (signal_4879), .Q (signal_4880) ) ;
    buf_clk cell_3345 ( .C (clk), .D (signal_4887), .Q (signal_4888) ) ;
    buf_clk cell_3353 ( .C (clk), .D (signal_4895), .Q (signal_4896) ) ;
    buf_clk cell_3361 ( .C (clk), .D (signal_4903), .Q (signal_4904) ) ;
    buf_clk cell_3369 ( .C (clk), .D (signal_4911), .Q (signal_4912) ) ;
    buf_clk cell_3377 ( .C (clk), .D (signal_4919), .Q (signal_4920) ) ;
    buf_clk cell_3385 ( .C (clk), .D (signal_4927), .Q (signal_4928) ) ;
    buf_clk cell_3393 ( .C (clk), .D (signal_4935), .Q (signal_4936) ) ;
    buf_clk cell_3401 ( .C (clk), .D (signal_4943), .Q (signal_4944) ) ;
    buf_clk cell_3409 ( .C (clk), .D (signal_4951), .Q (signal_4952) ) ;
    buf_clk cell_3417 ( .C (clk), .D (signal_4959), .Q (signal_4960) ) ;
    buf_clk cell_3425 ( .C (clk), .D (signal_4967), .Q (signal_4968) ) ;
    buf_clk cell_3433 ( .C (clk), .D (signal_4975), .Q (signal_4976) ) ;
    buf_clk cell_3441 ( .C (clk), .D (signal_4983), .Q (signal_4984) ) ;
    buf_clk cell_3449 ( .C (clk), .D (signal_4991), .Q (signal_4992) ) ;
    buf_clk cell_3457 ( .C (clk), .D (signal_4999), .Q (signal_5000) ) ;
    buf_clk cell_3465 ( .C (clk), .D (signal_5007), .Q (signal_5008) ) ;
    buf_clk cell_3473 ( .C (clk), .D (signal_5015), .Q (signal_5016) ) ;
    buf_clk cell_3481 ( .C (clk), .D (signal_5023), .Q (signal_5024) ) ;
    buf_clk cell_3489 ( .C (clk), .D (signal_5031), .Q (signal_5032) ) ;
    buf_clk cell_3497 ( .C (clk), .D (signal_5039), .Q (signal_5040) ) ;
    buf_clk cell_3505 ( .C (clk), .D (signal_5047), .Q (signal_5048) ) ;
    buf_clk cell_3513 ( .C (clk), .D (signal_5055), .Q (signal_5056) ) ;
    buf_clk cell_3521 ( .C (clk), .D (signal_5063), .Q (signal_5064) ) ;
    buf_clk cell_3529 ( .C (clk), .D (signal_5071), .Q (signal_5072) ) ;
    buf_clk cell_3537 ( .C (clk), .D (signal_5079), .Q (signal_5080) ) ;
    buf_clk cell_3545 ( .C (clk), .D (signal_5087), .Q (signal_5088) ) ;
    buf_clk cell_3553 ( .C (clk), .D (signal_5095), .Q (signal_5096) ) ;
    buf_clk cell_3561 ( .C (clk), .D (signal_5103), .Q (signal_5104) ) ;
    buf_clk cell_3569 ( .C (clk), .D (signal_5111), .Q (signal_5112) ) ;
    buf_clk cell_3577 ( .C (clk), .D (signal_5119), .Q (signal_5120) ) ;
    buf_clk cell_3585 ( .C (clk), .D (signal_5127), .Q (signal_5128) ) ;
    buf_clk cell_3593 ( .C (clk), .D (signal_5135), .Q (signal_5136) ) ;
    buf_clk cell_3601 ( .C (clk), .D (signal_5143), .Q (signal_5144) ) ;
    buf_clk cell_3609 ( .C (clk), .D (signal_5151), .Q (signal_5152) ) ;
    buf_clk cell_3617 ( .C (clk), .D (signal_5159), .Q (signal_5160) ) ;
    buf_clk cell_3625 ( .C (clk), .D (signal_5167), .Q (signal_5168) ) ;
    buf_clk cell_3633 ( .C (clk), .D (signal_5175), .Q (signal_5176) ) ;
    buf_clk cell_3641 ( .C (clk), .D (signal_5183), .Q (signal_5184) ) ;
    buf_clk cell_3649 ( .C (clk), .D (signal_5191), .Q (signal_5192) ) ;
    buf_clk cell_3657 ( .C (clk), .D (signal_5199), .Q (signal_5200) ) ;
    buf_clk cell_3665 ( .C (clk), .D (signal_5207), .Q (signal_5208) ) ;
    buf_clk cell_3673 ( .C (clk), .D (signal_5215), .Q (signal_5216) ) ;
    buf_clk cell_3681 ( .C (clk), .D (signal_5223), .Q (signal_5224) ) ;
    buf_clk cell_3689 ( .C (clk), .D (signal_5231), .Q (signal_5232) ) ;
    buf_clk cell_3697 ( .C (clk), .D (signal_5239), .Q (signal_5240) ) ;
    buf_clk cell_3705 ( .C (clk), .D (signal_5247), .Q (signal_5248) ) ;
    buf_clk cell_3713 ( .C (clk), .D (signal_5255), .Q (signal_5256) ) ;
    buf_clk cell_3721 ( .C (clk), .D (signal_5263), .Q (signal_5264) ) ;
    buf_clk cell_3729 ( .C (clk), .D (signal_5271), .Q (signal_5272) ) ;
    buf_clk cell_3737 ( .C (clk), .D (signal_5279), .Q (signal_5280) ) ;
    buf_clk cell_3745 ( .C (clk), .D (signal_5287), .Q (signal_5288) ) ;
    buf_clk cell_3753 ( .C (clk), .D (signal_5295), .Q (signal_5296) ) ;
    buf_clk cell_3761 ( .C (clk), .D (signal_5303), .Q (signal_5304) ) ;
    buf_clk cell_3769 ( .C (clk), .D (signal_5311), .Q (signal_5312) ) ;
    buf_clk cell_3777 ( .C (clk), .D (signal_5319), .Q (signal_5320) ) ;
    buf_clk cell_3785 ( .C (clk), .D (signal_5327), .Q (signal_5328) ) ;
    buf_clk cell_3793 ( .C (clk), .D (signal_5335), .Q (signal_5336) ) ;
    buf_clk cell_3801 ( .C (clk), .D (signal_5343), .Q (signal_5344) ) ;
    buf_clk cell_3809 ( .C (clk), .D (signal_5351), .Q (signal_5352) ) ;
    buf_clk cell_3817 ( .C (clk), .D (signal_5359), .Q (signal_5360) ) ;
    buf_clk cell_3825 ( .C (clk), .D (signal_5367), .Q (signal_5368) ) ;
    buf_clk cell_3833 ( .C (clk), .D (signal_5375), .Q (signal_5376) ) ;
    buf_clk cell_3841 ( .C (clk), .D (signal_5383), .Q (signal_5384) ) ;
    buf_clk cell_3849 ( .C (clk), .D (signal_5391), .Q (signal_5392) ) ;
    buf_clk cell_3857 ( .C (clk), .D (signal_5399), .Q (signal_5400) ) ;
    buf_clk cell_3865 ( .C (clk), .D (signal_5407), .Q (signal_5408) ) ;
    buf_clk cell_3873 ( .C (clk), .D (signal_5415), .Q (signal_5416) ) ;
    buf_clk cell_3881 ( .C (clk), .D (signal_5423), .Q (signal_5424) ) ;
    buf_clk cell_3889 ( .C (clk), .D (signal_5431), .Q (signal_5432) ) ;
    buf_clk cell_3897 ( .C (clk), .D (signal_5439), .Q (signal_5440) ) ;
    buf_clk cell_3905 ( .C (clk), .D (signal_5447), .Q (signal_5448) ) ;
    buf_clk cell_3913 ( .C (clk), .D (signal_5455), .Q (signal_5456) ) ;
    buf_clk cell_3921 ( .C (clk), .D (signal_5463), .Q (signal_5464) ) ;
    buf_clk cell_3929 ( .C (clk), .D (signal_5471), .Q (signal_5472) ) ;
    buf_clk cell_3937 ( .C (clk), .D (signal_5479), .Q (signal_5480) ) ;
    buf_clk cell_3945 ( .C (clk), .D (signal_5487), .Q (signal_5488) ) ;
    buf_clk cell_3953 ( .C (clk), .D (signal_5495), .Q (signal_5496) ) ;
    buf_clk cell_3961 ( .C (clk), .D (signal_5503), .Q (signal_5504) ) ;
    buf_clk cell_3969 ( .C (clk), .D (signal_5511), .Q (signal_5512) ) ;
    buf_clk cell_3977 ( .C (clk), .D (signal_5519), .Q (signal_5520) ) ;
    buf_clk cell_3985 ( .C (clk), .D (signal_5527), .Q (signal_5528) ) ;
    buf_clk cell_3993 ( .C (clk), .D (signal_5535), .Q (signal_5536) ) ;
    buf_clk cell_4001 ( .C (clk), .D (signal_5543), .Q (signal_5544) ) ;
    buf_clk cell_4009 ( .C (clk), .D (signal_5551), .Q (signal_5552) ) ;
    buf_clk cell_4017 ( .C (clk), .D (signal_5559), .Q (signal_5560) ) ;
    buf_clk cell_4025 ( .C (clk), .D (signal_5567), .Q (signal_5568) ) ;
    buf_clk cell_4033 ( .C (clk), .D (signal_5575), .Q (signal_5576) ) ;
    buf_clk cell_4041 ( .C (clk), .D (signal_5583), .Q (signal_5584) ) ;
    buf_clk cell_4049 ( .C (clk), .D (signal_5591), .Q (signal_5592) ) ;
    buf_clk cell_4057 ( .C (clk), .D (signal_5599), .Q (signal_5600) ) ;
    buf_clk cell_4065 ( .C (clk), .D (signal_5607), .Q (signal_5608) ) ;
    buf_clk cell_4073 ( .C (clk), .D (signal_5615), .Q (signal_5616) ) ;
    buf_clk cell_4081 ( .C (clk), .D (signal_5623), .Q (signal_5624) ) ;
    buf_clk cell_4089 ( .C (clk), .D (signal_5631), .Q (signal_5632) ) ;
    buf_clk cell_4097 ( .C (clk), .D (signal_5639), .Q (signal_5640) ) ;
    buf_clk cell_4105 ( .C (clk), .D (signal_5647), .Q (signal_5648) ) ;
    buf_clk cell_4113 ( .C (clk), .D (signal_5655), .Q (signal_5656) ) ;
    buf_clk cell_4121 ( .C (clk), .D (signal_5663), .Q (signal_5664) ) ;
    buf_clk cell_4129 ( .C (clk), .D (signal_5671), .Q (signal_5672) ) ;
    buf_clk cell_4131 ( .C (clk), .D (signal_5673), .Q (signal_5674) ) ;
    buf_clk cell_4139 ( .C (clk), .D (signal_5681), .Q (signal_5682) ) ;
    buf_clk cell_4147 ( .C (clk), .D (signal_5689), .Q (signal_5690) ) ;
    buf_clk cell_4155 ( .C (clk), .D (signal_5697), .Q (signal_5698) ) ;
    buf_clk cell_4163 ( .C (clk), .D (signal_5705), .Q (signal_5706) ) ;
    buf_clk cell_4171 ( .C (clk), .D (signal_5713), .Q (signal_5714) ) ;
    buf_clk cell_4179 ( .C (clk), .D (signal_5721), .Q (signal_5722) ) ;
    buf_clk cell_4187 ( .C (clk), .D (signal_5729), .Q (signal_5730) ) ;
    buf_clk cell_4195 ( .C (clk), .D (signal_5737), .Q (signal_5738) ) ;
    buf_clk cell_4203 ( .C (clk), .D (signal_5745), .Q (signal_5746) ) ;
    buf_clk cell_4211 ( .C (clk), .D (signal_5753), .Q (signal_5754) ) ;
    buf_clk cell_4219 ( .C (clk), .D (signal_5761), .Q (signal_5762) ) ;
    buf_clk cell_4227 ( .C (clk), .D (signal_5769), .Q (signal_5770) ) ;
    buf_clk cell_4235 ( .C (clk), .D (signal_5777), .Q (signal_5778) ) ;
    buf_clk cell_4243 ( .C (clk), .D (signal_5785), .Q (signal_5786) ) ;
    buf_clk cell_4251 ( .C (clk), .D (signal_5793), .Q (signal_5794) ) ;
    buf_clk cell_4259 ( .C (clk), .D (signal_5801), .Q (signal_5802) ) ;
    buf_clk cell_4267 ( .C (clk), .D (signal_5809), .Q (signal_5810) ) ;
    buf_clk cell_4275 ( .C (clk), .D (signal_5817), .Q (signal_5818) ) ;
    buf_clk cell_4283 ( .C (clk), .D (signal_5825), .Q (signal_5826) ) ;
    buf_clk cell_4291 ( .C (clk), .D (signal_5833), .Q (signal_5834) ) ;
    buf_clk cell_4299 ( .C (clk), .D (signal_5841), .Q (signal_5842) ) ;
    buf_clk cell_4307 ( .C (clk), .D (signal_5849), .Q (signal_5850) ) ;
    buf_clk cell_4315 ( .C (clk), .D (signal_5857), .Q (signal_5858) ) ;
    buf_clk cell_4323 ( .C (clk), .D (signal_5865), .Q (signal_5866) ) ;
    buf_clk cell_4331 ( .C (clk), .D (signal_5873), .Q (signal_5874) ) ;
    buf_clk cell_4339 ( .C (clk), .D (signal_5881), .Q (signal_5882) ) ;
    buf_clk cell_4347 ( .C (clk), .D (signal_5889), .Q (signal_5890) ) ;
    buf_clk cell_4355 ( .C (clk), .D (signal_5897), .Q (signal_5898) ) ;
    buf_clk cell_4363 ( .C (clk), .D (signal_5905), .Q (signal_5906) ) ;
    buf_clk cell_4371 ( .C (clk), .D (signal_5913), .Q (signal_5914) ) ;
    buf_clk cell_4379 ( .C (clk), .D (signal_5921), .Q (signal_5922) ) ;
    buf_clk cell_4387 ( .C (clk), .D (signal_5929), .Q (signal_5930) ) ;
    buf_clk cell_4395 ( .C (clk), .D (signal_5937), .Q (signal_5938) ) ;
    buf_clk cell_4403 ( .C (clk), .D (signal_5945), .Q (signal_5946) ) ;
    buf_clk cell_4411 ( .C (clk), .D (signal_5953), .Q (signal_5954) ) ;
    buf_clk cell_4419 ( .C (clk), .D (signal_5961), .Q (signal_5962) ) ;
    buf_clk cell_4427 ( .C (clk), .D (signal_5969), .Q (signal_5970) ) ;
    buf_clk cell_4435 ( .C (clk), .D (signal_5977), .Q (signal_5978) ) ;
    buf_clk cell_4443 ( .C (clk), .D (signal_5985), .Q (signal_5986) ) ;
    buf_clk cell_4451 ( .C (clk), .D (signal_5993), .Q (signal_5994) ) ;
    buf_clk cell_4459 ( .C (clk), .D (signal_6001), .Q (signal_6002) ) ;
    buf_clk cell_4467 ( .C (clk), .D (signal_6009), .Q (signal_6010) ) ;
    buf_clk cell_4475 ( .C (clk), .D (signal_6017), .Q (signal_6018) ) ;
    buf_clk cell_4483 ( .C (clk), .D (signal_6025), .Q (signal_6026) ) ;
    buf_clk cell_4491 ( .C (clk), .D (signal_6033), .Q (signal_6034) ) ;
    buf_clk cell_4499 ( .C (clk), .D (signal_6041), .Q (signal_6042) ) ;
    buf_clk cell_4507 ( .C (clk), .D (signal_6049), .Q (signal_6050) ) ;
    buf_clk cell_4515 ( .C (clk), .D (signal_6057), .Q (signal_6058) ) ;
    buf_clk cell_4523 ( .C (clk), .D (signal_6065), .Q (signal_6066) ) ;
    buf_clk cell_4531 ( .C (clk), .D (signal_6073), .Q (signal_6074) ) ;
    buf_clk cell_4539 ( .C (clk), .D (signal_6081), .Q (signal_6082) ) ;
    buf_clk cell_4547 ( .C (clk), .D (signal_6089), .Q (signal_6090) ) ;
    buf_clk cell_4555 ( .C (clk), .D (signal_6097), .Q (signal_6098) ) ;
    buf_clk cell_4563 ( .C (clk), .D (signal_6105), .Q (signal_6106) ) ;
    buf_clk cell_4571 ( .C (clk), .D (signal_6113), .Q (signal_6114) ) ;
    buf_clk cell_4579 ( .C (clk), .D (signal_6121), .Q (signal_6122) ) ;
    buf_clk cell_4587 ( .C (clk), .D (signal_6129), .Q (signal_6130) ) ;
    buf_clk cell_4595 ( .C (clk), .D (signal_6137), .Q (signal_6138) ) ;
    buf_clk cell_4603 ( .C (clk), .D (signal_6145), .Q (signal_6146) ) ;
    buf_clk cell_4611 ( .C (clk), .D (signal_6153), .Q (signal_6154) ) ;
    buf_clk cell_4619 ( .C (clk), .D (signal_6161), .Q (signal_6162) ) ;
    buf_clk cell_4627 ( .C (clk), .D (signal_6169), .Q (signal_6170) ) ;
    buf_clk cell_4635 ( .C (clk), .D (signal_6177), .Q (signal_6178) ) ;
    buf_clk cell_4643 ( .C (clk), .D (signal_6185), .Q (signal_6186) ) ;
    buf_clk cell_4645 ( .C (clk), .D (signal_6187), .Q (signal_6188) ) ;
    buf_clk cell_4845 ( .C (clk), .D (signal_6387), .Q (signal_6388) ) ;
    buf_clk cell_4853 ( .C (clk), .D (signal_6395), .Q (signal_6396) ) ;
    buf_clk cell_4861 ( .C (clk), .D (signal_6403), .Q (signal_6404) ) ;
    buf_clk cell_4869 ( .C (clk), .D (signal_6411), .Q (signal_6412) ) ;
    buf_clk cell_4871 ( .C (clk), .D (signal_6413), .Q (signal_6414) ) ;
    buf_clk cell_4873 ( .C (clk), .D (signal_6415), .Q (signal_6416) ) ;
    buf_clk cell_4875 ( .C (clk), .D (signal_6417), .Q (signal_6418) ) ;
    buf_clk cell_4877 ( .C (clk), .D (signal_6419), .Q (signal_6420) ) ;
    buf_clk cell_4879 ( .C (clk), .D (signal_6421), .Q (signal_6422) ) ;
    buf_clk cell_4881 ( .C (clk), .D (signal_6423), .Q (signal_6424) ) ;
    buf_clk cell_4883 ( .C (clk), .D (signal_6425), .Q (signal_6426) ) ;
    buf_clk cell_4885 ( .C (clk), .D (signal_6427), .Q (signal_6428) ) ;
    buf_clk cell_4887 ( .C (clk), .D (signal_6429), .Q (signal_6430) ) ;
    buf_clk cell_4889 ( .C (clk), .D (signal_6431), .Q (signal_6432) ) ;
    buf_clk cell_4891 ( .C (clk), .D (signal_6433), .Q (signal_6434) ) ;
    buf_clk cell_4893 ( .C (clk), .D (signal_6435), .Q (signal_6436) ) ;
    buf_clk cell_4895 ( .C (clk), .D (signal_6437), .Q (signal_6438) ) ;
    buf_clk cell_4897 ( .C (clk), .D (signal_6439), .Q (signal_6440) ) ;
    buf_clk cell_4899 ( .C (clk), .D (signal_6441), .Q (signal_6442) ) ;
    buf_clk cell_4901 ( .C (clk), .D (signal_6443), .Q (signal_6444) ) ;
    buf_clk cell_4903 ( .C (clk), .D (signal_6445), .Q (signal_6446) ) ;
    buf_clk cell_4905 ( .C (clk), .D (signal_6447), .Q (signal_6448) ) ;
    buf_clk cell_4907 ( .C (clk), .D (signal_6449), .Q (signal_6450) ) ;
    buf_clk cell_4909 ( .C (clk), .D (signal_6451), .Q (signal_6452) ) ;
    buf_clk cell_4911 ( .C (clk), .D (signal_6453), .Q (signal_6454) ) ;
    buf_clk cell_4913 ( .C (clk), .D (signal_6455), .Q (signal_6456) ) ;
    buf_clk cell_4915 ( .C (clk), .D (signal_6457), .Q (signal_6458) ) ;
    buf_clk cell_4917 ( .C (clk), .D (signal_6459), .Q (signal_6460) ) ;
    buf_clk cell_4919 ( .C (clk), .D (signal_6461), .Q (signal_6462) ) ;
    buf_clk cell_4921 ( .C (clk), .D (signal_6463), .Q (signal_6464) ) ;
    buf_clk cell_4923 ( .C (clk), .D (signal_6465), .Q (signal_6466) ) ;
    buf_clk cell_4925 ( .C (clk), .D (signal_6467), .Q (signal_6468) ) ;
    buf_clk cell_4927 ( .C (clk), .D (signal_6469), .Q (signal_6470) ) ;
    buf_clk cell_4929 ( .C (clk), .D (signal_6471), .Q (signal_6472) ) ;
    buf_clk cell_4931 ( .C (clk), .D (signal_6473), .Q (signal_6474) ) ;
    buf_clk cell_4933 ( .C (clk), .D (signal_6475), .Q (signal_6476) ) ;
    buf_clk cell_4935 ( .C (clk), .D (signal_6477), .Q (signal_6478) ) ;
    buf_clk cell_4937 ( .C (clk), .D (signal_6479), .Q (signal_6480) ) ;
    buf_clk cell_4939 ( .C (clk), .D (signal_6481), .Q (signal_6482) ) ;
    buf_clk cell_4941 ( .C (clk), .D (signal_6483), .Q (signal_6484) ) ;
    buf_clk cell_4943 ( .C (clk), .D (signal_6485), .Q (signal_6486) ) ;
    buf_clk cell_4945 ( .C (clk), .D (signal_6487), .Q (signal_6488) ) ;
    buf_clk cell_4947 ( .C (clk), .D (signal_6489), .Q (signal_6490) ) ;
    buf_clk cell_4949 ( .C (clk), .D (signal_6491), .Q (signal_6492) ) ;
    buf_clk cell_4951 ( .C (clk), .D (signal_6493), .Q (signal_6494) ) ;
    buf_clk cell_4953 ( .C (clk), .D (signal_6495), .Q (signal_6496) ) ;
    buf_clk cell_4955 ( .C (clk), .D (signal_6497), .Q (signal_6498) ) ;
    buf_clk cell_4957 ( .C (clk), .D (signal_6499), .Q (signal_6500) ) ;
    buf_clk cell_4959 ( .C (clk), .D (signal_6501), .Q (signal_6502) ) ;
    buf_clk cell_4961 ( .C (clk), .D (signal_6503), .Q (signal_6504) ) ;
    buf_clk cell_4963 ( .C (clk), .D (signal_6505), .Q (signal_6506) ) ;
    buf_clk cell_4965 ( .C (clk), .D (signal_6507), .Q (signal_6508) ) ;
    buf_clk cell_4967 ( .C (clk), .D (signal_6509), .Q (signal_6510) ) ;
    buf_clk cell_4969 ( .C (clk), .D (signal_6511), .Q (signal_6512) ) ;
    buf_clk cell_4971 ( .C (clk), .D (signal_6513), .Q (signal_6514) ) ;
    buf_clk cell_4973 ( .C (clk), .D (signal_6515), .Q (signal_6516) ) ;
    buf_clk cell_4975 ( .C (clk), .D (signal_6517), .Q (signal_6518) ) ;
    buf_clk cell_4977 ( .C (clk), .D (signal_6519), .Q (signal_6520) ) ;
    buf_clk cell_4979 ( .C (clk), .D (signal_6521), .Q (signal_6522) ) ;
    buf_clk cell_4981 ( .C (clk), .D (signal_6523), .Q (signal_6524) ) ;
    buf_clk cell_4983 ( .C (clk), .D (signal_6525), .Q (signal_6526) ) ;
    buf_clk cell_4985 ( .C (clk), .D (signal_6527), .Q (signal_6528) ) ;
    buf_clk cell_4987 ( .C (clk), .D (signal_6529), .Q (signal_6530) ) ;
    buf_clk cell_4989 ( .C (clk), .D (signal_6531), .Q (signal_6532) ) ;
    buf_clk cell_4991 ( .C (clk), .D (signal_6533), .Q (signal_6534) ) ;
    buf_clk cell_4993 ( .C (clk), .D (signal_6535), .Q (signal_6536) ) ;
    buf_clk cell_4995 ( .C (clk), .D (signal_6537), .Q (signal_6538) ) ;
    buf_clk cell_4997 ( .C (clk), .D (signal_6539), .Q (signal_6540) ) ;

    /* register cells */
    DFF_X1 cell_82 ( .CK (clk), .D (signal_6388), .Q (signal_927), .QN () ) ;
    DFF_X1 cell_84 ( .CK (clk), .D (signal_6396), .Q (signal_926), .QN () ) ;
    DFF_X1 cell_86 ( .CK (clk), .D (signal_6404), .Q (signal_925), .QN () ) ;
    DFF_X1 cell_88 ( .CK (clk), .D (signal_6412), .Q (signal_924), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_537 ( .clk (clk), .D ({signal_2777, signal_460}), .Q ({signal_2052, signal_1375}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_540 ( .clk (clk), .D ({signal_6416, signal_6414}), .Q ({signal_2224, signal_1374}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_543 ( .clk (clk), .D ({signal_2691, signal_464}), .Q ({signal_1841, signal_1373}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_546 ( .clk (clk), .D ({signal_6420, signal_6418}), .Q ({signal_1846, signal_1372}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_549 ( .clk (clk), .D ({signal_2778, signal_468}), .Q ({signal_2072, signal_1371}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_552 ( .clk (clk), .D ({signal_6424, signal_6422}), .Q ({signal_2233, signal_1370}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_555 ( .clk (clk), .D ({signal_2692, signal_472}), .Q ({signal_1836, signal_1369}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_558 ( .clk (clk), .D ({signal_6428, signal_6426}), .Q ({signal_1828, signal_1368}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_561 ( .clk (clk), .D ({signal_2779, signal_476}), .Q ({signal_2135, signal_1367}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_564 ( .clk (clk), .D ({signal_6432, signal_6430}), .Q ({signal_2266, signal_1366}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_567 ( .clk (clk), .D ({signal_2693, signal_480}), .Q ({signal_1839, signal_1365}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_570 ( .clk (clk), .D ({signal_6436, signal_6434}), .Q ({signal_1888, signal_1364}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_573 ( .clk (clk), .D ({signal_2780, signal_484}), .Q ({signal_2128, signal_1363}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_576 ( .clk (clk), .D ({signal_6440, signal_6438}), .Q ({signal_2261, signal_1362}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_579 ( .clk (clk), .D ({signal_2694, signal_488}), .Q ({signal_1883, signal_1361}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_582 ( .clk (clk), .D ({signal_6444, signal_6442}), .Q ({signal_1885, signal_1360}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_585 ( .clk (clk), .D ({signal_2791, signal_492}), .Q ({signal_2121, signal_1359}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_588 ( .clk (clk), .D ({signal_6448, signal_6446}), .Q ({signal_2256, signal_1358}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_591 ( .clk (clk), .D ({signal_2695, signal_496}), .Q ({signal_1878, signal_1357}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_594 ( .clk (clk), .D ({signal_6452, signal_6450}), .Q ({signal_1880, signal_1356}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_597 ( .clk (clk), .D ({signal_2792, signal_500}), .Q ({signal_2113, signal_1355}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_600 ( .clk (clk), .D ({signal_6456, signal_6454}), .Q ({signal_2250, signal_1354}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_603 ( .clk (clk), .D ({signal_2696, signal_504}), .Q ({signal_1873, signal_1353}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_606 ( .clk (clk), .D ({signal_6460, signal_6458}), .Q ({signal_1875, signal_1352}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_609 ( .clk (clk), .D ({signal_2781, signal_508}), .Q ({signal_2106, signal_1351}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_612 ( .clk (clk), .D ({signal_6464, signal_6462}), .Q ({signal_2245, signal_1350}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_615 ( .clk (clk), .D ({signal_2697, signal_512}), .Q ({signal_1868, signal_1349}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_618 ( .clk (clk), .D ({signal_6468, signal_6466}), .Q ({signal_1870, signal_1348}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_621 ( .clk (clk), .D ({signal_2782, signal_516}), .Q ({signal_2067, signal_1347}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_624 ( .clk (clk), .D ({signal_6472, signal_6470}), .Q ({signal_2239, signal_1346}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_627 ( .clk (clk), .D ({signal_2698, signal_520}), .Q ({signal_2098, signal_1345}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_630 ( .clk (clk), .D ({signal_6476, signal_6474}), .Q ({signal_1834, signal_1344}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_633 ( .clk (clk), .D ({signal_2783, signal_524}), .Q ({signal_2070, signal_1343}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_636 ( .clk (clk), .D ({signal_6480, signal_6478}), .Q ({signal_2219, signal_1342}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_639 ( .clk (clk), .D ({signal_2699, signal_528}), .Q ({signal_2018, signal_1341}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_642 ( .clk (clk), .D ({signal_6484, signal_6482}), .Q ({signal_1843, signal_1340}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_645 ( .clk (clk), .D ({signal_2784, signal_532}), .Q ({signal_2056, signal_1339}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_648 ( .clk (clk), .D ({signal_6488, signal_6486}), .Q ({signal_2211, signal_1338}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_651 ( .clk (clk), .D ({signal_2700, signal_536}), .Q ({signal_2035, signal_1337}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_654 ( .clk (clk), .D ({signal_6492, signal_6490}), .Q ({signal_1860, signal_1336}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_657 ( .clk (clk), .D ({signal_2785, signal_540}), .Q ({signal_2064, signal_1335}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_660 ( .clk (clk), .D ({signal_6496, signal_6494}), .Q ({signal_2191, signal_1334}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_663 ( .clk (clk), .D ({signal_2701, signal_544}), .Q ({signal_2033, signal_1333}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_666 ( .clk (clk), .D ({signal_6500, signal_6498}), .Q ({signal_1830, signal_1332}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_669 ( .clk (clk), .D ({signal_2786, signal_548}), .Q ({signal_2043, signal_1331}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_672 ( .clk (clk), .D ({signal_6504, signal_6502}), .Q ({signal_2202, signal_1330}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_675 ( .clk (clk), .D ({signal_2702, signal_552}), .Q ({signal_2059, signal_1329}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_678 ( .clk (clk), .D ({signal_6508, signal_6506}), .Q ({signal_1854, signal_1328}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_681 ( .clk (clk), .D ({signal_2787, signal_556}), .Q ({signal_2094, signal_1327}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_684 ( .clk (clk), .D ({signal_6512, signal_6510}), .Q ({signal_2205, signal_1326}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_687 ( .clk (clk), .D ({signal_2703, signal_560}), .Q ({signal_2022, signal_1325}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_690 ( .clk (clk), .D ({signal_6516, signal_6514}), .Q ({signal_1856, signal_1324}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_693 ( .clk (clk), .D ({signal_2793, signal_564}), .Q ({signal_2024, signal_1323}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_696 ( .clk (clk), .D ({signal_6520, signal_6518}), .Q ({signal_2230, signal_1322}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_699 ( .clk (clk), .D ({signal_2704, signal_568}), .Q ({signal_2030, signal_1321}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_702 ( .clk (clk), .D ({signal_6524, signal_6522}), .Q ({signal_1850, signal_1320}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_705 ( .clk (clk), .D ({signal_2796, signal_572}), .Q ({signal_2045, signal_1319}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_708 ( .clk (clk), .D ({signal_6528, signal_6526}), .Q ({signal_2226, signal_1318}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_711 ( .clk (clk), .D ({signal_2705, signal_576}), .Q ({signal_2038, signal_1317}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_714 ( .clk (clk), .D ({signal_6532, signal_6530}), .Q ({signal_1832, signal_1316}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_717 ( .clk (clk), .D ({signal_2797, signal_580}), .Q ({signal_2075, signal_1315}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_720 ( .clk (clk), .D ({signal_6536, signal_6534}), .Q ({signal_2217, signal_1314}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_723 ( .clk (clk), .D ({signal_2706, signal_584}), .Q ({signal_2026, signal_1313}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_726 ( .clk (clk), .D ({signal_6540, signal_6538}), .Q ({signal_1862, signal_1312}) ) ;
endmodule
