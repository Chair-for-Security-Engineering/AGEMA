/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_Pipeline_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input [339:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_161 ;
    wire new_AGEMA_signal_162 ;
    wire new_AGEMA_signal_167 ;
    wire new_AGEMA_signal_168 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_181 ;
    wire new_AGEMA_signal_182 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;
    wire new_AGEMA_signal_593 ;
    wire new_AGEMA_signal_594 ;
    wire new_AGEMA_signal_595 ;
    wire new_AGEMA_signal_596 ;
    wire new_AGEMA_signal_597 ;
    wire new_AGEMA_signal_598 ;
    wire new_AGEMA_signal_599 ;
    wire new_AGEMA_signal_600 ;
    wire new_AGEMA_signal_601 ;
    wire new_AGEMA_signal_602 ;
    wire new_AGEMA_signal_603 ;
    wire new_AGEMA_signal_604 ;
    wire new_AGEMA_signal_605 ;
    wire new_AGEMA_signal_606 ;
    wire new_AGEMA_signal_607 ;
    wire new_AGEMA_signal_608 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;
    wire new_AGEMA_signal_656 ;
    wire new_AGEMA_signal_657 ;
    wire new_AGEMA_signal_658 ;
    wire new_AGEMA_signal_659 ;
    wire new_AGEMA_signal_660 ;
    wire new_AGEMA_signal_661 ;
    wire new_AGEMA_signal_662 ;
    wire new_AGEMA_signal_663 ;
    wire new_AGEMA_signal_664 ;
    wire new_AGEMA_signal_665 ;
    wire new_AGEMA_signal_666 ;
    wire new_AGEMA_signal_667 ;
    wire new_AGEMA_signal_668 ;
    wire new_AGEMA_signal_669 ;
    wire new_AGEMA_signal_670 ;
    wire new_AGEMA_signal_671 ;
    wire new_AGEMA_signal_672 ;
    wire new_AGEMA_signal_673 ;
    wire new_AGEMA_signal_674 ;
    wire new_AGEMA_signal_675 ;
    wire new_AGEMA_signal_676 ;
    wire new_AGEMA_signal_677 ;
    wire new_AGEMA_signal_678 ;
    wire new_AGEMA_signal_679 ;
    wire new_AGEMA_signal_680 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T1_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T2_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T3_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T4_U1 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T5_U1 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T6_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .c ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T7_U1 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T8_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .c ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, T8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T9_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .c ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T10_U1 ( .a ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .b ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .c ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T11_U1 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T12_U1 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T13_U1 ( .a ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .b ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}), .c ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, new_AGEMA_signal_231, T13}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T14_U1 ( .a ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .b ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}), .c ({new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, new_AGEMA_signal_263, T14}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T15_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .b ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}), .c ({new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T15}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T16_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}), .c ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T17_U1 ( .a ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}), .b ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .c ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T18_U1 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, new_AGEMA_signal_215, T18}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T19_U1 ( .a ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, new_AGEMA_signal_215, T18}), .c ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T20_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}), .c ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T21_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, T21}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T22_U1 ( .a ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, T21}), .c ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T23_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .b ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}), .c ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, new_AGEMA_signal_275, T23}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T24_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .b ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}), .c ({new_AGEMA_signal_310, new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, T24}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T25_U1 ( .a ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}), .b ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}), .c ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, new_AGEMA_signal_311, T25}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T26_U1 ( .a ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .b ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .c ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, new_AGEMA_signal_279, T26}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_T27_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}), .c ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, new_AGEMA_signal_251, T27}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_136 ( .C (clk), .D (T14), .Q (new_AGEMA_signal_1067) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C (clk), .D (new_AGEMA_signal_263), .Q (new_AGEMA_signal_1069) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C (clk), .D (new_AGEMA_signal_264), .Q (new_AGEMA_signal_1071) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C (clk), .D (new_AGEMA_signal_265), .Q (new_AGEMA_signal_1073) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C (clk), .D (new_AGEMA_signal_266), .Q (new_AGEMA_signal_1075) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C (clk), .D (T26), .Q (new_AGEMA_signal_1077) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C (clk), .D (new_AGEMA_signal_279), .Q (new_AGEMA_signal_1079) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C (clk), .D (new_AGEMA_signal_280), .Q (new_AGEMA_signal_1081) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C (clk), .D (new_AGEMA_signal_281), .Q (new_AGEMA_signal_1083) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C (clk), .D (new_AGEMA_signal_282), .Q (new_AGEMA_signal_1085) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C (clk), .D (T24), .Q (new_AGEMA_signal_1087) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C (clk), .D (new_AGEMA_signal_307), .Q (new_AGEMA_signal_1089) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C (clk), .D (new_AGEMA_signal_308), .Q (new_AGEMA_signal_1091) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C (clk), .D (new_AGEMA_signal_309), .Q (new_AGEMA_signal_1093) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C (clk), .D (new_AGEMA_signal_310), .Q (new_AGEMA_signal_1095) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C (clk), .D (T25), .Q (new_AGEMA_signal_1097) ) ;
    buf_clk new_AGEMA_reg_buffer_168 ( .C (clk), .D (new_AGEMA_signal_311), .Q (new_AGEMA_signal_1099) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C (clk), .D (new_AGEMA_signal_312), .Q (new_AGEMA_signal_1101) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C (clk), .D (new_AGEMA_signal_313), .Q (new_AGEMA_signal_1103) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C (clk), .D (new_AGEMA_signal_314), .Q (new_AGEMA_signal_1105) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C (clk), .D (T6), .Q (new_AGEMA_signal_1187) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C (clk), .D (new_AGEMA_signal_223), .Q (new_AGEMA_signal_1193) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C (clk), .D (new_AGEMA_signal_224), .Q (new_AGEMA_signal_1199) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C (clk), .D (new_AGEMA_signal_225), .Q (new_AGEMA_signal_1205) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C (clk), .D (new_AGEMA_signal_226), .Q (new_AGEMA_signal_1211) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C (clk), .D (T8), .Q (new_AGEMA_signal_1217) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C (clk), .D (new_AGEMA_signal_255), .Q (new_AGEMA_signal_1223) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C (clk), .D (new_AGEMA_signal_256), .Q (new_AGEMA_signal_1229) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C (clk), .D (new_AGEMA_signal_257), .Q (new_AGEMA_signal_1235) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C (clk), .D (new_AGEMA_signal_258), .Q (new_AGEMA_signal_1241) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C (clk), .D (X_s0[0]), .Q (new_AGEMA_signal_1247) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C (clk), .D (X_s1[0]), .Q (new_AGEMA_signal_1253) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C (clk), .D (X_s2[0]), .Q (new_AGEMA_signal_1259) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C (clk), .D (X_s3[0]), .Q (new_AGEMA_signal_1265) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C (clk), .D (X_s4[0]), .Q (new_AGEMA_signal_1271) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C (clk), .D (T16), .Q (new_AGEMA_signal_1277) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C (clk), .D (new_AGEMA_signal_239), .Q (new_AGEMA_signal_1283) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C (clk), .D (new_AGEMA_signal_240), .Q (new_AGEMA_signal_1289) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C (clk), .D (new_AGEMA_signal_241), .Q (new_AGEMA_signal_1295) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C (clk), .D (new_AGEMA_signal_242), .Q (new_AGEMA_signal_1301) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C (clk), .D (T9), .Q (new_AGEMA_signal_1307) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C (clk), .D (new_AGEMA_signal_227), .Q (new_AGEMA_signal_1313) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C (clk), .D (new_AGEMA_signal_228), .Q (new_AGEMA_signal_1319) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C (clk), .D (new_AGEMA_signal_229), .Q (new_AGEMA_signal_1325) ) ;
    buf_clk new_AGEMA_reg_buffer_400 ( .C (clk), .D (new_AGEMA_signal_230), .Q (new_AGEMA_signal_1331) ) ;
    buf_clk new_AGEMA_reg_buffer_406 ( .C (clk), .D (T17), .Q (new_AGEMA_signal_1337) ) ;
    buf_clk new_AGEMA_reg_buffer_412 ( .C (clk), .D (new_AGEMA_signal_267), .Q (new_AGEMA_signal_1343) ) ;
    buf_clk new_AGEMA_reg_buffer_418 ( .C (clk), .D (new_AGEMA_signal_268), .Q (new_AGEMA_signal_1349) ) ;
    buf_clk new_AGEMA_reg_buffer_424 ( .C (clk), .D (new_AGEMA_signal_269), .Q (new_AGEMA_signal_1355) ) ;
    buf_clk new_AGEMA_reg_buffer_430 ( .C (clk), .D (new_AGEMA_signal_270), .Q (new_AGEMA_signal_1361) ) ;
    buf_clk new_AGEMA_reg_buffer_436 ( .C (clk), .D (T15), .Q (new_AGEMA_signal_1367) ) ;
    buf_clk new_AGEMA_reg_buffer_442 ( .C (clk), .D (new_AGEMA_signal_235), .Q (new_AGEMA_signal_1373) ) ;
    buf_clk new_AGEMA_reg_buffer_448 ( .C (clk), .D (new_AGEMA_signal_236), .Q (new_AGEMA_signal_1379) ) ;
    buf_clk new_AGEMA_reg_buffer_454 ( .C (clk), .D (new_AGEMA_signal_237), .Q (new_AGEMA_signal_1385) ) ;
    buf_clk new_AGEMA_reg_buffer_460 ( .C (clk), .D (new_AGEMA_signal_238), .Q (new_AGEMA_signal_1391) ) ;
    buf_clk new_AGEMA_reg_buffer_466 ( .C (clk), .D (T27), .Q (new_AGEMA_signal_1397) ) ;
    buf_clk new_AGEMA_reg_buffer_472 ( .C (clk), .D (new_AGEMA_signal_251), .Q (new_AGEMA_signal_1403) ) ;
    buf_clk new_AGEMA_reg_buffer_478 ( .C (clk), .D (new_AGEMA_signal_252), .Q (new_AGEMA_signal_1409) ) ;
    buf_clk new_AGEMA_reg_buffer_484 ( .C (clk), .D (new_AGEMA_signal_253), .Q (new_AGEMA_signal_1415) ) ;
    buf_clk new_AGEMA_reg_buffer_490 ( .C (clk), .D (new_AGEMA_signal_254), .Q (new_AGEMA_signal_1421) ) ;
    buf_clk new_AGEMA_reg_buffer_496 ( .C (clk), .D (T10), .Q (new_AGEMA_signal_1427) ) ;
    buf_clk new_AGEMA_reg_buffer_502 ( .C (clk), .D (new_AGEMA_signal_259), .Q (new_AGEMA_signal_1433) ) ;
    buf_clk new_AGEMA_reg_buffer_508 ( .C (clk), .D (new_AGEMA_signal_260), .Q (new_AGEMA_signal_1439) ) ;
    buf_clk new_AGEMA_reg_buffer_514 ( .C (clk), .D (new_AGEMA_signal_261), .Q (new_AGEMA_signal_1445) ) ;
    buf_clk new_AGEMA_reg_buffer_520 ( .C (clk), .D (new_AGEMA_signal_262), .Q (new_AGEMA_signal_1451) ) ;
    buf_clk new_AGEMA_reg_buffer_526 ( .C (clk), .D (T13), .Q (new_AGEMA_signal_1457) ) ;
    buf_clk new_AGEMA_reg_buffer_532 ( .C (clk), .D (new_AGEMA_signal_231), .Q (new_AGEMA_signal_1463) ) ;
    buf_clk new_AGEMA_reg_buffer_538 ( .C (clk), .D (new_AGEMA_signal_232), .Q (new_AGEMA_signal_1469) ) ;
    buf_clk new_AGEMA_reg_buffer_544 ( .C (clk), .D (new_AGEMA_signal_233), .Q (new_AGEMA_signal_1475) ) ;
    buf_clk new_AGEMA_reg_buffer_550 ( .C (clk), .D (new_AGEMA_signal_234), .Q (new_AGEMA_signal_1481) ) ;
    buf_clk new_AGEMA_reg_buffer_556 ( .C (clk), .D (T23), .Q (new_AGEMA_signal_1487) ) ;
    buf_clk new_AGEMA_reg_buffer_562 ( .C (clk), .D (new_AGEMA_signal_275), .Q (new_AGEMA_signal_1493) ) ;
    buf_clk new_AGEMA_reg_buffer_568 ( .C (clk), .D (new_AGEMA_signal_276), .Q (new_AGEMA_signal_1499) ) ;
    buf_clk new_AGEMA_reg_buffer_574 ( .C (clk), .D (new_AGEMA_signal_277), .Q (new_AGEMA_signal_1505) ) ;
    buf_clk new_AGEMA_reg_buffer_580 ( .C (clk), .D (new_AGEMA_signal_278), .Q (new_AGEMA_signal_1511) ) ;
    buf_clk new_AGEMA_reg_buffer_586 ( .C (clk), .D (T19), .Q (new_AGEMA_signal_1517) ) ;
    buf_clk new_AGEMA_reg_buffer_592 ( .C (clk), .D (new_AGEMA_signal_243), .Q (new_AGEMA_signal_1523) ) ;
    buf_clk new_AGEMA_reg_buffer_598 ( .C (clk), .D (new_AGEMA_signal_244), .Q (new_AGEMA_signal_1529) ) ;
    buf_clk new_AGEMA_reg_buffer_604 ( .C (clk), .D (new_AGEMA_signal_245), .Q (new_AGEMA_signal_1535) ) ;
    buf_clk new_AGEMA_reg_buffer_610 ( .C (clk), .D (new_AGEMA_signal_246), .Q (new_AGEMA_signal_1541) ) ;
    buf_clk new_AGEMA_reg_buffer_616 ( .C (clk), .D (T3), .Q (new_AGEMA_signal_1547) ) ;
    buf_clk new_AGEMA_reg_buffer_622 ( .C (clk), .D (new_AGEMA_signal_175), .Q (new_AGEMA_signal_1553) ) ;
    buf_clk new_AGEMA_reg_buffer_628 ( .C (clk), .D (new_AGEMA_signal_176), .Q (new_AGEMA_signal_1559) ) ;
    buf_clk new_AGEMA_reg_buffer_634 ( .C (clk), .D (new_AGEMA_signal_177), .Q (new_AGEMA_signal_1565) ) ;
    buf_clk new_AGEMA_reg_buffer_640 ( .C (clk), .D (new_AGEMA_signal_178), .Q (new_AGEMA_signal_1571) ) ;
    buf_clk new_AGEMA_reg_buffer_646 ( .C (clk), .D (T22), .Q (new_AGEMA_signal_1577) ) ;
    buf_clk new_AGEMA_reg_buffer_652 ( .C (clk), .D (new_AGEMA_signal_247), .Q (new_AGEMA_signal_1583) ) ;
    buf_clk new_AGEMA_reg_buffer_658 ( .C (clk), .D (new_AGEMA_signal_248), .Q (new_AGEMA_signal_1589) ) ;
    buf_clk new_AGEMA_reg_buffer_664 ( .C (clk), .D (new_AGEMA_signal_249), .Q (new_AGEMA_signal_1595) ) ;
    buf_clk new_AGEMA_reg_buffer_670 ( .C (clk), .D (new_AGEMA_signal_250), .Q (new_AGEMA_signal_1601) ) ;
    buf_clk new_AGEMA_reg_buffer_676 ( .C (clk), .D (T20), .Q (new_AGEMA_signal_1607) ) ;
    buf_clk new_AGEMA_reg_buffer_682 ( .C (clk), .D (new_AGEMA_signal_271), .Q (new_AGEMA_signal_1613) ) ;
    buf_clk new_AGEMA_reg_buffer_688 ( .C (clk), .D (new_AGEMA_signal_272), .Q (new_AGEMA_signal_1619) ) ;
    buf_clk new_AGEMA_reg_buffer_694 ( .C (clk), .D (new_AGEMA_signal_273), .Q (new_AGEMA_signal_1625) ) ;
    buf_clk new_AGEMA_reg_buffer_700 ( .C (clk), .D (new_AGEMA_signal_274), .Q (new_AGEMA_signal_1631) ) ;
    buf_clk new_AGEMA_reg_buffer_706 ( .C (clk), .D (T1), .Q (new_AGEMA_signal_1637) ) ;
    buf_clk new_AGEMA_reg_buffer_712 ( .C (clk), .D (new_AGEMA_signal_159), .Q (new_AGEMA_signal_1643) ) ;
    buf_clk new_AGEMA_reg_buffer_718 ( .C (clk), .D (new_AGEMA_signal_160), .Q (new_AGEMA_signal_1649) ) ;
    buf_clk new_AGEMA_reg_buffer_724 ( .C (clk), .D (new_AGEMA_signal_161), .Q (new_AGEMA_signal_1655) ) ;
    buf_clk new_AGEMA_reg_buffer_730 ( .C (clk), .D (new_AGEMA_signal_162), .Q (new_AGEMA_signal_1661) ) ;
    buf_clk new_AGEMA_reg_buffer_736 ( .C (clk), .D (T4), .Q (new_AGEMA_signal_1667) ) ;
    buf_clk new_AGEMA_reg_buffer_742 ( .C (clk), .D (new_AGEMA_signal_179), .Q (new_AGEMA_signal_1673) ) ;
    buf_clk new_AGEMA_reg_buffer_748 ( .C (clk), .D (new_AGEMA_signal_180), .Q (new_AGEMA_signal_1679) ) ;
    buf_clk new_AGEMA_reg_buffer_754 ( .C (clk), .D (new_AGEMA_signal_181), .Q (new_AGEMA_signal_1685) ) ;
    buf_clk new_AGEMA_reg_buffer_760 ( .C (clk), .D (new_AGEMA_signal_182), .Q (new_AGEMA_signal_1691) ) ;
    buf_clk new_AGEMA_reg_buffer_766 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_1697) ) ;
    buf_clk new_AGEMA_reg_buffer_772 ( .C (clk), .D (new_AGEMA_signal_167), .Q (new_AGEMA_signal_1703) ) ;
    buf_clk new_AGEMA_reg_buffer_778 ( .C (clk), .D (new_AGEMA_signal_168), .Q (new_AGEMA_signal_1709) ) ;
    buf_clk new_AGEMA_reg_buffer_784 ( .C (clk), .D (new_AGEMA_signal_169), .Q (new_AGEMA_signal_1715) ) ;
    buf_clk new_AGEMA_reg_buffer_790 ( .C (clk), .D (new_AGEMA_signal_170), .Q (new_AGEMA_signal_1721) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M1_U1 ( .a ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, new_AGEMA_signal_231, T13}), .b ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M2_U1 ( .a ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, new_AGEMA_signal_275, T23}), .b ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, T8}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, M2}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M3_U1 ( .a ({new_AGEMA_signal_1076, new_AGEMA_signal_1074, new_AGEMA_signal_1072, new_AGEMA_signal_1070, new_AGEMA_signal_1068}), .b ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}), .c ({new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M3}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M4_U1 ( .a ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, new_AGEMA_signal_287, M4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M5_U1 ( .a ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, new_AGEMA_signal_287, M4}), .b ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}), .c ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, new_AGEMA_signal_323, M5}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M6_U1 ( .a ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .b ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M7_U1 ( .a ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}), .b ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}), .clk (clk), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M7}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M8_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1084, new_AGEMA_signal_1082, new_AGEMA_signal_1080, new_AGEMA_signal_1078}), .b ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}), .c ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, M8}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M9_U1 ( .a ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}), .b ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M10_U1 ( .a ({new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M9}), .b ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}), .c ({new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M10}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M11_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T15}), .clk (clk), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M12_U1 ( .a ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}), .b ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, new_AGEMA_signal_251, T27}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, M12}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M13_U1 ( .a ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, M12}), .b ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}), .c ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M14_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .b ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, M14}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M15_U1 ( .a ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, M14}), .b ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}), .c ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M16_U1 ( .a ({new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M3}), .b ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, M2}), .c ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, M16}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M17_U1 ( .a ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, new_AGEMA_signal_323, M5}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1094, new_AGEMA_signal_1092, new_AGEMA_signal_1090, new_AGEMA_signal_1088}), .c ({new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M17}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M18_U1 ( .a ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, M8}), .b ({new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M7}), .c ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, new_AGEMA_signal_359, M18}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M19_U1 ( .a ({new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M10}), .b ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}), .c ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, M19}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M20_U1 ( .a ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, M16}), .b ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}), .c ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M21_U1 ( .a ({new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M17}), .b ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}), .c ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M22_U1 ( .a ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, new_AGEMA_signal_359, M18}), .b ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}), .c ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M23_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, M19}), .b ({new_AGEMA_signal_1106, new_AGEMA_signal_1104, new_AGEMA_signal_1102, new_AGEMA_signal_1100, new_AGEMA_signal_1098}), .c ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M24_U1 ( .a ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .b ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .c ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, new_AGEMA_signal_395, M24}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M27_U1 ( .a ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .b ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .c ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C (clk), .D (new_AGEMA_signal_1067), .Q (new_AGEMA_signal_1068) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C (clk), .D (new_AGEMA_signal_1069), .Q (new_AGEMA_signal_1070) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C (clk), .D (new_AGEMA_signal_1071), .Q (new_AGEMA_signal_1072) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C (clk), .D (new_AGEMA_signal_1073), .Q (new_AGEMA_signal_1074) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C (clk), .D (new_AGEMA_signal_1075), .Q (new_AGEMA_signal_1076) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C (clk), .D (new_AGEMA_signal_1077), .Q (new_AGEMA_signal_1078) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C (clk), .D (new_AGEMA_signal_1079), .Q (new_AGEMA_signal_1080) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C (clk), .D (new_AGEMA_signal_1081), .Q (new_AGEMA_signal_1082) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C (clk), .D (new_AGEMA_signal_1083), .Q (new_AGEMA_signal_1084) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C (clk), .D (new_AGEMA_signal_1085), .Q (new_AGEMA_signal_1086) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C (clk), .D (new_AGEMA_signal_1087), .Q (new_AGEMA_signal_1088) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C (clk), .D (new_AGEMA_signal_1089), .Q (new_AGEMA_signal_1090) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C (clk), .D (new_AGEMA_signal_1091), .Q (new_AGEMA_signal_1092) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C (clk), .D (new_AGEMA_signal_1093), .Q (new_AGEMA_signal_1094) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C (clk), .D (new_AGEMA_signal_1095), .Q (new_AGEMA_signal_1096) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C (clk), .D (new_AGEMA_signal_1097), .Q (new_AGEMA_signal_1098) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C (clk), .D (new_AGEMA_signal_1099), .Q (new_AGEMA_signal_1100) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C (clk), .D (new_AGEMA_signal_1101), .Q (new_AGEMA_signal_1102) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C (clk), .D (new_AGEMA_signal_1103), .Q (new_AGEMA_signal_1104) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C (clk), .D (new_AGEMA_signal_1105), .Q (new_AGEMA_signal_1106) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C (clk), .D (new_AGEMA_signal_1187), .Q (new_AGEMA_signal_1188) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C (clk), .D (new_AGEMA_signal_1193), .Q (new_AGEMA_signal_1194) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C (clk), .D (new_AGEMA_signal_1199), .Q (new_AGEMA_signal_1200) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C (clk), .D (new_AGEMA_signal_1205), .Q (new_AGEMA_signal_1206) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C (clk), .D (new_AGEMA_signal_1211), .Q (new_AGEMA_signal_1212) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C (clk), .D (new_AGEMA_signal_1217), .Q (new_AGEMA_signal_1218) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C (clk), .D (new_AGEMA_signal_1223), .Q (new_AGEMA_signal_1224) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C (clk), .D (new_AGEMA_signal_1229), .Q (new_AGEMA_signal_1230) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C (clk), .D (new_AGEMA_signal_1235), .Q (new_AGEMA_signal_1236) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C (clk), .D (new_AGEMA_signal_1241), .Q (new_AGEMA_signal_1242) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C (clk), .D (new_AGEMA_signal_1247), .Q (new_AGEMA_signal_1248) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C (clk), .D (new_AGEMA_signal_1253), .Q (new_AGEMA_signal_1254) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C (clk), .D (new_AGEMA_signal_1259), .Q (new_AGEMA_signal_1260) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C (clk), .D (new_AGEMA_signal_1265), .Q (new_AGEMA_signal_1266) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C (clk), .D (new_AGEMA_signal_1271), .Q (new_AGEMA_signal_1272) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C (clk), .D (new_AGEMA_signal_1277), .Q (new_AGEMA_signal_1278) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C (clk), .D (new_AGEMA_signal_1283), .Q (new_AGEMA_signal_1284) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C (clk), .D (new_AGEMA_signal_1289), .Q (new_AGEMA_signal_1290) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C (clk), .D (new_AGEMA_signal_1295), .Q (new_AGEMA_signal_1296) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C (clk), .D (new_AGEMA_signal_1301), .Q (new_AGEMA_signal_1302) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C (clk), .D (new_AGEMA_signal_1307), .Q (new_AGEMA_signal_1308) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C (clk), .D (new_AGEMA_signal_1313), .Q (new_AGEMA_signal_1314) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C (clk), .D (new_AGEMA_signal_1319), .Q (new_AGEMA_signal_1320) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C (clk), .D (new_AGEMA_signal_1325), .Q (new_AGEMA_signal_1326) ) ;
    buf_clk new_AGEMA_reg_buffer_401 ( .C (clk), .D (new_AGEMA_signal_1331), .Q (new_AGEMA_signal_1332) ) ;
    buf_clk new_AGEMA_reg_buffer_407 ( .C (clk), .D (new_AGEMA_signal_1337), .Q (new_AGEMA_signal_1338) ) ;
    buf_clk new_AGEMA_reg_buffer_413 ( .C (clk), .D (new_AGEMA_signal_1343), .Q (new_AGEMA_signal_1344) ) ;
    buf_clk new_AGEMA_reg_buffer_419 ( .C (clk), .D (new_AGEMA_signal_1349), .Q (new_AGEMA_signal_1350) ) ;
    buf_clk new_AGEMA_reg_buffer_425 ( .C (clk), .D (new_AGEMA_signal_1355), .Q (new_AGEMA_signal_1356) ) ;
    buf_clk new_AGEMA_reg_buffer_431 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_1362) ) ;
    buf_clk new_AGEMA_reg_buffer_437 ( .C (clk), .D (new_AGEMA_signal_1367), .Q (new_AGEMA_signal_1368) ) ;
    buf_clk new_AGEMA_reg_buffer_443 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_1374) ) ;
    buf_clk new_AGEMA_reg_buffer_449 ( .C (clk), .D (new_AGEMA_signal_1379), .Q (new_AGEMA_signal_1380) ) ;
    buf_clk new_AGEMA_reg_buffer_455 ( .C (clk), .D (new_AGEMA_signal_1385), .Q (new_AGEMA_signal_1386) ) ;
    buf_clk new_AGEMA_reg_buffer_461 ( .C (clk), .D (new_AGEMA_signal_1391), .Q (new_AGEMA_signal_1392) ) ;
    buf_clk new_AGEMA_reg_buffer_467 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_1398) ) ;
    buf_clk new_AGEMA_reg_buffer_473 ( .C (clk), .D (new_AGEMA_signal_1403), .Q (new_AGEMA_signal_1404) ) ;
    buf_clk new_AGEMA_reg_buffer_479 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_1410) ) ;
    buf_clk new_AGEMA_reg_buffer_485 ( .C (clk), .D (new_AGEMA_signal_1415), .Q (new_AGEMA_signal_1416) ) ;
    buf_clk new_AGEMA_reg_buffer_491 ( .C (clk), .D (new_AGEMA_signal_1421), .Q (new_AGEMA_signal_1422) ) ;
    buf_clk new_AGEMA_reg_buffer_497 ( .C (clk), .D (new_AGEMA_signal_1427), .Q (new_AGEMA_signal_1428) ) ;
    buf_clk new_AGEMA_reg_buffer_503 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_1434) ) ;
    buf_clk new_AGEMA_reg_buffer_509 ( .C (clk), .D (new_AGEMA_signal_1439), .Q (new_AGEMA_signal_1440) ) ;
    buf_clk new_AGEMA_reg_buffer_515 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_1446) ) ;
    buf_clk new_AGEMA_reg_buffer_521 ( .C (clk), .D (new_AGEMA_signal_1451), .Q (new_AGEMA_signal_1452) ) ;
    buf_clk new_AGEMA_reg_buffer_527 ( .C (clk), .D (new_AGEMA_signal_1457), .Q (new_AGEMA_signal_1458) ) ;
    buf_clk new_AGEMA_reg_buffer_533 ( .C (clk), .D (new_AGEMA_signal_1463), .Q (new_AGEMA_signal_1464) ) ;
    buf_clk new_AGEMA_reg_buffer_539 ( .C (clk), .D (new_AGEMA_signal_1469), .Q (new_AGEMA_signal_1470) ) ;
    buf_clk new_AGEMA_reg_buffer_545 ( .C (clk), .D (new_AGEMA_signal_1475), .Q (new_AGEMA_signal_1476) ) ;
    buf_clk new_AGEMA_reg_buffer_551 ( .C (clk), .D (new_AGEMA_signal_1481), .Q (new_AGEMA_signal_1482) ) ;
    buf_clk new_AGEMA_reg_buffer_557 ( .C (clk), .D (new_AGEMA_signal_1487), .Q (new_AGEMA_signal_1488) ) ;
    buf_clk new_AGEMA_reg_buffer_563 ( .C (clk), .D (new_AGEMA_signal_1493), .Q (new_AGEMA_signal_1494) ) ;
    buf_clk new_AGEMA_reg_buffer_569 ( .C (clk), .D (new_AGEMA_signal_1499), .Q (new_AGEMA_signal_1500) ) ;
    buf_clk new_AGEMA_reg_buffer_575 ( .C (clk), .D (new_AGEMA_signal_1505), .Q (new_AGEMA_signal_1506) ) ;
    buf_clk new_AGEMA_reg_buffer_581 ( .C (clk), .D (new_AGEMA_signal_1511), .Q (new_AGEMA_signal_1512) ) ;
    buf_clk new_AGEMA_reg_buffer_587 ( .C (clk), .D (new_AGEMA_signal_1517), .Q (new_AGEMA_signal_1518) ) ;
    buf_clk new_AGEMA_reg_buffer_593 ( .C (clk), .D (new_AGEMA_signal_1523), .Q (new_AGEMA_signal_1524) ) ;
    buf_clk new_AGEMA_reg_buffer_599 ( .C (clk), .D (new_AGEMA_signal_1529), .Q (new_AGEMA_signal_1530) ) ;
    buf_clk new_AGEMA_reg_buffer_605 ( .C (clk), .D (new_AGEMA_signal_1535), .Q (new_AGEMA_signal_1536) ) ;
    buf_clk new_AGEMA_reg_buffer_611 ( .C (clk), .D (new_AGEMA_signal_1541), .Q (new_AGEMA_signal_1542) ) ;
    buf_clk new_AGEMA_reg_buffer_617 ( .C (clk), .D (new_AGEMA_signal_1547), .Q (new_AGEMA_signal_1548) ) ;
    buf_clk new_AGEMA_reg_buffer_623 ( .C (clk), .D (new_AGEMA_signal_1553), .Q (new_AGEMA_signal_1554) ) ;
    buf_clk new_AGEMA_reg_buffer_629 ( .C (clk), .D (new_AGEMA_signal_1559), .Q (new_AGEMA_signal_1560) ) ;
    buf_clk new_AGEMA_reg_buffer_635 ( .C (clk), .D (new_AGEMA_signal_1565), .Q (new_AGEMA_signal_1566) ) ;
    buf_clk new_AGEMA_reg_buffer_641 ( .C (clk), .D (new_AGEMA_signal_1571), .Q (new_AGEMA_signal_1572) ) ;
    buf_clk new_AGEMA_reg_buffer_647 ( .C (clk), .D (new_AGEMA_signal_1577), .Q (new_AGEMA_signal_1578) ) ;
    buf_clk new_AGEMA_reg_buffer_653 ( .C (clk), .D (new_AGEMA_signal_1583), .Q (new_AGEMA_signal_1584) ) ;
    buf_clk new_AGEMA_reg_buffer_659 ( .C (clk), .D (new_AGEMA_signal_1589), .Q (new_AGEMA_signal_1590) ) ;
    buf_clk new_AGEMA_reg_buffer_665 ( .C (clk), .D (new_AGEMA_signal_1595), .Q (new_AGEMA_signal_1596) ) ;
    buf_clk new_AGEMA_reg_buffer_671 ( .C (clk), .D (new_AGEMA_signal_1601), .Q (new_AGEMA_signal_1602) ) ;
    buf_clk new_AGEMA_reg_buffer_677 ( .C (clk), .D (new_AGEMA_signal_1607), .Q (new_AGEMA_signal_1608) ) ;
    buf_clk new_AGEMA_reg_buffer_683 ( .C (clk), .D (new_AGEMA_signal_1613), .Q (new_AGEMA_signal_1614) ) ;
    buf_clk new_AGEMA_reg_buffer_689 ( .C (clk), .D (new_AGEMA_signal_1619), .Q (new_AGEMA_signal_1620) ) ;
    buf_clk new_AGEMA_reg_buffer_695 ( .C (clk), .D (new_AGEMA_signal_1625), .Q (new_AGEMA_signal_1626) ) ;
    buf_clk new_AGEMA_reg_buffer_701 ( .C (clk), .D (new_AGEMA_signal_1631), .Q (new_AGEMA_signal_1632) ) ;
    buf_clk new_AGEMA_reg_buffer_707 ( .C (clk), .D (new_AGEMA_signal_1637), .Q (new_AGEMA_signal_1638) ) ;
    buf_clk new_AGEMA_reg_buffer_713 ( .C (clk), .D (new_AGEMA_signal_1643), .Q (new_AGEMA_signal_1644) ) ;
    buf_clk new_AGEMA_reg_buffer_719 ( .C (clk), .D (new_AGEMA_signal_1649), .Q (new_AGEMA_signal_1650) ) ;
    buf_clk new_AGEMA_reg_buffer_725 ( .C (clk), .D (new_AGEMA_signal_1655), .Q (new_AGEMA_signal_1656) ) ;
    buf_clk new_AGEMA_reg_buffer_731 ( .C (clk), .D (new_AGEMA_signal_1661), .Q (new_AGEMA_signal_1662) ) ;
    buf_clk new_AGEMA_reg_buffer_737 ( .C (clk), .D (new_AGEMA_signal_1667), .Q (new_AGEMA_signal_1668) ) ;
    buf_clk new_AGEMA_reg_buffer_743 ( .C (clk), .D (new_AGEMA_signal_1673), .Q (new_AGEMA_signal_1674) ) ;
    buf_clk new_AGEMA_reg_buffer_749 ( .C (clk), .D (new_AGEMA_signal_1679), .Q (new_AGEMA_signal_1680) ) ;
    buf_clk new_AGEMA_reg_buffer_755 ( .C (clk), .D (new_AGEMA_signal_1685), .Q (new_AGEMA_signal_1686) ) ;
    buf_clk new_AGEMA_reg_buffer_761 ( .C (clk), .D (new_AGEMA_signal_1691), .Q (new_AGEMA_signal_1692) ) ;
    buf_clk new_AGEMA_reg_buffer_767 ( .C (clk), .D (new_AGEMA_signal_1697), .Q (new_AGEMA_signal_1698) ) ;
    buf_clk new_AGEMA_reg_buffer_773 ( .C (clk), .D (new_AGEMA_signal_1703), .Q (new_AGEMA_signal_1704) ) ;
    buf_clk new_AGEMA_reg_buffer_779 ( .C (clk), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_1710) ) ;
    buf_clk new_AGEMA_reg_buffer_785 ( .C (clk), .D (new_AGEMA_signal_1715), .Q (new_AGEMA_signal_1716) ) ;
    buf_clk new_AGEMA_reg_buffer_791 ( .C (clk), .D (new_AGEMA_signal_1721), .Q (new_AGEMA_signal_1722) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_176 ( .C (clk), .D (M21), .Q (new_AGEMA_signal_1107) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C (clk), .D (new_AGEMA_signal_371), .Q (new_AGEMA_signal_1109) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C (clk), .D (new_AGEMA_signal_372), .Q (new_AGEMA_signal_1111) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C (clk), .D (new_AGEMA_signal_373), .Q (new_AGEMA_signal_1113) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C (clk), .D (new_AGEMA_signal_374), .Q (new_AGEMA_signal_1115) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C (clk), .D (M23), .Q (new_AGEMA_signal_1117) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C (clk), .D (new_AGEMA_signal_379), .Q (new_AGEMA_signal_1119) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C (clk), .D (new_AGEMA_signal_380), .Q (new_AGEMA_signal_1121) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C (clk), .D (new_AGEMA_signal_381), .Q (new_AGEMA_signal_1123) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C (clk), .D (new_AGEMA_signal_382), .Q (new_AGEMA_signal_1125) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C (clk), .D (M27), .Q (new_AGEMA_signal_1127) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C (clk), .D (new_AGEMA_signal_387), .Q (new_AGEMA_signal_1129) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C (clk), .D (new_AGEMA_signal_388), .Q (new_AGEMA_signal_1131) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C (clk), .D (new_AGEMA_signal_389), .Q (new_AGEMA_signal_1133) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C (clk), .D (new_AGEMA_signal_390), .Q (new_AGEMA_signal_1135) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C (clk), .D (M24), .Q (new_AGEMA_signal_1137) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C (clk), .D (new_AGEMA_signal_395), .Q (new_AGEMA_signal_1139) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C (clk), .D (new_AGEMA_signal_396), .Q (new_AGEMA_signal_1141) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C (clk), .D (new_AGEMA_signal_397), .Q (new_AGEMA_signal_1143) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C (clk), .D (new_AGEMA_signal_398), .Q (new_AGEMA_signal_1145) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C (clk), .D (new_AGEMA_signal_1188), .Q (new_AGEMA_signal_1189) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_1195) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C (clk), .D (new_AGEMA_signal_1200), .Q (new_AGEMA_signal_1201) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_1207) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C (clk), .D (new_AGEMA_signal_1212), .Q (new_AGEMA_signal_1213) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C (clk), .D (new_AGEMA_signal_1218), .Q (new_AGEMA_signal_1219) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C (clk), .D (new_AGEMA_signal_1224), .Q (new_AGEMA_signal_1225) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C (clk), .D (new_AGEMA_signal_1230), .Q (new_AGEMA_signal_1231) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C (clk), .D (new_AGEMA_signal_1236), .Q (new_AGEMA_signal_1237) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_1243) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C (clk), .D (new_AGEMA_signal_1248), .Q (new_AGEMA_signal_1249) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_1255) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C (clk), .D (new_AGEMA_signal_1260), .Q (new_AGEMA_signal_1261) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C (clk), .D (new_AGEMA_signal_1266), .Q (new_AGEMA_signal_1267) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C (clk), .D (new_AGEMA_signal_1272), .Q (new_AGEMA_signal_1273) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_1279) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C (clk), .D (new_AGEMA_signal_1284), .Q (new_AGEMA_signal_1285) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_1291) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C (clk), .D (new_AGEMA_signal_1296), .Q (new_AGEMA_signal_1297) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C (clk), .D (new_AGEMA_signal_1302), .Q (new_AGEMA_signal_1303) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C (clk), .D (new_AGEMA_signal_1308), .Q (new_AGEMA_signal_1309) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C (clk), .D (new_AGEMA_signal_1314), .Q (new_AGEMA_signal_1315) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C (clk), .D (new_AGEMA_signal_1320), .Q (new_AGEMA_signal_1321) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C (clk), .D (new_AGEMA_signal_1326), .Q (new_AGEMA_signal_1327) ) ;
    buf_clk new_AGEMA_reg_buffer_402 ( .C (clk), .D (new_AGEMA_signal_1332), .Q (new_AGEMA_signal_1333) ) ;
    buf_clk new_AGEMA_reg_buffer_408 ( .C (clk), .D (new_AGEMA_signal_1338), .Q (new_AGEMA_signal_1339) ) ;
    buf_clk new_AGEMA_reg_buffer_414 ( .C (clk), .D (new_AGEMA_signal_1344), .Q (new_AGEMA_signal_1345) ) ;
    buf_clk new_AGEMA_reg_buffer_420 ( .C (clk), .D (new_AGEMA_signal_1350), .Q (new_AGEMA_signal_1351) ) ;
    buf_clk new_AGEMA_reg_buffer_426 ( .C (clk), .D (new_AGEMA_signal_1356), .Q (new_AGEMA_signal_1357) ) ;
    buf_clk new_AGEMA_reg_buffer_432 ( .C (clk), .D (new_AGEMA_signal_1362), .Q (new_AGEMA_signal_1363) ) ;
    buf_clk new_AGEMA_reg_buffer_438 ( .C (clk), .D (new_AGEMA_signal_1368), .Q (new_AGEMA_signal_1369) ) ;
    buf_clk new_AGEMA_reg_buffer_444 ( .C (clk), .D (new_AGEMA_signal_1374), .Q (new_AGEMA_signal_1375) ) ;
    buf_clk new_AGEMA_reg_buffer_450 ( .C (clk), .D (new_AGEMA_signal_1380), .Q (new_AGEMA_signal_1381) ) ;
    buf_clk new_AGEMA_reg_buffer_456 ( .C (clk), .D (new_AGEMA_signal_1386), .Q (new_AGEMA_signal_1387) ) ;
    buf_clk new_AGEMA_reg_buffer_462 ( .C (clk), .D (new_AGEMA_signal_1392), .Q (new_AGEMA_signal_1393) ) ;
    buf_clk new_AGEMA_reg_buffer_468 ( .C (clk), .D (new_AGEMA_signal_1398), .Q (new_AGEMA_signal_1399) ) ;
    buf_clk new_AGEMA_reg_buffer_474 ( .C (clk), .D (new_AGEMA_signal_1404), .Q (new_AGEMA_signal_1405) ) ;
    buf_clk new_AGEMA_reg_buffer_480 ( .C (clk), .D (new_AGEMA_signal_1410), .Q (new_AGEMA_signal_1411) ) ;
    buf_clk new_AGEMA_reg_buffer_486 ( .C (clk), .D (new_AGEMA_signal_1416), .Q (new_AGEMA_signal_1417) ) ;
    buf_clk new_AGEMA_reg_buffer_492 ( .C (clk), .D (new_AGEMA_signal_1422), .Q (new_AGEMA_signal_1423) ) ;
    buf_clk new_AGEMA_reg_buffer_498 ( .C (clk), .D (new_AGEMA_signal_1428), .Q (new_AGEMA_signal_1429) ) ;
    buf_clk new_AGEMA_reg_buffer_504 ( .C (clk), .D (new_AGEMA_signal_1434), .Q (new_AGEMA_signal_1435) ) ;
    buf_clk new_AGEMA_reg_buffer_510 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_1441) ) ;
    buf_clk new_AGEMA_reg_buffer_516 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_1447) ) ;
    buf_clk new_AGEMA_reg_buffer_522 ( .C (clk), .D (new_AGEMA_signal_1452), .Q (new_AGEMA_signal_1453) ) ;
    buf_clk new_AGEMA_reg_buffer_528 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_1459) ) ;
    buf_clk new_AGEMA_reg_buffer_534 ( .C (clk), .D (new_AGEMA_signal_1464), .Q (new_AGEMA_signal_1465) ) ;
    buf_clk new_AGEMA_reg_buffer_540 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_1471) ) ;
    buf_clk new_AGEMA_reg_buffer_546 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_1477) ) ;
    buf_clk new_AGEMA_reg_buffer_552 ( .C (clk), .D (new_AGEMA_signal_1482), .Q (new_AGEMA_signal_1483) ) ;
    buf_clk new_AGEMA_reg_buffer_558 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_1489) ) ;
    buf_clk new_AGEMA_reg_buffer_564 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_1495) ) ;
    buf_clk new_AGEMA_reg_buffer_570 ( .C (clk), .D (new_AGEMA_signal_1500), .Q (new_AGEMA_signal_1501) ) ;
    buf_clk new_AGEMA_reg_buffer_576 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_1507) ) ;
    buf_clk new_AGEMA_reg_buffer_582 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_1513) ) ;
    buf_clk new_AGEMA_reg_buffer_588 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_1519) ) ;
    buf_clk new_AGEMA_reg_buffer_594 ( .C (clk), .D (new_AGEMA_signal_1524), .Q (new_AGEMA_signal_1525) ) ;
    buf_clk new_AGEMA_reg_buffer_600 ( .C (clk), .D (new_AGEMA_signal_1530), .Q (new_AGEMA_signal_1531) ) ;
    buf_clk new_AGEMA_reg_buffer_606 ( .C (clk), .D (new_AGEMA_signal_1536), .Q (new_AGEMA_signal_1537) ) ;
    buf_clk new_AGEMA_reg_buffer_612 ( .C (clk), .D (new_AGEMA_signal_1542), .Q (new_AGEMA_signal_1543) ) ;
    buf_clk new_AGEMA_reg_buffer_618 ( .C (clk), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_1549) ) ;
    buf_clk new_AGEMA_reg_buffer_624 ( .C (clk), .D (new_AGEMA_signal_1554), .Q (new_AGEMA_signal_1555) ) ;
    buf_clk new_AGEMA_reg_buffer_630 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_1561) ) ;
    buf_clk new_AGEMA_reg_buffer_636 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_1567) ) ;
    buf_clk new_AGEMA_reg_buffer_642 ( .C (clk), .D (new_AGEMA_signal_1572), .Q (new_AGEMA_signal_1573) ) ;
    buf_clk new_AGEMA_reg_buffer_648 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_1579) ) ;
    buf_clk new_AGEMA_reg_buffer_654 ( .C (clk), .D (new_AGEMA_signal_1584), .Q (new_AGEMA_signal_1585) ) ;
    buf_clk new_AGEMA_reg_buffer_660 ( .C (clk), .D (new_AGEMA_signal_1590), .Q (new_AGEMA_signal_1591) ) ;
    buf_clk new_AGEMA_reg_buffer_666 ( .C (clk), .D (new_AGEMA_signal_1596), .Q (new_AGEMA_signal_1597) ) ;
    buf_clk new_AGEMA_reg_buffer_672 ( .C (clk), .D (new_AGEMA_signal_1602), .Q (new_AGEMA_signal_1603) ) ;
    buf_clk new_AGEMA_reg_buffer_678 ( .C (clk), .D (new_AGEMA_signal_1608), .Q (new_AGEMA_signal_1609) ) ;
    buf_clk new_AGEMA_reg_buffer_684 ( .C (clk), .D (new_AGEMA_signal_1614), .Q (new_AGEMA_signal_1615) ) ;
    buf_clk new_AGEMA_reg_buffer_690 ( .C (clk), .D (new_AGEMA_signal_1620), .Q (new_AGEMA_signal_1621) ) ;
    buf_clk new_AGEMA_reg_buffer_696 ( .C (clk), .D (new_AGEMA_signal_1626), .Q (new_AGEMA_signal_1627) ) ;
    buf_clk new_AGEMA_reg_buffer_702 ( .C (clk), .D (new_AGEMA_signal_1632), .Q (new_AGEMA_signal_1633) ) ;
    buf_clk new_AGEMA_reg_buffer_708 ( .C (clk), .D (new_AGEMA_signal_1638), .Q (new_AGEMA_signal_1639) ) ;
    buf_clk new_AGEMA_reg_buffer_714 ( .C (clk), .D (new_AGEMA_signal_1644), .Q (new_AGEMA_signal_1645) ) ;
    buf_clk new_AGEMA_reg_buffer_720 ( .C (clk), .D (new_AGEMA_signal_1650), .Q (new_AGEMA_signal_1651) ) ;
    buf_clk new_AGEMA_reg_buffer_726 ( .C (clk), .D (new_AGEMA_signal_1656), .Q (new_AGEMA_signal_1657) ) ;
    buf_clk new_AGEMA_reg_buffer_732 ( .C (clk), .D (new_AGEMA_signal_1662), .Q (new_AGEMA_signal_1663) ) ;
    buf_clk new_AGEMA_reg_buffer_738 ( .C (clk), .D (new_AGEMA_signal_1668), .Q (new_AGEMA_signal_1669) ) ;
    buf_clk new_AGEMA_reg_buffer_744 ( .C (clk), .D (new_AGEMA_signal_1674), .Q (new_AGEMA_signal_1675) ) ;
    buf_clk new_AGEMA_reg_buffer_750 ( .C (clk), .D (new_AGEMA_signal_1680), .Q (new_AGEMA_signal_1681) ) ;
    buf_clk new_AGEMA_reg_buffer_756 ( .C (clk), .D (new_AGEMA_signal_1686), .Q (new_AGEMA_signal_1687) ) ;
    buf_clk new_AGEMA_reg_buffer_762 ( .C (clk), .D (new_AGEMA_signal_1692), .Q (new_AGEMA_signal_1693) ) ;
    buf_clk new_AGEMA_reg_buffer_768 ( .C (clk), .D (new_AGEMA_signal_1698), .Q (new_AGEMA_signal_1699) ) ;
    buf_clk new_AGEMA_reg_buffer_774 ( .C (clk), .D (new_AGEMA_signal_1704), .Q (new_AGEMA_signal_1705) ) ;
    buf_clk new_AGEMA_reg_buffer_780 ( .C (clk), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_1711) ) ;
    buf_clk new_AGEMA_reg_buffer_786 ( .C (clk), .D (new_AGEMA_signal_1716), .Q (new_AGEMA_signal_1717) ) ;
    buf_clk new_AGEMA_reg_buffer_792 ( .C (clk), .D (new_AGEMA_signal_1722), .Q (new_AGEMA_signal_1723) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M25_U1 ( .a ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .b ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .clk (clk), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M26_U1 ( .a ({new_AGEMA_signal_1116, new_AGEMA_signal_1114, new_AGEMA_signal_1112, new_AGEMA_signal_1110, new_AGEMA_signal_1108}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, M26}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M28_U1 ( .a ({new_AGEMA_signal_1126, new_AGEMA_signal_1124, new_AGEMA_signal_1122, new_AGEMA_signal_1120, new_AGEMA_signal_1118}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M28}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M31_U1 ( .a ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .b ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .clk (clk), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, new_AGEMA_signal_407, M31}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M33_U1 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1134, new_AGEMA_signal_1132, new_AGEMA_signal_1130, new_AGEMA_signal_1128}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, M33}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M34_U1 ( .a ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .b ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M34}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M36_U1 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1144, new_AGEMA_signal_1142, new_AGEMA_signal_1140, new_AGEMA_signal_1138}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, new_AGEMA_signal_431, M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C (clk), .D (new_AGEMA_signal_1107), .Q (new_AGEMA_signal_1108) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C (clk), .D (new_AGEMA_signal_1109), .Q (new_AGEMA_signal_1110) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C (clk), .D (new_AGEMA_signal_1111), .Q (new_AGEMA_signal_1112) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C (clk), .D (new_AGEMA_signal_1113), .Q (new_AGEMA_signal_1114) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C (clk), .D (new_AGEMA_signal_1115), .Q (new_AGEMA_signal_1116) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C (clk), .D (new_AGEMA_signal_1117), .Q (new_AGEMA_signal_1118) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C (clk), .D (new_AGEMA_signal_1119), .Q (new_AGEMA_signal_1120) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C (clk), .D (new_AGEMA_signal_1121), .Q (new_AGEMA_signal_1122) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C (clk), .D (new_AGEMA_signal_1123), .Q (new_AGEMA_signal_1124) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C (clk), .D (new_AGEMA_signal_1125), .Q (new_AGEMA_signal_1126) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C (clk), .D (new_AGEMA_signal_1127), .Q (new_AGEMA_signal_1128) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C (clk), .D (new_AGEMA_signal_1129), .Q (new_AGEMA_signal_1130) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C (clk), .D (new_AGEMA_signal_1131), .Q (new_AGEMA_signal_1132) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C (clk), .D (new_AGEMA_signal_1133), .Q (new_AGEMA_signal_1134) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C (clk), .D (new_AGEMA_signal_1135), .Q (new_AGEMA_signal_1136) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C (clk), .D (new_AGEMA_signal_1137), .Q (new_AGEMA_signal_1138) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C (clk), .D (new_AGEMA_signal_1139), .Q (new_AGEMA_signal_1140) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C (clk), .D (new_AGEMA_signal_1141), .Q (new_AGEMA_signal_1142) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C (clk), .D (new_AGEMA_signal_1143), .Q (new_AGEMA_signal_1144) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C (clk), .D (new_AGEMA_signal_1145), .Q (new_AGEMA_signal_1146) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C (clk), .D (new_AGEMA_signal_1189), .Q (new_AGEMA_signal_1190) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C (clk), .D (new_AGEMA_signal_1195), .Q (new_AGEMA_signal_1196) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C (clk), .D (new_AGEMA_signal_1201), .Q (new_AGEMA_signal_1202) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C (clk), .D (new_AGEMA_signal_1207), .Q (new_AGEMA_signal_1208) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C (clk), .D (new_AGEMA_signal_1213), .Q (new_AGEMA_signal_1214) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C (clk), .D (new_AGEMA_signal_1219), .Q (new_AGEMA_signal_1220) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C (clk), .D (new_AGEMA_signal_1225), .Q (new_AGEMA_signal_1226) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C (clk), .D (new_AGEMA_signal_1231), .Q (new_AGEMA_signal_1232) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C (clk), .D (new_AGEMA_signal_1237), .Q (new_AGEMA_signal_1238) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C (clk), .D (new_AGEMA_signal_1243), .Q (new_AGEMA_signal_1244) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C (clk), .D (new_AGEMA_signal_1249), .Q (new_AGEMA_signal_1250) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C (clk), .D (new_AGEMA_signal_1255), .Q (new_AGEMA_signal_1256) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C (clk), .D (new_AGEMA_signal_1261), .Q (new_AGEMA_signal_1262) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C (clk), .D (new_AGEMA_signal_1267), .Q (new_AGEMA_signal_1268) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C (clk), .D (new_AGEMA_signal_1273), .Q (new_AGEMA_signal_1274) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C (clk), .D (new_AGEMA_signal_1279), .Q (new_AGEMA_signal_1280) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C (clk), .D (new_AGEMA_signal_1285), .Q (new_AGEMA_signal_1286) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C (clk), .D (new_AGEMA_signal_1291), .Q (new_AGEMA_signal_1292) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C (clk), .D (new_AGEMA_signal_1297), .Q (new_AGEMA_signal_1298) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C (clk), .D (new_AGEMA_signal_1303), .Q (new_AGEMA_signal_1304) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C (clk), .D (new_AGEMA_signal_1309), .Q (new_AGEMA_signal_1310) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C (clk), .D (new_AGEMA_signal_1315), .Q (new_AGEMA_signal_1316) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C (clk), .D (new_AGEMA_signal_1321), .Q (new_AGEMA_signal_1322) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C (clk), .D (new_AGEMA_signal_1327), .Q (new_AGEMA_signal_1328) ) ;
    buf_clk new_AGEMA_reg_buffer_403 ( .C (clk), .D (new_AGEMA_signal_1333), .Q (new_AGEMA_signal_1334) ) ;
    buf_clk new_AGEMA_reg_buffer_409 ( .C (clk), .D (new_AGEMA_signal_1339), .Q (new_AGEMA_signal_1340) ) ;
    buf_clk new_AGEMA_reg_buffer_415 ( .C (clk), .D (new_AGEMA_signal_1345), .Q (new_AGEMA_signal_1346) ) ;
    buf_clk new_AGEMA_reg_buffer_421 ( .C (clk), .D (new_AGEMA_signal_1351), .Q (new_AGEMA_signal_1352) ) ;
    buf_clk new_AGEMA_reg_buffer_427 ( .C (clk), .D (new_AGEMA_signal_1357), .Q (new_AGEMA_signal_1358) ) ;
    buf_clk new_AGEMA_reg_buffer_433 ( .C (clk), .D (new_AGEMA_signal_1363), .Q (new_AGEMA_signal_1364) ) ;
    buf_clk new_AGEMA_reg_buffer_439 ( .C (clk), .D (new_AGEMA_signal_1369), .Q (new_AGEMA_signal_1370) ) ;
    buf_clk new_AGEMA_reg_buffer_445 ( .C (clk), .D (new_AGEMA_signal_1375), .Q (new_AGEMA_signal_1376) ) ;
    buf_clk new_AGEMA_reg_buffer_451 ( .C (clk), .D (new_AGEMA_signal_1381), .Q (new_AGEMA_signal_1382) ) ;
    buf_clk new_AGEMA_reg_buffer_457 ( .C (clk), .D (new_AGEMA_signal_1387), .Q (new_AGEMA_signal_1388) ) ;
    buf_clk new_AGEMA_reg_buffer_463 ( .C (clk), .D (new_AGEMA_signal_1393), .Q (new_AGEMA_signal_1394) ) ;
    buf_clk new_AGEMA_reg_buffer_469 ( .C (clk), .D (new_AGEMA_signal_1399), .Q (new_AGEMA_signal_1400) ) ;
    buf_clk new_AGEMA_reg_buffer_475 ( .C (clk), .D (new_AGEMA_signal_1405), .Q (new_AGEMA_signal_1406) ) ;
    buf_clk new_AGEMA_reg_buffer_481 ( .C (clk), .D (new_AGEMA_signal_1411), .Q (new_AGEMA_signal_1412) ) ;
    buf_clk new_AGEMA_reg_buffer_487 ( .C (clk), .D (new_AGEMA_signal_1417), .Q (new_AGEMA_signal_1418) ) ;
    buf_clk new_AGEMA_reg_buffer_493 ( .C (clk), .D (new_AGEMA_signal_1423), .Q (new_AGEMA_signal_1424) ) ;
    buf_clk new_AGEMA_reg_buffer_499 ( .C (clk), .D (new_AGEMA_signal_1429), .Q (new_AGEMA_signal_1430) ) ;
    buf_clk new_AGEMA_reg_buffer_505 ( .C (clk), .D (new_AGEMA_signal_1435), .Q (new_AGEMA_signal_1436) ) ;
    buf_clk new_AGEMA_reg_buffer_511 ( .C (clk), .D (new_AGEMA_signal_1441), .Q (new_AGEMA_signal_1442) ) ;
    buf_clk new_AGEMA_reg_buffer_517 ( .C (clk), .D (new_AGEMA_signal_1447), .Q (new_AGEMA_signal_1448) ) ;
    buf_clk new_AGEMA_reg_buffer_523 ( .C (clk), .D (new_AGEMA_signal_1453), .Q (new_AGEMA_signal_1454) ) ;
    buf_clk new_AGEMA_reg_buffer_529 ( .C (clk), .D (new_AGEMA_signal_1459), .Q (new_AGEMA_signal_1460) ) ;
    buf_clk new_AGEMA_reg_buffer_535 ( .C (clk), .D (new_AGEMA_signal_1465), .Q (new_AGEMA_signal_1466) ) ;
    buf_clk new_AGEMA_reg_buffer_541 ( .C (clk), .D (new_AGEMA_signal_1471), .Q (new_AGEMA_signal_1472) ) ;
    buf_clk new_AGEMA_reg_buffer_547 ( .C (clk), .D (new_AGEMA_signal_1477), .Q (new_AGEMA_signal_1478) ) ;
    buf_clk new_AGEMA_reg_buffer_553 ( .C (clk), .D (new_AGEMA_signal_1483), .Q (new_AGEMA_signal_1484) ) ;
    buf_clk new_AGEMA_reg_buffer_559 ( .C (clk), .D (new_AGEMA_signal_1489), .Q (new_AGEMA_signal_1490) ) ;
    buf_clk new_AGEMA_reg_buffer_565 ( .C (clk), .D (new_AGEMA_signal_1495), .Q (new_AGEMA_signal_1496) ) ;
    buf_clk new_AGEMA_reg_buffer_571 ( .C (clk), .D (new_AGEMA_signal_1501), .Q (new_AGEMA_signal_1502) ) ;
    buf_clk new_AGEMA_reg_buffer_577 ( .C (clk), .D (new_AGEMA_signal_1507), .Q (new_AGEMA_signal_1508) ) ;
    buf_clk new_AGEMA_reg_buffer_583 ( .C (clk), .D (new_AGEMA_signal_1513), .Q (new_AGEMA_signal_1514) ) ;
    buf_clk new_AGEMA_reg_buffer_589 ( .C (clk), .D (new_AGEMA_signal_1519), .Q (new_AGEMA_signal_1520) ) ;
    buf_clk new_AGEMA_reg_buffer_595 ( .C (clk), .D (new_AGEMA_signal_1525), .Q (new_AGEMA_signal_1526) ) ;
    buf_clk new_AGEMA_reg_buffer_601 ( .C (clk), .D (new_AGEMA_signal_1531), .Q (new_AGEMA_signal_1532) ) ;
    buf_clk new_AGEMA_reg_buffer_607 ( .C (clk), .D (new_AGEMA_signal_1537), .Q (new_AGEMA_signal_1538) ) ;
    buf_clk new_AGEMA_reg_buffer_613 ( .C (clk), .D (new_AGEMA_signal_1543), .Q (new_AGEMA_signal_1544) ) ;
    buf_clk new_AGEMA_reg_buffer_619 ( .C (clk), .D (new_AGEMA_signal_1549), .Q (new_AGEMA_signal_1550) ) ;
    buf_clk new_AGEMA_reg_buffer_625 ( .C (clk), .D (new_AGEMA_signal_1555), .Q (new_AGEMA_signal_1556) ) ;
    buf_clk new_AGEMA_reg_buffer_631 ( .C (clk), .D (new_AGEMA_signal_1561), .Q (new_AGEMA_signal_1562) ) ;
    buf_clk new_AGEMA_reg_buffer_637 ( .C (clk), .D (new_AGEMA_signal_1567), .Q (new_AGEMA_signal_1568) ) ;
    buf_clk new_AGEMA_reg_buffer_643 ( .C (clk), .D (new_AGEMA_signal_1573), .Q (new_AGEMA_signal_1574) ) ;
    buf_clk new_AGEMA_reg_buffer_649 ( .C (clk), .D (new_AGEMA_signal_1579), .Q (new_AGEMA_signal_1580) ) ;
    buf_clk new_AGEMA_reg_buffer_655 ( .C (clk), .D (new_AGEMA_signal_1585), .Q (new_AGEMA_signal_1586) ) ;
    buf_clk new_AGEMA_reg_buffer_661 ( .C (clk), .D (new_AGEMA_signal_1591), .Q (new_AGEMA_signal_1592) ) ;
    buf_clk new_AGEMA_reg_buffer_667 ( .C (clk), .D (new_AGEMA_signal_1597), .Q (new_AGEMA_signal_1598) ) ;
    buf_clk new_AGEMA_reg_buffer_673 ( .C (clk), .D (new_AGEMA_signal_1603), .Q (new_AGEMA_signal_1604) ) ;
    buf_clk new_AGEMA_reg_buffer_679 ( .C (clk), .D (new_AGEMA_signal_1609), .Q (new_AGEMA_signal_1610) ) ;
    buf_clk new_AGEMA_reg_buffer_685 ( .C (clk), .D (new_AGEMA_signal_1615), .Q (new_AGEMA_signal_1616) ) ;
    buf_clk new_AGEMA_reg_buffer_691 ( .C (clk), .D (new_AGEMA_signal_1621), .Q (new_AGEMA_signal_1622) ) ;
    buf_clk new_AGEMA_reg_buffer_697 ( .C (clk), .D (new_AGEMA_signal_1627), .Q (new_AGEMA_signal_1628) ) ;
    buf_clk new_AGEMA_reg_buffer_703 ( .C (clk), .D (new_AGEMA_signal_1633), .Q (new_AGEMA_signal_1634) ) ;
    buf_clk new_AGEMA_reg_buffer_709 ( .C (clk), .D (new_AGEMA_signal_1639), .Q (new_AGEMA_signal_1640) ) ;
    buf_clk new_AGEMA_reg_buffer_715 ( .C (clk), .D (new_AGEMA_signal_1645), .Q (new_AGEMA_signal_1646) ) ;
    buf_clk new_AGEMA_reg_buffer_721 ( .C (clk), .D (new_AGEMA_signal_1651), .Q (new_AGEMA_signal_1652) ) ;
    buf_clk new_AGEMA_reg_buffer_727 ( .C (clk), .D (new_AGEMA_signal_1657), .Q (new_AGEMA_signal_1658) ) ;
    buf_clk new_AGEMA_reg_buffer_733 ( .C (clk), .D (new_AGEMA_signal_1663), .Q (new_AGEMA_signal_1664) ) ;
    buf_clk new_AGEMA_reg_buffer_739 ( .C (clk), .D (new_AGEMA_signal_1669), .Q (new_AGEMA_signal_1670) ) ;
    buf_clk new_AGEMA_reg_buffer_745 ( .C (clk), .D (new_AGEMA_signal_1675), .Q (new_AGEMA_signal_1676) ) ;
    buf_clk new_AGEMA_reg_buffer_751 ( .C (clk), .D (new_AGEMA_signal_1681), .Q (new_AGEMA_signal_1682) ) ;
    buf_clk new_AGEMA_reg_buffer_757 ( .C (clk), .D (new_AGEMA_signal_1687), .Q (new_AGEMA_signal_1688) ) ;
    buf_clk new_AGEMA_reg_buffer_763 ( .C (clk), .D (new_AGEMA_signal_1693), .Q (new_AGEMA_signal_1694) ) ;
    buf_clk new_AGEMA_reg_buffer_769 ( .C (clk), .D (new_AGEMA_signal_1699), .Q (new_AGEMA_signal_1700) ) ;
    buf_clk new_AGEMA_reg_buffer_775 ( .C (clk), .D (new_AGEMA_signal_1705), .Q (new_AGEMA_signal_1706) ) ;
    buf_clk new_AGEMA_reg_buffer_781 ( .C (clk), .D (new_AGEMA_signal_1711), .Q (new_AGEMA_signal_1712) ) ;
    buf_clk new_AGEMA_reg_buffer_787 ( .C (clk), .D (new_AGEMA_signal_1717), .Q (new_AGEMA_signal_1718) ) ;
    buf_clk new_AGEMA_reg_buffer_793 ( .C (clk), .D (new_AGEMA_signal_1723), .Q (new_AGEMA_signal_1724) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_216 ( .C (clk), .D (new_AGEMA_signal_1108), .Q (new_AGEMA_signal_1147) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C (clk), .D (new_AGEMA_signal_1110), .Q (new_AGEMA_signal_1149) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C (clk), .D (new_AGEMA_signal_1112), .Q (new_AGEMA_signal_1151) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C (clk), .D (new_AGEMA_signal_1114), .Q (new_AGEMA_signal_1153) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C (clk), .D (new_AGEMA_signal_1116), .Q (new_AGEMA_signal_1155) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C (clk), .D (M33), .Q (new_AGEMA_signal_1157) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C (clk), .D (new_AGEMA_signal_411), .Q (new_AGEMA_signal_1159) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C (clk), .D (new_AGEMA_signal_412), .Q (new_AGEMA_signal_1161) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C (clk), .D (new_AGEMA_signal_413), .Q (new_AGEMA_signal_1163) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C (clk), .D (new_AGEMA_signal_414), .Q (new_AGEMA_signal_1165) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C (clk), .D (new_AGEMA_signal_1118), .Q (new_AGEMA_signal_1167) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C (clk), .D (new_AGEMA_signal_1120), .Q (new_AGEMA_signal_1169) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C (clk), .D (new_AGEMA_signal_1122), .Q (new_AGEMA_signal_1171) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C (clk), .D (new_AGEMA_signal_1124), .Q (new_AGEMA_signal_1173) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C (clk), .D (new_AGEMA_signal_1126), .Q (new_AGEMA_signal_1175) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C (clk), .D (M36), .Q (new_AGEMA_signal_1177) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C (clk), .D (new_AGEMA_signal_431), .Q (new_AGEMA_signal_1179) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C (clk), .D (new_AGEMA_signal_432), .Q (new_AGEMA_signal_1181) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C (clk), .D (new_AGEMA_signal_433), .Q (new_AGEMA_signal_1183) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C (clk), .D (new_AGEMA_signal_434), .Q (new_AGEMA_signal_1185) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C (clk), .D (new_AGEMA_signal_1190), .Q (new_AGEMA_signal_1191) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C (clk), .D (new_AGEMA_signal_1196), .Q (new_AGEMA_signal_1197) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C (clk), .D (new_AGEMA_signal_1202), .Q (new_AGEMA_signal_1203) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C (clk), .D (new_AGEMA_signal_1208), .Q (new_AGEMA_signal_1209) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C (clk), .D (new_AGEMA_signal_1214), .Q (new_AGEMA_signal_1215) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C (clk), .D (new_AGEMA_signal_1220), .Q (new_AGEMA_signal_1221) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C (clk), .D (new_AGEMA_signal_1226), .Q (new_AGEMA_signal_1227) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C (clk), .D (new_AGEMA_signal_1232), .Q (new_AGEMA_signal_1233) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C (clk), .D (new_AGEMA_signal_1238), .Q (new_AGEMA_signal_1239) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C (clk), .D (new_AGEMA_signal_1244), .Q (new_AGEMA_signal_1245) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C (clk), .D (new_AGEMA_signal_1250), .Q (new_AGEMA_signal_1251) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C (clk), .D (new_AGEMA_signal_1256), .Q (new_AGEMA_signal_1257) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C (clk), .D (new_AGEMA_signal_1262), .Q (new_AGEMA_signal_1263) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C (clk), .D (new_AGEMA_signal_1268), .Q (new_AGEMA_signal_1269) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C (clk), .D (new_AGEMA_signal_1274), .Q (new_AGEMA_signal_1275) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C (clk), .D (new_AGEMA_signal_1280), .Q (new_AGEMA_signal_1281) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C (clk), .D (new_AGEMA_signal_1286), .Q (new_AGEMA_signal_1287) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C (clk), .D (new_AGEMA_signal_1292), .Q (new_AGEMA_signal_1293) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C (clk), .D (new_AGEMA_signal_1298), .Q (new_AGEMA_signal_1299) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C (clk), .D (new_AGEMA_signal_1304), .Q (new_AGEMA_signal_1305) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C (clk), .D (new_AGEMA_signal_1310), .Q (new_AGEMA_signal_1311) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C (clk), .D (new_AGEMA_signal_1316), .Q (new_AGEMA_signal_1317) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C (clk), .D (new_AGEMA_signal_1322), .Q (new_AGEMA_signal_1323) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C (clk), .D (new_AGEMA_signal_1328), .Q (new_AGEMA_signal_1329) ) ;
    buf_clk new_AGEMA_reg_buffer_404 ( .C (clk), .D (new_AGEMA_signal_1334), .Q (new_AGEMA_signal_1335) ) ;
    buf_clk new_AGEMA_reg_buffer_410 ( .C (clk), .D (new_AGEMA_signal_1340), .Q (new_AGEMA_signal_1341) ) ;
    buf_clk new_AGEMA_reg_buffer_416 ( .C (clk), .D (new_AGEMA_signal_1346), .Q (new_AGEMA_signal_1347) ) ;
    buf_clk new_AGEMA_reg_buffer_422 ( .C (clk), .D (new_AGEMA_signal_1352), .Q (new_AGEMA_signal_1353) ) ;
    buf_clk new_AGEMA_reg_buffer_428 ( .C (clk), .D (new_AGEMA_signal_1358), .Q (new_AGEMA_signal_1359) ) ;
    buf_clk new_AGEMA_reg_buffer_434 ( .C (clk), .D (new_AGEMA_signal_1364), .Q (new_AGEMA_signal_1365) ) ;
    buf_clk new_AGEMA_reg_buffer_440 ( .C (clk), .D (new_AGEMA_signal_1370), .Q (new_AGEMA_signal_1371) ) ;
    buf_clk new_AGEMA_reg_buffer_446 ( .C (clk), .D (new_AGEMA_signal_1376), .Q (new_AGEMA_signal_1377) ) ;
    buf_clk new_AGEMA_reg_buffer_452 ( .C (clk), .D (new_AGEMA_signal_1382), .Q (new_AGEMA_signal_1383) ) ;
    buf_clk new_AGEMA_reg_buffer_458 ( .C (clk), .D (new_AGEMA_signal_1388), .Q (new_AGEMA_signal_1389) ) ;
    buf_clk new_AGEMA_reg_buffer_464 ( .C (clk), .D (new_AGEMA_signal_1394), .Q (new_AGEMA_signal_1395) ) ;
    buf_clk new_AGEMA_reg_buffer_470 ( .C (clk), .D (new_AGEMA_signal_1400), .Q (new_AGEMA_signal_1401) ) ;
    buf_clk new_AGEMA_reg_buffer_476 ( .C (clk), .D (new_AGEMA_signal_1406), .Q (new_AGEMA_signal_1407) ) ;
    buf_clk new_AGEMA_reg_buffer_482 ( .C (clk), .D (new_AGEMA_signal_1412), .Q (new_AGEMA_signal_1413) ) ;
    buf_clk new_AGEMA_reg_buffer_488 ( .C (clk), .D (new_AGEMA_signal_1418), .Q (new_AGEMA_signal_1419) ) ;
    buf_clk new_AGEMA_reg_buffer_494 ( .C (clk), .D (new_AGEMA_signal_1424), .Q (new_AGEMA_signal_1425) ) ;
    buf_clk new_AGEMA_reg_buffer_500 ( .C (clk), .D (new_AGEMA_signal_1430), .Q (new_AGEMA_signal_1431) ) ;
    buf_clk new_AGEMA_reg_buffer_506 ( .C (clk), .D (new_AGEMA_signal_1436), .Q (new_AGEMA_signal_1437) ) ;
    buf_clk new_AGEMA_reg_buffer_512 ( .C (clk), .D (new_AGEMA_signal_1442), .Q (new_AGEMA_signal_1443) ) ;
    buf_clk new_AGEMA_reg_buffer_518 ( .C (clk), .D (new_AGEMA_signal_1448), .Q (new_AGEMA_signal_1449) ) ;
    buf_clk new_AGEMA_reg_buffer_524 ( .C (clk), .D (new_AGEMA_signal_1454), .Q (new_AGEMA_signal_1455) ) ;
    buf_clk new_AGEMA_reg_buffer_530 ( .C (clk), .D (new_AGEMA_signal_1460), .Q (new_AGEMA_signal_1461) ) ;
    buf_clk new_AGEMA_reg_buffer_536 ( .C (clk), .D (new_AGEMA_signal_1466), .Q (new_AGEMA_signal_1467) ) ;
    buf_clk new_AGEMA_reg_buffer_542 ( .C (clk), .D (new_AGEMA_signal_1472), .Q (new_AGEMA_signal_1473) ) ;
    buf_clk new_AGEMA_reg_buffer_548 ( .C (clk), .D (new_AGEMA_signal_1478), .Q (new_AGEMA_signal_1479) ) ;
    buf_clk new_AGEMA_reg_buffer_554 ( .C (clk), .D (new_AGEMA_signal_1484), .Q (new_AGEMA_signal_1485) ) ;
    buf_clk new_AGEMA_reg_buffer_560 ( .C (clk), .D (new_AGEMA_signal_1490), .Q (new_AGEMA_signal_1491) ) ;
    buf_clk new_AGEMA_reg_buffer_566 ( .C (clk), .D (new_AGEMA_signal_1496), .Q (new_AGEMA_signal_1497) ) ;
    buf_clk new_AGEMA_reg_buffer_572 ( .C (clk), .D (new_AGEMA_signal_1502), .Q (new_AGEMA_signal_1503) ) ;
    buf_clk new_AGEMA_reg_buffer_578 ( .C (clk), .D (new_AGEMA_signal_1508), .Q (new_AGEMA_signal_1509) ) ;
    buf_clk new_AGEMA_reg_buffer_584 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_1515) ) ;
    buf_clk new_AGEMA_reg_buffer_590 ( .C (clk), .D (new_AGEMA_signal_1520), .Q (new_AGEMA_signal_1521) ) ;
    buf_clk new_AGEMA_reg_buffer_596 ( .C (clk), .D (new_AGEMA_signal_1526), .Q (new_AGEMA_signal_1527) ) ;
    buf_clk new_AGEMA_reg_buffer_602 ( .C (clk), .D (new_AGEMA_signal_1532), .Q (new_AGEMA_signal_1533) ) ;
    buf_clk new_AGEMA_reg_buffer_608 ( .C (clk), .D (new_AGEMA_signal_1538), .Q (new_AGEMA_signal_1539) ) ;
    buf_clk new_AGEMA_reg_buffer_614 ( .C (clk), .D (new_AGEMA_signal_1544), .Q (new_AGEMA_signal_1545) ) ;
    buf_clk new_AGEMA_reg_buffer_620 ( .C (clk), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_1551) ) ;
    buf_clk new_AGEMA_reg_buffer_626 ( .C (clk), .D (new_AGEMA_signal_1556), .Q (new_AGEMA_signal_1557) ) ;
    buf_clk new_AGEMA_reg_buffer_632 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_1563) ) ;
    buf_clk new_AGEMA_reg_buffer_638 ( .C (clk), .D (new_AGEMA_signal_1568), .Q (new_AGEMA_signal_1569) ) ;
    buf_clk new_AGEMA_reg_buffer_644 ( .C (clk), .D (new_AGEMA_signal_1574), .Q (new_AGEMA_signal_1575) ) ;
    buf_clk new_AGEMA_reg_buffer_650 ( .C (clk), .D (new_AGEMA_signal_1580), .Q (new_AGEMA_signal_1581) ) ;
    buf_clk new_AGEMA_reg_buffer_656 ( .C (clk), .D (new_AGEMA_signal_1586), .Q (new_AGEMA_signal_1587) ) ;
    buf_clk new_AGEMA_reg_buffer_662 ( .C (clk), .D (new_AGEMA_signal_1592), .Q (new_AGEMA_signal_1593) ) ;
    buf_clk new_AGEMA_reg_buffer_668 ( .C (clk), .D (new_AGEMA_signal_1598), .Q (new_AGEMA_signal_1599) ) ;
    buf_clk new_AGEMA_reg_buffer_674 ( .C (clk), .D (new_AGEMA_signal_1604), .Q (new_AGEMA_signal_1605) ) ;
    buf_clk new_AGEMA_reg_buffer_680 ( .C (clk), .D (new_AGEMA_signal_1610), .Q (new_AGEMA_signal_1611) ) ;
    buf_clk new_AGEMA_reg_buffer_686 ( .C (clk), .D (new_AGEMA_signal_1616), .Q (new_AGEMA_signal_1617) ) ;
    buf_clk new_AGEMA_reg_buffer_692 ( .C (clk), .D (new_AGEMA_signal_1622), .Q (new_AGEMA_signal_1623) ) ;
    buf_clk new_AGEMA_reg_buffer_698 ( .C (clk), .D (new_AGEMA_signal_1628), .Q (new_AGEMA_signal_1629) ) ;
    buf_clk new_AGEMA_reg_buffer_704 ( .C (clk), .D (new_AGEMA_signal_1634), .Q (new_AGEMA_signal_1635) ) ;
    buf_clk new_AGEMA_reg_buffer_710 ( .C (clk), .D (new_AGEMA_signal_1640), .Q (new_AGEMA_signal_1641) ) ;
    buf_clk new_AGEMA_reg_buffer_716 ( .C (clk), .D (new_AGEMA_signal_1646), .Q (new_AGEMA_signal_1647) ) ;
    buf_clk new_AGEMA_reg_buffer_722 ( .C (clk), .D (new_AGEMA_signal_1652), .Q (new_AGEMA_signal_1653) ) ;
    buf_clk new_AGEMA_reg_buffer_728 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_1659) ) ;
    buf_clk new_AGEMA_reg_buffer_734 ( .C (clk), .D (new_AGEMA_signal_1664), .Q (new_AGEMA_signal_1665) ) ;
    buf_clk new_AGEMA_reg_buffer_740 ( .C (clk), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_1671) ) ;
    buf_clk new_AGEMA_reg_buffer_746 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_1677) ) ;
    buf_clk new_AGEMA_reg_buffer_752 ( .C (clk), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_1683) ) ;
    buf_clk new_AGEMA_reg_buffer_758 ( .C (clk), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_1689) ) ;
    buf_clk new_AGEMA_reg_buffer_764 ( .C (clk), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_1695) ) ;
    buf_clk new_AGEMA_reg_buffer_770 ( .C (clk), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_1701) ) ;
    buf_clk new_AGEMA_reg_buffer_776 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_1707) ) ;
    buf_clk new_AGEMA_reg_buffer_782 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_1713) ) ;
    buf_clk new_AGEMA_reg_buffer_788 ( .C (clk), .D (new_AGEMA_signal_1718), .Q (new_AGEMA_signal_1719) ) ;
    buf_clk new_AGEMA_reg_buffer_794 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_1725) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M29_U1 ( .a ({new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M28}), .b ({new_AGEMA_signal_1136, new_AGEMA_signal_1134, new_AGEMA_signal_1132, new_AGEMA_signal_1130, new_AGEMA_signal_1128}), .clk (clk), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M29}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M30_U1 ( .a ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, M26}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1144, new_AGEMA_signal_1142, new_AGEMA_signal_1140, new_AGEMA_signal_1138}), .clk (clk), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, new_AGEMA_signal_419, M30}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M32_U1 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1134, new_AGEMA_signal_1132, new_AGEMA_signal_1130, new_AGEMA_signal_1128}), .b ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, new_AGEMA_signal_407, M31}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, M32}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M35_U1 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1144, new_AGEMA_signal_1142, new_AGEMA_signal_1140, new_AGEMA_signal_1138}), .b ({new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M34}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M35}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M37_U1 ( .a ({new_AGEMA_signal_1156, new_AGEMA_signal_1154, new_AGEMA_signal_1152, new_AGEMA_signal_1150, new_AGEMA_signal_1148}), .b ({new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M29}), .c ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M38_U1 ( .a ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, M32}), .b ({new_AGEMA_signal_1166, new_AGEMA_signal_1164, new_AGEMA_signal_1162, new_AGEMA_signal_1160, new_AGEMA_signal_1158}), .c ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M39_U1 ( .a ({new_AGEMA_signal_1176, new_AGEMA_signal_1174, new_AGEMA_signal_1172, new_AGEMA_signal_1170, new_AGEMA_signal_1168}), .b ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, new_AGEMA_signal_419, M30}), .c ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M40_U1 ( .a ({new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M35}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1184, new_AGEMA_signal_1182, new_AGEMA_signal_1180, new_AGEMA_signal_1178}), .c ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M41_U1 ( .a ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .c ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M42_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .c ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M43_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .c ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M44_U1 ( .a ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .c ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_M45_U1 ( .a ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .b ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .c ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C (clk), .D (new_AGEMA_signal_1147), .Q (new_AGEMA_signal_1148) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C (clk), .D (new_AGEMA_signal_1149), .Q (new_AGEMA_signal_1150) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C (clk), .D (new_AGEMA_signal_1151), .Q (new_AGEMA_signal_1152) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C (clk), .D (new_AGEMA_signal_1153), .Q (new_AGEMA_signal_1154) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C (clk), .D (new_AGEMA_signal_1155), .Q (new_AGEMA_signal_1156) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C (clk), .D (new_AGEMA_signal_1157), .Q (new_AGEMA_signal_1158) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C (clk), .D (new_AGEMA_signal_1159), .Q (new_AGEMA_signal_1160) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C (clk), .D (new_AGEMA_signal_1161), .Q (new_AGEMA_signal_1162) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C (clk), .D (new_AGEMA_signal_1163), .Q (new_AGEMA_signal_1164) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C (clk), .D (new_AGEMA_signal_1165), .Q (new_AGEMA_signal_1166) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C (clk), .D (new_AGEMA_signal_1167), .Q (new_AGEMA_signal_1168) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C (clk), .D (new_AGEMA_signal_1169), .Q (new_AGEMA_signal_1170) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C (clk), .D (new_AGEMA_signal_1171), .Q (new_AGEMA_signal_1172) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C (clk), .D (new_AGEMA_signal_1173), .Q (new_AGEMA_signal_1174) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C (clk), .D (new_AGEMA_signal_1175), .Q (new_AGEMA_signal_1176) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C (clk), .D (new_AGEMA_signal_1177), .Q (new_AGEMA_signal_1178) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C (clk), .D (new_AGEMA_signal_1179), .Q (new_AGEMA_signal_1180) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C (clk), .D (new_AGEMA_signal_1181), .Q (new_AGEMA_signal_1182) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C (clk), .D (new_AGEMA_signal_1183), .Q (new_AGEMA_signal_1184) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C (clk), .D (new_AGEMA_signal_1185), .Q (new_AGEMA_signal_1186) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C (clk), .D (new_AGEMA_signal_1191), .Q (new_AGEMA_signal_1192) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C (clk), .D (new_AGEMA_signal_1197), .Q (new_AGEMA_signal_1198) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C (clk), .D (new_AGEMA_signal_1203), .Q (new_AGEMA_signal_1204) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C (clk), .D (new_AGEMA_signal_1209), .Q (new_AGEMA_signal_1210) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C (clk), .D (new_AGEMA_signal_1215), .Q (new_AGEMA_signal_1216) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C (clk), .D (new_AGEMA_signal_1221), .Q (new_AGEMA_signal_1222) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C (clk), .D (new_AGEMA_signal_1227), .Q (new_AGEMA_signal_1228) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C (clk), .D (new_AGEMA_signal_1233), .Q (new_AGEMA_signal_1234) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C (clk), .D (new_AGEMA_signal_1239), .Q (new_AGEMA_signal_1240) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C (clk), .D (new_AGEMA_signal_1245), .Q (new_AGEMA_signal_1246) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C (clk), .D (new_AGEMA_signal_1251), .Q (new_AGEMA_signal_1252) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C (clk), .D (new_AGEMA_signal_1257), .Q (new_AGEMA_signal_1258) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C (clk), .D (new_AGEMA_signal_1263), .Q (new_AGEMA_signal_1264) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_1270) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C (clk), .D (new_AGEMA_signal_1275), .Q (new_AGEMA_signal_1276) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_1282) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C (clk), .D (new_AGEMA_signal_1287), .Q (new_AGEMA_signal_1288) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C (clk), .D (new_AGEMA_signal_1293), .Q (new_AGEMA_signal_1294) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C (clk), .D (new_AGEMA_signal_1299), .Q (new_AGEMA_signal_1300) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C (clk), .D (new_AGEMA_signal_1305), .Q (new_AGEMA_signal_1306) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C (clk), .D (new_AGEMA_signal_1311), .Q (new_AGEMA_signal_1312) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C (clk), .D (new_AGEMA_signal_1317), .Q (new_AGEMA_signal_1318) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C (clk), .D (new_AGEMA_signal_1323), .Q (new_AGEMA_signal_1324) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C (clk), .D (new_AGEMA_signal_1329), .Q (new_AGEMA_signal_1330) ) ;
    buf_clk new_AGEMA_reg_buffer_405 ( .C (clk), .D (new_AGEMA_signal_1335), .Q (new_AGEMA_signal_1336) ) ;
    buf_clk new_AGEMA_reg_buffer_411 ( .C (clk), .D (new_AGEMA_signal_1341), .Q (new_AGEMA_signal_1342) ) ;
    buf_clk new_AGEMA_reg_buffer_417 ( .C (clk), .D (new_AGEMA_signal_1347), .Q (new_AGEMA_signal_1348) ) ;
    buf_clk new_AGEMA_reg_buffer_423 ( .C (clk), .D (new_AGEMA_signal_1353), .Q (new_AGEMA_signal_1354) ) ;
    buf_clk new_AGEMA_reg_buffer_429 ( .C (clk), .D (new_AGEMA_signal_1359), .Q (new_AGEMA_signal_1360) ) ;
    buf_clk new_AGEMA_reg_buffer_435 ( .C (clk), .D (new_AGEMA_signal_1365), .Q (new_AGEMA_signal_1366) ) ;
    buf_clk new_AGEMA_reg_buffer_441 ( .C (clk), .D (new_AGEMA_signal_1371), .Q (new_AGEMA_signal_1372) ) ;
    buf_clk new_AGEMA_reg_buffer_447 ( .C (clk), .D (new_AGEMA_signal_1377), .Q (new_AGEMA_signal_1378) ) ;
    buf_clk new_AGEMA_reg_buffer_453 ( .C (clk), .D (new_AGEMA_signal_1383), .Q (new_AGEMA_signal_1384) ) ;
    buf_clk new_AGEMA_reg_buffer_459 ( .C (clk), .D (new_AGEMA_signal_1389), .Q (new_AGEMA_signal_1390) ) ;
    buf_clk new_AGEMA_reg_buffer_465 ( .C (clk), .D (new_AGEMA_signal_1395), .Q (new_AGEMA_signal_1396) ) ;
    buf_clk new_AGEMA_reg_buffer_471 ( .C (clk), .D (new_AGEMA_signal_1401), .Q (new_AGEMA_signal_1402) ) ;
    buf_clk new_AGEMA_reg_buffer_477 ( .C (clk), .D (new_AGEMA_signal_1407), .Q (new_AGEMA_signal_1408) ) ;
    buf_clk new_AGEMA_reg_buffer_483 ( .C (clk), .D (new_AGEMA_signal_1413), .Q (new_AGEMA_signal_1414) ) ;
    buf_clk new_AGEMA_reg_buffer_489 ( .C (clk), .D (new_AGEMA_signal_1419), .Q (new_AGEMA_signal_1420) ) ;
    buf_clk new_AGEMA_reg_buffer_495 ( .C (clk), .D (new_AGEMA_signal_1425), .Q (new_AGEMA_signal_1426) ) ;
    buf_clk new_AGEMA_reg_buffer_501 ( .C (clk), .D (new_AGEMA_signal_1431), .Q (new_AGEMA_signal_1432) ) ;
    buf_clk new_AGEMA_reg_buffer_507 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_1438) ) ;
    buf_clk new_AGEMA_reg_buffer_513 ( .C (clk), .D (new_AGEMA_signal_1443), .Q (new_AGEMA_signal_1444) ) ;
    buf_clk new_AGEMA_reg_buffer_519 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_1450) ) ;
    buf_clk new_AGEMA_reg_buffer_525 ( .C (clk), .D (new_AGEMA_signal_1455), .Q (new_AGEMA_signal_1456) ) ;
    buf_clk new_AGEMA_reg_buffer_531 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_1462) ) ;
    buf_clk new_AGEMA_reg_buffer_537 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_1468) ) ;
    buf_clk new_AGEMA_reg_buffer_543 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_1474) ) ;
    buf_clk new_AGEMA_reg_buffer_549 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_1480) ) ;
    buf_clk new_AGEMA_reg_buffer_555 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_1486) ) ;
    buf_clk new_AGEMA_reg_buffer_561 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_1492) ) ;
    buf_clk new_AGEMA_reg_buffer_567 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_1498) ) ;
    buf_clk new_AGEMA_reg_buffer_573 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_1504) ) ;
    buf_clk new_AGEMA_reg_buffer_579 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_1510) ) ;
    buf_clk new_AGEMA_reg_buffer_585 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_1516) ) ;
    buf_clk new_AGEMA_reg_buffer_591 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_1522) ) ;
    buf_clk new_AGEMA_reg_buffer_597 ( .C (clk), .D (new_AGEMA_signal_1527), .Q (new_AGEMA_signal_1528) ) ;
    buf_clk new_AGEMA_reg_buffer_603 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_1534) ) ;
    buf_clk new_AGEMA_reg_buffer_609 ( .C (clk), .D (new_AGEMA_signal_1539), .Q (new_AGEMA_signal_1540) ) ;
    buf_clk new_AGEMA_reg_buffer_615 ( .C (clk), .D (new_AGEMA_signal_1545), .Q (new_AGEMA_signal_1546) ) ;
    buf_clk new_AGEMA_reg_buffer_621 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_1552) ) ;
    buf_clk new_AGEMA_reg_buffer_627 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_1558) ) ;
    buf_clk new_AGEMA_reg_buffer_633 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_1564) ) ;
    buf_clk new_AGEMA_reg_buffer_639 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_1570) ) ;
    buf_clk new_AGEMA_reg_buffer_645 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_1576) ) ;
    buf_clk new_AGEMA_reg_buffer_651 ( .C (clk), .D (new_AGEMA_signal_1581), .Q (new_AGEMA_signal_1582) ) ;
    buf_clk new_AGEMA_reg_buffer_657 ( .C (clk), .D (new_AGEMA_signal_1587), .Q (new_AGEMA_signal_1588) ) ;
    buf_clk new_AGEMA_reg_buffer_663 ( .C (clk), .D (new_AGEMA_signal_1593), .Q (new_AGEMA_signal_1594) ) ;
    buf_clk new_AGEMA_reg_buffer_669 ( .C (clk), .D (new_AGEMA_signal_1599), .Q (new_AGEMA_signal_1600) ) ;
    buf_clk new_AGEMA_reg_buffer_675 ( .C (clk), .D (new_AGEMA_signal_1605), .Q (new_AGEMA_signal_1606) ) ;
    buf_clk new_AGEMA_reg_buffer_681 ( .C (clk), .D (new_AGEMA_signal_1611), .Q (new_AGEMA_signal_1612) ) ;
    buf_clk new_AGEMA_reg_buffer_687 ( .C (clk), .D (new_AGEMA_signal_1617), .Q (new_AGEMA_signal_1618) ) ;
    buf_clk new_AGEMA_reg_buffer_693 ( .C (clk), .D (new_AGEMA_signal_1623), .Q (new_AGEMA_signal_1624) ) ;
    buf_clk new_AGEMA_reg_buffer_699 ( .C (clk), .D (new_AGEMA_signal_1629), .Q (new_AGEMA_signal_1630) ) ;
    buf_clk new_AGEMA_reg_buffer_705 ( .C (clk), .D (new_AGEMA_signal_1635), .Q (new_AGEMA_signal_1636) ) ;
    buf_clk new_AGEMA_reg_buffer_711 ( .C (clk), .D (new_AGEMA_signal_1641), .Q (new_AGEMA_signal_1642) ) ;
    buf_clk new_AGEMA_reg_buffer_717 ( .C (clk), .D (new_AGEMA_signal_1647), .Q (new_AGEMA_signal_1648) ) ;
    buf_clk new_AGEMA_reg_buffer_723 ( .C (clk), .D (new_AGEMA_signal_1653), .Q (new_AGEMA_signal_1654) ) ;
    buf_clk new_AGEMA_reg_buffer_729 ( .C (clk), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_1660) ) ;
    buf_clk new_AGEMA_reg_buffer_735 ( .C (clk), .D (new_AGEMA_signal_1665), .Q (new_AGEMA_signal_1666) ) ;
    buf_clk new_AGEMA_reg_buffer_741 ( .C (clk), .D (new_AGEMA_signal_1671), .Q (new_AGEMA_signal_1672) ) ;
    buf_clk new_AGEMA_reg_buffer_747 ( .C (clk), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_1678) ) ;
    buf_clk new_AGEMA_reg_buffer_753 ( .C (clk), .D (new_AGEMA_signal_1683), .Q (new_AGEMA_signal_1684) ) ;
    buf_clk new_AGEMA_reg_buffer_759 ( .C (clk), .D (new_AGEMA_signal_1689), .Q (new_AGEMA_signal_1690) ) ;
    buf_clk new_AGEMA_reg_buffer_765 ( .C (clk), .D (new_AGEMA_signal_1695), .Q (new_AGEMA_signal_1696) ) ;
    buf_clk new_AGEMA_reg_buffer_771 ( .C (clk), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_1702) ) ;
    buf_clk new_AGEMA_reg_buffer_777 ( .C (clk), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_1708) ) ;
    buf_clk new_AGEMA_reg_buffer_783 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_1714) ) ;
    buf_clk new_AGEMA_reg_buffer_789 ( .C (clk), .D (new_AGEMA_signal_1719), .Q (new_AGEMA_signal_1720) ) ;
    buf_clk new_AGEMA_reg_buffer_795 ( .C (clk), .D (new_AGEMA_signal_1725), .Q (new_AGEMA_signal_1726) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M46_U1 ( .a ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}), .b ({new_AGEMA_signal_1216, new_AGEMA_signal_1210, new_AGEMA_signal_1204, new_AGEMA_signal_1198, new_AGEMA_signal_1192}), .clk (clk), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M47_U1 ( .a ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .b ({new_AGEMA_signal_1246, new_AGEMA_signal_1240, new_AGEMA_signal_1234, new_AGEMA_signal_1228, new_AGEMA_signal_1222}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, new_AGEMA_signal_467, M47}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M48_U1 ( .a ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1270, new_AGEMA_signal_1264, new_AGEMA_signal_1258, new_AGEMA_signal_1252}), .clk (clk), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M49_U1 ( .a ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}), .b ({new_AGEMA_signal_1306, new_AGEMA_signal_1300, new_AGEMA_signal_1294, new_AGEMA_signal_1288, new_AGEMA_signal_1282}), .clk (clk), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, M49}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M50_U1 ( .a ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .b ({new_AGEMA_signal_1336, new_AGEMA_signal_1330, new_AGEMA_signal_1324, new_AGEMA_signal_1318, new_AGEMA_signal_1312}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M51_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_1366, new_AGEMA_signal_1360, new_AGEMA_signal_1354, new_AGEMA_signal_1348, new_AGEMA_signal_1342}), .clk (clk), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M52_U1 ( .a ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .b ({new_AGEMA_signal_1396, new_AGEMA_signal_1390, new_AGEMA_signal_1384, new_AGEMA_signal_1378, new_AGEMA_signal_1372}), .clk (clk), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M53_U1 ( .a ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}), .b ({new_AGEMA_signal_1426, new_AGEMA_signal_1420, new_AGEMA_signal_1414, new_AGEMA_signal_1408, new_AGEMA_signal_1402}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M54_U1 ( .a ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .b ({new_AGEMA_signal_1456, new_AGEMA_signal_1450, new_AGEMA_signal_1444, new_AGEMA_signal_1438, new_AGEMA_signal_1432}), .clk (clk), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, new_AGEMA_signal_515, M54}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M55_U1 ( .a ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}), .b ({new_AGEMA_signal_1486, new_AGEMA_signal_1480, new_AGEMA_signal_1474, new_AGEMA_signal_1468, new_AGEMA_signal_1462}), .clk (clk), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M56_U1 ( .a ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .b ({new_AGEMA_signal_1516, new_AGEMA_signal_1510, new_AGEMA_signal_1504, new_AGEMA_signal_1498, new_AGEMA_signal_1492}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M57_U1 ( .a ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .b ({new_AGEMA_signal_1546, new_AGEMA_signal_1540, new_AGEMA_signal_1534, new_AGEMA_signal_1528, new_AGEMA_signal_1522}), .clk (clk), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, M57}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M58_U1 ( .a ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1570, new_AGEMA_signal_1564, new_AGEMA_signal_1558, new_AGEMA_signal_1552}), .clk (clk), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M59_U1 ( .a ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1600, new_AGEMA_signal_1594, new_AGEMA_signal_1588, new_AGEMA_signal_1582}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, new_AGEMA_signal_491, M59}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M60_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1630, new_AGEMA_signal_1624, new_AGEMA_signal_1618, new_AGEMA_signal_1612}), .clk (clk), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, M60}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M61_U1 ( .a ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1660, new_AGEMA_signal_1654, new_AGEMA_signal_1648, new_AGEMA_signal_1642}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M62_U1 ( .a ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}), .b ({new_AGEMA_signal_1696, new_AGEMA_signal_1690, new_AGEMA_signal_1684, new_AGEMA_signal_1678, new_AGEMA_signal_1672}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND_M63_U1 ( .a ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1720, new_AGEMA_signal_1714, new_AGEMA_signal_1708, new_AGEMA_signal_1702}), .clk (clk), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, M63}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L0_U1 ( .a ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .b ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}), .c ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L1_U1 ( .a ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}), .b ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}), .c ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L2_U1 ( .a ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}), .b ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}), .c ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L3_U1 ( .a ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, new_AGEMA_signal_467, M47}), .b ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}), .c ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L4_U1 ( .a ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, new_AGEMA_signal_515, M54}), .b ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}), .c ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L5_U1 ( .a ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, M49}), .b ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .c ({new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, L5}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L6_U1 ( .a ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}), .b ({new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, L5}), .c ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L7_U1 ( .a ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}), .b ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}), .c ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L8_U1 ( .a ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}), .b ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, new_AGEMA_signal_491, M59}), .c ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L9_U1 ( .a ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}), .b ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}), .c ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L10_U1 ( .a ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}), .b ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}), .c ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L11_U1 ( .a ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, M60}), .b ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}), .c ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L12_U1 ( .a ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}), .b ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}), .c ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, L12}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L13_U1 ( .a ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .c ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, new_AGEMA_signal_623, L13}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L14_U1 ( .a ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}), .b ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .c ({new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, new_AGEMA_signal_571, L14}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L15_U1 ( .a ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, new_AGEMA_signal_575, L15}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L16_U1 ( .a ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .c ({new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, L16}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L17_U1 ( .a ({new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, M57}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, L17}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L18_U1 ( .a ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}), .b ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}), .c ({new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, new_AGEMA_signal_583, L18}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L19_U1 ( .a ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, M63}), .b ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}), .c ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, new_AGEMA_signal_611, L19}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L20_U1 ( .a ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, new_AGEMA_signal_631, L20}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L21_U1 ( .a ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .b ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}), .c ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, new_AGEMA_signal_635, L21}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L22_U1 ( .a ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}), .b ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, L12}), .c ({new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, L22}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L23_U1 ( .a ({new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, new_AGEMA_signal_583, L18}), .b ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}), .c ({new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, new_AGEMA_signal_619, L23}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L24_U1 ( .a ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, new_AGEMA_signal_575, L15}), .b ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}), .c ({new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, L24}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L25_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}), .c ({new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, new_AGEMA_signal_643, L25}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L26_U1 ( .a ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}), .b ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}), .c ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, new_AGEMA_signal_647, L26}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L27_U1 ( .a ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}), .b ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}), .c ({new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, L27}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L28_U1 ( .a ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}), .b ({new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, new_AGEMA_signal_571, L14}), .c ({new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, new_AGEMA_signal_655, L28}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_L29_U1 ( .a ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}), .b ({new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, L17}), .c ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, new_AGEMA_signal_659, L29}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S0_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, L24}), .c ({new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, new_AGEMA_signal_667, O[7]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S1_U1 ( .a ({new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, L16}), .b ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, new_AGEMA_signal_647, L26}), .c ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, new_AGEMA_signal_671, O[6]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S2_U1 ( .a ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, new_AGEMA_signal_611, L19}), .b ({new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, new_AGEMA_signal_655, L28}), .c ({new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, O[5]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S3_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, new_AGEMA_signal_635, L21}), .c ({new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, new_AGEMA_signal_679, O[4]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S4_U1 ( .a ({new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, new_AGEMA_signal_631, L20}), .b ({new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, L22}), .c ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, new_AGEMA_signal_683, O[3]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S5_U1 ( .a ({new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, new_AGEMA_signal_643, L25}), .b ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, new_AGEMA_signal_659, L29}), .c ({new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, O[2]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S6_U1 ( .a ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, new_AGEMA_signal_623, L13}), .b ({new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, L27}), .c ({new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, new_AGEMA_signal_691, O[1]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR_S7_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, new_AGEMA_signal_619, L23}), .c ({new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, O[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_7_ ( .clk (clk), .D ({new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, new_AGEMA_signal_667, O[7]}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_6_ ( .clk (clk), .D ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, new_AGEMA_signal_671, O[6]}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_5_ ( .clk (clk), .D ({new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, O[5]}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_4_ ( .clk (clk), .D ({new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, new_AGEMA_signal_679, O[4]}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, new_AGEMA_signal_683, O[3]}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, O[2]}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, new_AGEMA_signal_691, O[1]}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, O[0]}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
