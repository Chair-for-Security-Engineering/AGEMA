/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDsylvan_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [4283:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;

    /* cells in depth 0 */
    MUX2_X1 cell_176 ( .S ( 1'b1 ), .A ( 1'b1 ), .B ( 1'b0 ), .Z ( signal_192 ) ) ;
    MUX2_X1 cell_177 ( .S ( 1'b1 ), .A ( 1'b0 ), .B ( 1'b1 ), .Z ( signal_193 ) ) ;

    /* cells in depth 1 */
    buf_clk cell_892 ( .C ( clk ), .D ( X_s0[1] ), .Q ( signal_7374 ) ) ;
    buf_clk cell_894 ( .C ( clk ), .D ( X_s1[1] ), .Q ( signal_7376 ) ) ;
    buf_clk cell_896 ( .C ( clk ), .D ( X_s2[1] ), .Q ( signal_7378 ) ) ;
    buf_clk cell_898 ( .C ( clk ), .D ( X_s3[1] ), .Q ( signal_7380 ) ) ;
    buf_clk cell_900 ( .C ( clk ), .D ( signal_193 ), .Q ( signal_7382 ) ) ;
    buf_clk cell_902 ( .C ( clk ), .D ( signal_192 ), .Q ( signal_7384 ) ) ;
    buf_clk cell_904 ( .C ( clk ), .D ( X_s0[2] ), .Q ( signal_7386 ) ) ;
    buf_clk cell_906 ( .C ( clk ), .D ( X_s1[2] ), .Q ( signal_7388 ) ) ;
    buf_clk cell_908 ( .C ( clk ), .D ( X_s2[2] ), .Q ( signal_7390 ) ) ;
    buf_clk cell_910 ( .C ( clk ), .D ( X_s3[2] ), .Q ( signal_7392 ) ) ;
    buf_clk cell_1084 ( .C ( clk ), .D ( X_s0[3] ), .Q ( signal_7566 ) ) ;
    buf_clk cell_1090 ( .C ( clk ), .D ( X_s1[3] ), .Q ( signal_7572 ) ) ;
    buf_clk cell_1096 ( .C ( clk ), .D ( X_s2[3] ), .Q ( signal_7578 ) ) ;
    buf_clk cell_1102 ( .C ( clk ), .D ( X_s3[3] ), .Q ( signal_7584 ) ) ;
    buf_clk cell_1124 ( .C ( clk ), .D ( X_s0[4] ), .Q ( signal_7606 ) ) ;
    buf_clk cell_1132 ( .C ( clk ), .D ( X_s1[4] ), .Q ( signal_7614 ) ) ;
    buf_clk cell_1140 ( .C ( clk ), .D ( X_s2[4] ), .Q ( signal_7622 ) ) ;
    buf_clk cell_1148 ( .C ( clk ), .D ( X_s3[4] ), .Q ( signal_7630 ) ) ;
    buf_clk cell_1156 ( .C ( clk ), .D ( X_s0[5] ), .Q ( signal_7638 ) ) ;
    buf_clk cell_1166 ( .C ( clk ), .D ( X_s1[5] ), .Q ( signal_7648 ) ) ;
    buf_clk cell_1176 ( .C ( clk ), .D ( X_s2[5] ), .Q ( signal_7658 ) ) ;
    buf_clk cell_1186 ( .C ( clk ), .D ( X_s3[5] ), .Q ( signal_7668 ) ) ;
    buf_clk cell_1196 ( .C ( clk ), .D ( X_s0[6] ), .Q ( signal_7678 ) ) ;
    buf_clk cell_1208 ( .C ( clk ), .D ( X_s1[6] ), .Q ( signal_7690 ) ) ;
    buf_clk cell_1220 ( .C ( clk ), .D ( X_s2[6] ), .Q ( signal_7702 ) ) ;
    buf_clk cell_1232 ( .C ( clk ), .D ( X_s3[6] ), .Q ( signal_7714 ) ) ;
    buf_clk cell_1244 ( .C ( clk ), .D ( X_s0[7] ), .Q ( signal_7726 ) ) ;
    buf_clk cell_1258 ( .C ( clk ), .D ( X_s1[7] ), .Q ( signal_7740 ) ) ;
    buf_clk cell_1272 ( .C ( clk ), .D ( X_s2[7] ), .Q ( signal_7754 ) ) ;
    buf_clk cell_1286 ( .C ( clk ), .D ( X_s3[7] ), .Q ( signal_7768 ) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_178 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_905, signal_904, signal_903, signal_194}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_179 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_908, signal_907, signal_906, signal_195}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_180 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_914, signal_913, signal_912, signal_196}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_181 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_917, signal_916, signal_915, signal_197}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_182 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_920, signal_919, signal_918, signal_198}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_183 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_923, signal_922, signal_921, signal_199}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_184 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_926, signal_925, signal_924, signal_200}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_185 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, signal_193}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_929, signal_928, signal_927, signal_201}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_186 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_932, signal_931, signal_930, signal_202}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_187 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_935, signal_934, signal_933, signal_203}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_188 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_938, signal_937, signal_936, signal_204}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_189 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_941, signal_940, signal_939, signal_205}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_190 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, signal_193}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_944, signal_943, signal_942, signal_206}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_192 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, signal_193}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_950, signal_949, signal_948, signal_208}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_193 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_953, signal_952, signal_951, signal_209}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_194 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_956, signal_955, signal_954, signal_210}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_195 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, signal_193}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_959, signal_958, signal_957, signal_211}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_198 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_968, signal_967, signal_966, signal_214}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_202 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, signal_193}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_980, signal_979, signal_978, signal_218}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_203 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_983, signal_982, signal_981, signal_219}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_207 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_995, signal_994, signal_993, signal_223}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_209 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_193}), .a ({1'b0, 1'b0, 1'b0, signal_192}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_1001, signal_1000, signal_999, signal_225}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_215 ( .s ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0, signal_192}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_1019, signal_1018, signal_1017, signal_231}) ) ;
    buf_clk cell_893 ( .C ( clk ), .D ( signal_7374 ), .Q ( signal_7375 ) ) ;
    buf_clk cell_895 ( .C ( clk ), .D ( signal_7376 ), .Q ( signal_7377 ) ) ;
    buf_clk cell_897 ( .C ( clk ), .D ( signal_7378 ), .Q ( signal_7379 ) ) ;
    buf_clk cell_899 ( .C ( clk ), .D ( signal_7380 ), .Q ( signal_7381 ) ) ;
    buf_clk cell_901 ( .C ( clk ), .D ( signal_7382 ), .Q ( signal_7383 ) ) ;
    buf_clk cell_903 ( .C ( clk ), .D ( signal_7384 ), .Q ( signal_7385 ) ) ;
    buf_clk cell_905 ( .C ( clk ), .D ( signal_7386 ), .Q ( signal_7387 ) ) ;
    buf_clk cell_907 ( .C ( clk ), .D ( signal_7388 ), .Q ( signal_7389 ) ) ;
    buf_clk cell_909 ( .C ( clk ), .D ( signal_7390 ), .Q ( signal_7391 ) ) ;
    buf_clk cell_911 ( .C ( clk ), .D ( signal_7392 ), .Q ( signal_7393 ) ) ;
    buf_clk cell_1085 ( .C ( clk ), .D ( signal_7566 ), .Q ( signal_7567 ) ) ;
    buf_clk cell_1091 ( .C ( clk ), .D ( signal_7572 ), .Q ( signal_7573 ) ) ;
    buf_clk cell_1097 ( .C ( clk ), .D ( signal_7578 ), .Q ( signal_7579 ) ) ;
    buf_clk cell_1103 ( .C ( clk ), .D ( signal_7584 ), .Q ( signal_7585 ) ) ;
    buf_clk cell_1125 ( .C ( clk ), .D ( signal_7606 ), .Q ( signal_7607 ) ) ;
    buf_clk cell_1133 ( .C ( clk ), .D ( signal_7614 ), .Q ( signal_7615 ) ) ;
    buf_clk cell_1141 ( .C ( clk ), .D ( signal_7622 ), .Q ( signal_7623 ) ) ;
    buf_clk cell_1149 ( .C ( clk ), .D ( signal_7630 ), .Q ( signal_7631 ) ) ;
    buf_clk cell_1157 ( .C ( clk ), .D ( signal_7638 ), .Q ( signal_7639 ) ) ;
    buf_clk cell_1167 ( .C ( clk ), .D ( signal_7648 ), .Q ( signal_7649 ) ) ;
    buf_clk cell_1177 ( .C ( clk ), .D ( signal_7658 ), .Q ( signal_7659 ) ) ;
    buf_clk cell_1187 ( .C ( clk ), .D ( signal_7668 ), .Q ( signal_7669 ) ) ;
    buf_clk cell_1197 ( .C ( clk ), .D ( signal_7678 ), .Q ( signal_7679 ) ) ;
    buf_clk cell_1209 ( .C ( clk ), .D ( signal_7690 ), .Q ( signal_7691 ) ) ;
    buf_clk cell_1221 ( .C ( clk ), .D ( signal_7702 ), .Q ( signal_7703 ) ) ;
    buf_clk cell_1233 ( .C ( clk ), .D ( signal_7714 ), .Q ( signal_7715 ) ) ;
    buf_clk cell_1245 ( .C ( clk ), .D ( signal_7726 ), .Q ( signal_7727 ) ) ;
    buf_clk cell_1259 ( .C ( clk ), .D ( signal_7740 ), .Q ( signal_7741 ) ) ;
    buf_clk cell_1273 ( .C ( clk ), .D ( signal_7754 ), .Q ( signal_7755 ) ) ;
    buf_clk cell_1287 ( .C ( clk ), .D ( signal_7768 ), .Q ( signal_7769 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_912 ( .C ( clk ), .D ( signal_7387 ), .Q ( signal_7394 ) ) ;
    buf_clk cell_914 ( .C ( clk ), .D ( signal_7389 ), .Q ( signal_7396 ) ) ;
    buf_clk cell_916 ( .C ( clk ), .D ( signal_7391 ), .Q ( signal_7398 ) ) ;
    buf_clk cell_918 ( .C ( clk ), .D ( signal_7393 ), .Q ( signal_7400 ) ) ;
    buf_clk cell_920 ( .C ( clk ), .D ( signal_211 ), .Q ( signal_7402 ) ) ;
    buf_clk cell_922 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_7404 ) ) ;
    buf_clk cell_924 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_7406 ) ) ;
    buf_clk cell_926 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_7408 ) ) ;
    buf_clk cell_928 ( .C ( clk ), .D ( signal_196 ), .Q ( signal_7410 ) ) ;
    buf_clk cell_930 ( .C ( clk ), .D ( signal_912 ), .Q ( signal_7412 ) ) ;
    buf_clk cell_932 ( .C ( clk ), .D ( signal_913 ), .Q ( signal_7414 ) ) ;
    buf_clk cell_934 ( .C ( clk ), .D ( signal_914 ), .Q ( signal_7416 ) ) ;
    buf_clk cell_936 ( .C ( clk ), .D ( signal_214 ), .Q ( signal_7418 ) ) ;
    buf_clk cell_938 ( .C ( clk ), .D ( signal_966 ), .Q ( signal_7420 ) ) ;
    buf_clk cell_940 ( .C ( clk ), .D ( signal_967 ), .Q ( signal_7422 ) ) ;
    buf_clk cell_942 ( .C ( clk ), .D ( signal_968 ), .Q ( signal_7424 ) ) ;
    buf_clk cell_944 ( .C ( clk ), .D ( signal_218 ), .Q ( signal_7426 ) ) ;
    buf_clk cell_946 ( .C ( clk ), .D ( signal_978 ), .Q ( signal_7428 ) ) ;
    buf_clk cell_948 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_7430 ) ) ;
    buf_clk cell_950 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_7432 ) ) ;
    buf_clk cell_952 ( .C ( clk ), .D ( signal_200 ), .Q ( signal_7434 ) ) ;
    buf_clk cell_954 ( .C ( clk ), .D ( signal_924 ), .Q ( signal_7436 ) ) ;
    buf_clk cell_956 ( .C ( clk ), .D ( signal_925 ), .Q ( signal_7438 ) ) ;
    buf_clk cell_958 ( .C ( clk ), .D ( signal_926 ), .Q ( signal_7440 ) ) ;
    buf_clk cell_960 ( .C ( clk ), .D ( signal_7385 ), .Q ( signal_7442 ) ) ;
    buf_clk cell_962 ( .C ( clk ), .D ( signal_206 ), .Q ( signal_7444 ) ) ;
    buf_clk cell_964 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_7446 ) ) ;
    buf_clk cell_966 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_7448 ) ) ;
    buf_clk cell_968 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_7450 ) ) ;
    buf_clk cell_970 ( .C ( clk ), .D ( signal_194 ), .Q ( signal_7452 ) ) ;
    buf_clk cell_972 ( .C ( clk ), .D ( signal_903 ), .Q ( signal_7454 ) ) ;
    buf_clk cell_974 ( .C ( clk ), .D ( signal_904 ), .Q ( signal_7456 ) ) ;
    buf_clk cell_976 ( .C ( clk ), .D ( signal_905 ), .Q ( signal_7458 ) ) ;
    buf_clk cell_978 ( .C ( clk ), .D ( signal_208 ), .Q ( signal_7460 ) ) ;
    buf_clk cell_980 ( .C ( clk ), .D ( signal_948 ), .Q ( signal_7462 ) ) ;
    buf_clk cell_982 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_7464 ) ) ;
    buf_clk cell_984 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_7466 ) ) ;
    buf_clk cell_986 ( .C ( clk ), .D ( signal_209 ), .Q ( signal_7468 ) ) ;
    buf_clk cell_988 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_7470 ) ) ;
    buf_clk cell_990 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_7472 ) ) ;
    buf_clk cell_992 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_7474 ) ) ;
    buf_clk cell_994 ( .C ( clk ), .D ( signal_210 ), .Q ( signal_7476 ) ) ;
    buf_clk cell_996 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_7478 ) ) ;
    buf_clk cell_998 ( .C ( clk ), .D ( signal_955 ), .Q ( signal_7480 ) ) ;
    buf_clk cell_1000 ( .C ( clk ), .D ( signal_956 ), .Q ( signal_7482 ) ) ;
    buf_clk cell_1002 ( .C ( clk ), .D ( signal_7383 ), .Q ( signal_7484 ) ) ;
    buf_clk cell_1004 ( .C ( clk ), .D ( signal_205 ), .Q ( signal_7486 ) ) ;
    buf_clk cell_1006 ( .C ( clk ), .D ( signal_939 ), .Q ( signal_7488 ) ) ;
    buf_clk cell_1008 ( .C ( clk ), .D ( signal_940 ), .Q ( signal_7490 ) ) ;
    buf_clk cell_1010 ( .C ( clk ), .D ( signal_941 ), .Q ( signal_7492 ) ) ;
    buf_clk cell_1012 ( .C ( clk ), .D ( signal_198 ), .Q ( signal_7494 ) ) ;
    buf_clk cell_1014 ( .C ( clk ), .D ( signal_918 ), .Q ( signal_7496 ) ) ;
    buf_clk cell_1016 ( .C ( clk ), .D ( signal_919 ), .Q ( signal_7498 ) ) ;
    buf_clk cell_1018 ( .C ( clk ), .D ( signal_920 ), .Q ( signal_7500 ) ) ;
    buf_clk cell_1020 ( .C ( clk ), .D ( signal_219 ), .Q ( signal_7502 ) ) ;
    buf_clk cell_1022 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_7504 ) ) ;
    buf_clk cell_1024 ( .C ( clk ), .D ( signal_982 ), .Q ( signal_7506 ) ) ;
    buf_clk cell_1026 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_7508 ) ) ;
    buf_clk cell_1028 ( .C ( clk ), .D ( signal_197 ), .Q ( signal_7510 ) ) ;
    buf_clk cell_1030 ( .C ( clk ), .D ( signal_915 ), .Q ( signal_7512 ) ) ;
    buf_clk cell_1032 ( .C ( clk ), .D ( signal_916 ), .Q ( signal_7514 ) ) ;
    buf_clk cell_1034 ( .C ( clk ), .D ( signal_917 ), .Q ( signal_7516 ) ) ;
    buf_clk cell_1036 ( .C ( clk ), .D ( signal_204 ), .Q ( signal_7518 ) ) ;
    buf_clk cell_1038 ( .C ( clk ), .D ( signal_936 ), .Q ( signal_7520 ) ) ;
    buf_clk cell_1040 ( .C ( clk ), .D ( signal_937 ), .Q ( signal_7522 ) ) ;
    buf_clk cell_1042 ( .C ( clk ), .D ( signal_938 ), .Q ( signal_7524 ) ) ;
    buf_clk cell_1044 ( .C ( clk ), .D ( signal_223 ), .Q ( signal_7526 ) ) ;
    buf_clk cell_1046 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_7528 ) ) ;
    buf_clk cell_1048 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_7530 ) ) ;
    buf_clk cell_1050 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_7532 ) ) ;
    buf_clk cell_1052 ( .C ( clk ), .D ( signal_225 ), .Q ( signal_7534 ) ) ;
    buf_clk cell_1054 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_7536 ) ) ;
    buf_clk cell_1056 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_7538 ) ) ;
    buf_clk cell_1058 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_7540 ) ) ;
    buf_clk cell_1060 ( .C ( clk ), .D ( signal_201 ), .Q ( signal_7542 ) ) ;
    buf_clk cell_1062 ( .C ( clk ), .D ( signal_927 ), .Q ( signal_7544 ) ) ;
    buf_clk cell_1064 ( .C ( clk ), .D ( signal_928 ), .Q ( signal_7546 ) ) ;
    buf_clk cell_1066 ( .C ( clk ), .D ( signal_929 ), .Q ( signal_7548 ) ) ;
    buf_clk cell_1068 ( .C ( clk ), .D ( signal_231 ), .Q ( signal_7550 ) ) ;
    buf_clk cell_1070 ( .C ( clk ), .D ( signal_1017 ), .Q ( signal_7552 ) ) ;
    buf_clk cell_1072 ( .C ( clk ), .D ( signal_1018 ), .Q ( signal_7554 ) ) ;
    buf_clk cell_1074 ( .C ( clk ), .D ( signal_1019 ), .Q ( signal_7556 ) ) ;
    buf_clk cell_1076 ( .C ( clk ), .D ( signal_203 ), .Q ( signal_7558 ) ) ;
    buf_clk cell_1078 ( .C ( clk ), .D ( signal_933 ), .Q ( signal_7560 ) ) ;
    buf_clk cell_1080 ( .C ( clk ), .D ( signal_934 ), .Q ( signal_7562 ) ) ;
    buf_clk cell_1082 ( .C ( clk ), .D ( signal_935 ), .Q ( signal_7564 ) ) ;
    buf_clk cell_1086 ( .C ( clk ), .D ( signal_7567 ), .Q ( signal_7568 ) ) ;
    buf_clk cell_1092 ( .C ( clk ), .D ( signal_7573 ), .Q ( signal_7574 ) ) ;
    buf_clk cell_1098 ( .C ( clk ), .D ( signal_7579 ), .Q ( signal_7580 ) ) ;
    buf_clk cell_1104 ( .C ( clk ), .D ( signal_7585 ), .Q ( signal_7586 ) ) ;
    buf_clk cell_1126 ( .C ( clk ), .D ( signal_7607 ), .Q ( signal_7608 ) ) ;
    buf_clk cell_1134 ( .C ( clk ), .D ( signal_7615 ), .Q ( signal_7616 ) ) ;
    buf_clk cell_1142 ( .C ( clk ), .D ( signal_7623 ), .Q ( signal_7624 ) ) ;
    buf_clk cell_1150 ( .C ( clk ), .D ( signal_7631 ), .Q ( signal_7632 ) ) ;
    buf_clk cell_1158 ( .C ( clk ), .D ( signal_7639 ), .Q ( signal_7640 ) ) ;
    buf_clk cell_1168 ( .C ( clk ), .D ( signal_7649 ), .Q ( signal_7650 ) ) ;
    buf_clk cell_1178 ( .C ( clk ), .D ( signal_7659 ), .Q ( signal_7660 ) ) ;
    buf_clk cell_1188 ( .C ( clk ), .D ( signal_7669 ), .Q ( signal_7670 ) ) ;
    buf_clk cell_1198 ( .C ( clk ), .D ( signal_7679 ), .Q ( signal_7680 ) ) ;
    buf_clk cell_1210 ( .C ( clk ), .D ( signal_7691 ), .Q ( signal_7692 ) ) ;
    buf_clk cell_1222 ( .C ( clk ), .D ( signal_7703 ), .Q ( signal_7704 ) ) ;
    buf_clk cell_1234 ( .C ( clk ), .D ( signal_7715 ), .Q ( signal_7716 ) ) ;
    buf_clk cell_1246 ( .C ( clk ), .D ( signal_7727 ), .Q ( signal_7728 ) ) ;
    buf_clk cell_1260 ( .C ( clk ), .D ( signal_7741 ), .Q ( signal_7742 ) ) ;
    buf_clk cell_1274 ( .C ( clk ), .D ( signal_7755 ), .Q ( signal_7756 ) ) ;
    buf_clk cell_1288 ( .C ( clk ), .D ( signal_7769 ), .Q ( signal_7770 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_191 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_947, signal_946, signal_945, signal_207}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_196 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_962, signal_961, signal_960, signal_212}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_197 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_965, signal_964, signal_963, signal_213}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_199 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_971, signal_970, signal_969, signal_215}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_200 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_974, signal_973, signal_972, signal_216}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_201 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_977, signal_976, signal_975, signal_217}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_204 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_986, signal_985, signal_984, signal_220}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_205 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_989, signal_988, signal_987, signal_221}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_206 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_992, signal_991, signal_990, signal_222}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_208 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_998, signal_997, signal_996, signal_224}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_210 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_1004, signal_1003, signal_1002, signal_226}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_211 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_1007, signal_1006, signal_1005, signal_227}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_212 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_1010, signal_1009, signal_1008, signal_228}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_213 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_1013, signal_1012, signal_1011, signal_229}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_214 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_1016, signal_1015, signal_1014, signal_230}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_216 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_1022, signal_1021, signal_1020, signal_232}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_217 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_1025, signal_1024, signal_1023, signal_233}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_218 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_1028, signal_1027, signal_1026, signal_234}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_219 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_1031, signal_1030, signal_1029, signal_235}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_220 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_1034, signal_1033, signal_1032, signal_236}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_221 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_1037, signal_1036, signal_1035, signal_237}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_222 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_1040, signal_1039, signal_1038, signal_238}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_223 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_1043, signal_1042, signal_1041, signal_239}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_224 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_1046, signal_1045, signal_1044, signal_240}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_225 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_1049, signal_1048, signal_1047, signal_241}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_226 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_1052, signal_1051, signal_1050, signal_242}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_227 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_1055, signal_1054, signal_1053, signal_243}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_228 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_1058, signal_1057, signal_1056, signal_244}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_229 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_1061, signal_1060, signal_1059, signal_245}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_230 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_1064, signal_1063, signal_1062, signal_246}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_231 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_1067, signal_1066, signal_1065, signal_247}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_232 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_1070, signal_1069, signal_1068, signal_248}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_233 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_1073, signal_1072, signal_1071, signal_249}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_234 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_1076, signal_1075, signal_1074, signal_250}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_235 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_1079, signal_1078, signal_1077, signal_251}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_236 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_1082, signal_1081, signal_1080, signal_252}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_237 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_1085, signal_1084, signal_1083, signal_253}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_238 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_1088, signal_1087, signal_1086, signal_254}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_239 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_1091, signal_1090, signal_1089, signal_255}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_240 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_1094, signal_1093, signal_1092, signal_256}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_241 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_1097, signal_1096, signal_1095, signal_257}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_242 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_1100, signal_1099, signal_1098, signal_258}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_243 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_1103, signal_1102, signal_1101, signal_259}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_244 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_1106, signal_1105, signal_1104, signal_260}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_245 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_1109, signal_1108, signal_1107, signal_261}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_246 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_1112, signal_1111, signal_1110, signal_262}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_247 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_1115, signal_1114, signal_1113, signal_263}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_248 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_1118, signal_1117, signal_1116, signal_264}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_249 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_1121, signal_1120, signal_1119, signal_265}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_250 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_1124, signal_1123, signal_1122, signal_266}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_251 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_1127, signal_1126, signal_1125, signal_267}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_252 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_1130, signal_1129, signal_1128, signal_268}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_253 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_1133, signal_1132, signal_1131, signal_269}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_254 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_1136, signal_1135, signal_1134, signal_270}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_255 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_1139, signal_1138, signal_1137, signal_271}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_256 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_1142, signal_1141, signal_1140, signal_272}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_257 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_1145, signal_1144, signal_1143, signal_273}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_258 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_1148, signal_1147, signal_1146, signal_274}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_259 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_1151, signal_1150, signal_1149, signal_275}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_260 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_1154, signal_1153, signal_1152, signal_276}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_261 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_1157, signal_1156, signal_1155, signal_277}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_262 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_1160, signal_1159, signal_1158, signal_278}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_263 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_1163, signal_1162, signal_1161, signal_279}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_265 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_1172, signal_1171, signal_1170, signal_281}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_266 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_1175, signal_1174, signal_1173, signal_282}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_267 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_1178, signal_1177, signal_1176, signal_283}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_268 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_1181, signal_1180, signal_1179, signal_284}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_269 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_1184, signal_1183, signal_1182, signal_285}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_270 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_1187, signal_1186, signal_1185, signal_286}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_271 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_1190, signal_1189, signal_1188, signal_287}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_272 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_1193, signal_1192, signal_1191, signal_288}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_273 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_1196, signal_1195, signal_1194, signal_289}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_274 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_1199, signal_1198, signal_1197, signal_290}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_275 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_1202, signal_1201, signal_1200, signal_291}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_276 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_1205, signal_1204, signal_1203, signal_292}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_277 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_1208, signal_1207, signal_1206, signal_293}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_278 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_1211, signal_1210, signal_1209, signal_294}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_279 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_1214, signal_1213, signal_1212, signal_295}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_280 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_1217, signal_1216, signal_1215, signal_296}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_281 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_1220, signal_1219, signal_1218, signal_297}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_282 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_1223, signal_1222, signal_1221, signal_298}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_283 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_1226, signal_1225, signal_1224, signal_299}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_284 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_1229, signal_1228, signal_1227, signal_300}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_285 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_1232, signal_1231, signal_1230, signal_301}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_286 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_1235, signal_1234, signal_1233, signal_302}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_287 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_1238, signal_1237, signal_1236, signal_303}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_288 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_1241, signal_1240, signal_1239, signal_304}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_289 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1244, signal_1243, signal_1242, signal_305}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_290 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_1247, signal_1246, signal_1245, signal_306}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_291 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_1250, signal_1249, signal_1248, signal_307}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_292 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_1253, signal_1252, signal_1251, signal_308}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_293 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_1256, signal_1255, signal_1254, signal_309}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_294 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1259, signal_1258, signal_1257, signal_310}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_295 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_1262, signal_1261, signal_1260, signal_311}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_296 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_1265, signal_1264, signal_1263, signal_312}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_297 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_1268, signal_1267, signal_1266, signal_313}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_298 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_1271, signal_1270, signal_1269, signal_314}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_299 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1274, signal_1273, signal_1272, signal_315}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_300 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_1277, signal_1276, signal_1275, signal_316}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_301 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_1280, signal_1279, signal_1278, signal_317}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_302 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_1283, signal_1282, signal_1281, signal_318}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_303 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_1286, signal_1285, signal_1284, signal_319}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_304 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1289, signal_1288, signal_1287, signal_320}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_305 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_1292, signal_1291, signal_1290, signal_321}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_306 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_1295, signal_1294, signal_1293, signal_322}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_307 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_1298, signal_1297, signal_1296, signal_323}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_308 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_1301, signal_1300, signal_1299, signal_324}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_309 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1304, signal_1303, signal_1302, signal_325}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_310 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_1307, signal_1306, signal_1305, signal_326}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_311 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_1310, signal_1309, signal_1308, signal_327}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_312 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_1313, signal_1312, signal_1311, signal_328}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_313 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_1316, signal_1315, signal_1314, signal_329}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_314 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1319, signal_1318, signal_1317, signal_330}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_315 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_1322, signal_1321, signal_1320, signal_331}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_316 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_1325, signal_1324, signal_1323, signal_332}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_317 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_1328, signal_1327, signal_1326, signal_333}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_318 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_1331, signal_1330, signal_1329, signal_334}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_319 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1334, signal_1333, signal_1332, signal_335}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_320 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_1337, signal_1336, signal_1335, signal_336}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_321 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_1340, signal_1339, signal_1338, signal_337}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_323 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_1346, signal_1345, signal_1344, signal_339}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_324 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_1349, signal_1348, signal_1347, signal_340}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_326 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1355, signal_1354, signal_1353, signal_342}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_327 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_1358, signal_1357, signal_1356, signal_343}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_328 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_1361, signal_1360, signal_1359, signal_344}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_330 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_1367, signal_1366, signal_1365, signal_346}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_331 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_1370, signal_1369, signal_1368, signal_347}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_332 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1373, signal_1372, signal_1371, signal_348}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_333 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_1376, signal_1375, signal_1374, signal_349}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_334 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_1379, signal_1378, signal_1377, signal_350}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_335 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_1382, signal_1381, signal_1380, signal_351}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_336 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_1385, signal_1384, signal_1383, signal_352}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_337 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_929, signal_928, signal_927, signal_201}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1388, signal_1387, signal_1386, signal_353}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_338 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_1391, signal_1390, signal_1389, signal_354}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_339 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_1394, signal_1393, signal_1392, signal_355}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_340 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_1397, signal_1396, signal_1395, signal_356}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_341 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_1400, signal_1399, signal_1398, signal_357}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_342 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1403, signal_1402, signal_1401, signal_358}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_343 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_1406, signal_1405, signal_1404, signal_359}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_344 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_1409, signal_1408, signal_1407, signal_360}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_345 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_1412, signal_1411, signal_1410, signal_361}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_346 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_1415, signal_1414, signal_1413, signal_362}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_347 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_1418, signal_1417, signal_1416, signal_363}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_348 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_932, signal_931, signal_930, signal_202}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_1421, signal_1420, signal_1419, signal_364}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_349 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_1424, signal_1423, signal_1422, signal_365}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_350 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_1427, signal_1426, signal_1425, signal_366}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_351 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_950, signal_949, signal_948, signal_208}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_1430, signal_1429, signal_1428, signal_367}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_352 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_1433, signal_1432, signal_1431, signal_368}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_353 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_1436, signal_1435, signal_1434, signal_369}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_354 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_1439, signal_1438, signal_1437, signal_370}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_355 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_1442, signal_1441, signal_1440, signal_371}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_356 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_1445, signal_1444, signal_1443, signal_372}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_357 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_926, signal_925, signal_924, signal_200}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_1448, signal_1447, signal_1446, signal_373}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_358 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_1451, signal_1450, signal_1449, signal_374}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_359 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_1454, signal_1453, signal_1452, signal_375}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_360 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_1457, signal_1456, signal_1455, signal_376}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_361 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_1460, signal_1459, signal_1458, signal_377}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_362 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1463, signal_1462, signal_1461, signal_378}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_363 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_1466, signal_1465, signal_1464, signal_379}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_364 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_1469, signal_1468, signal_1467, signal_380}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_365 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_1472, signal_1471, signal_1470, signal_381}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_366 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_938, signal_937, signal_936, signal_204}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_1475, signal_1474, signal_1473, signal_382}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_367 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_923, signal_922, signal_921, signal_199}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1478, signal_1477, signal_1476, signal_383}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_368 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_1481, signal_1480, signal_1479, signal_384}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_369 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_944, signal_943, signal_942, signal_206}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_1484, signal_1483, signal_1482, signal_385}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_370 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_920, signal_919, signal_918, signal_198}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_1487, signal_1486, signal_1485, signal_386}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_371 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_1490, signal_1489, signal_1488, signal_387}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_372 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1493, signal_1492, signal_1491, signal_388}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_373 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_1496, signal_1495, signal_1494, signal_389}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_374 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_1499, signal_1498, signal_1497, signal_390}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_375 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_1502, signal_1501, signal_1500, signal_391}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_376 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_1505, signal_1504, signal_1503, signal_392}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_377 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1508, signal_1507, signal_1506, signal_393}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_378 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_1511, signal_1510, signal_1509, signal_394}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_379 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_1514, signal_1513, signal_1512, signal_395}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_380 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_926, signal_925, signal_924, signal_200}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_1517, signal_1516, signal_1515, signal_396}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_381 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_1520, signal_1519, signal_1518, signal_397}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_382 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_935, signal_934, signal_933, signal_203}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1523, signal_1522, signal_1521, signal_398}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_383 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_923, signal_922, signal_921, signal_199}), .a ({signal_950, signal_949, signal_948, signal_208}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_1526, signal_1525, signal_1524, signal_399}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_384 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({1'b0, 1'b0, 1'b0, signal_7385}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_1529, signal_1528, signal_1527, signal_400}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_385 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_941, signal_940, signal_939, signal_205}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_1532, signal_1531, signal_1530, signal_401}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_386 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_905, signal_904, signal_903, signal_194}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_1535, signal_1534, signal_1533, signal_402}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_387 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_908, signal_907, signal_906, signal_195}), .a ({signal_944, signal_943, signal_942, signal_206}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_1538, signal_1537, signal_1536, signal_403}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_388 ( .s ({signal_7393, signal_7391, signal_7389, signal_7387}), .b ({signal_980, signal_979, signal_978, signal_218}), .a ({signal_983, signal_982, signal_981, signal_219}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({signal_1541, signal_1540, signal_1539, signal_404}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_389 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_941, signal_940, signal_939, signal_205}), .a ({1'b0, 1'b0, 1'b0, signal_7383}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({signal_1544, signal_1543, signal_1542, signal_405}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_390 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7383}), .a ({signal_935, signal_934, signal_933, signal_203}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({signal_1547, signal_1546, signal_1545, signal_406}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_391 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_938, signal_937, signal_936, signal_204}), .a ({signal_905, signal_904, signal_903, signal_194}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({signal_1550, signal_1549, signal_1548, signal_407}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_392 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_920, signal_919, signal_918, signal_198}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_1553, signal_1552, signal_1551, signal_408}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_393 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({signal_929, signal_928, signal_927, signal_201}), .a ({signal_908, signal_907, signal_906, signal_195}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({signal_1556, signal_1555, signal_1554, signal_409}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_394 ( .s ({signal_7381, signal_7379, signal_7377, signal_7375}), .b ({1'b0, 1'b0, 1'b0, signal_7385}), .a ({signal_932, signal_931, signal_930, signal_202}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({signal_1559, signal_1558, signal_1557, signal_410}) ) ;
    buf_clk cell_913 ( .C ( clk ), .D ( signal_7394 ), .Q ( signal_7395 ) ) ;
    buf_clk cell_915 ( .C ( clk ), .D ( signal_7396 ), .Q ( signal_7397 ) ) ;
    buf_clk cell_917 ( .C ( clk ), .D ( signal_7398 ), .Q ( signal_7399 ) ) ;
    buf_clk cell_919 ( .C ( clk ), .D ( signal_7400 ), .Q ( signal_7401 ) ) ;
    buf_clk cell_921 ( .C ( clk ), .D ( signal_7402 ), .Q ( signal_7403 ) ) ;
    buf_clk cell_923 ( .C ( clk ), .D ( signal_7404 ), .Q ( signal_7405 ) ) ;
    buf_clk cell_925 ( .C ( clk ), .D ( signal_7406 ), .Q ( signal_7407 ) ) ;
    buf_clk cell_927 ( .C ( clk ), .D ( signal_7408 ), .Q ( signal_7409 ) ) ;
    buf_clk cell_929 ( .C ( clk ), .D ( signal_7410 ), .Q ( signal_7411 ) ) ;
    buf_clk cell_931 ( .C ( clk ), .D ( signal_7412 ), .Q ( signal_7413 ) ) ;
    buf_clk cell_933 ( .C ( clk ), .D ( signal_7414 ), .Q ( signal_7415 ) ) ;
    buf_clk cell_935 ( .C ( clk ), .D ( signal_7416 ), .Q ( signal_7417 ) ) ;
    buf_clk cell_937 ( .C ( clk ), .D ( signal_7418 ), .Q ( signal_7419 ) ) ;
    buf_clk cell_939 ( .C ( clk ), .D ( signal_7420 ), .Q ( signal_7421 ) ) ;
    buf_clk cell_941 ( .C ( clk ), .D ( signal_7422 ), .Q ( signal_7423 ) ) ;
    buf_clk cell_943 ( .C ( clk ), .D ( signal_7424 ), .Q ( signal_7425 ) ) ;
    buf_clk cell_945 ( .C ( clk ), .D ( signal_7426 ), .Q ( signal_7427 ) ) ;
    buf_clk cell_947 ( .C ( clk ), .D ( signal_7428 ), .Q ( signal_7429 ) ) ;
    buf_clk cell_949 ( .C ( clk ), .D ( signal_7430 ), .Q ( signal_7431 ) ) ;
    buf_clk cell_951 ( .C ( clk ), .D ( signal_7432 ), .Q ( signal_7433 ) ) ;
    buf_clk cell_953 ( .C ( clk ), .D ( signal_7434 ), .Q ( signal_7435 ) ) ;
    buf_clk cell_955 ( .C ( clk ), .D ( signal_7436 ), .Q ( signal_7437 ) ) ;
    buf_clk cell_957 ( .C ( clk ), .D ( signal_7438 ), .Q ( signal_7439 ) ) ;
    buf_clk cell_959 ( .C ( clk ), .D ( signal_7440 ), .Q ( signal_7441 ) ) ;
    buf_clk cell_961 ( .C ( clk ), .D ( signal_7442 ), .Q ( signal_7443 ) ) ;
    buf_clk cell_963 ( .C ( clk ), .D ( signal_7444 ), .Q ( signal_7445 ) ) ;
    buf_clk cell_965 ( .C ( clk ), .D ( signal_7446 ), .Q ( signal_7447 ) ) ;
    buf_clk cell_967 ( .C ( clk ), .D ( signal_7448 ), .Q ( signal_7449 ) ) ;
    buf_clk cell_969 ( .C ( clk ), .D ( signal_7450 ), .Q ( signal_7451 ) ) ;
    buf_clk cell_971 ( .C ( clk ), .D ( signal_7452 ), .Q ( signal_7453 ) ) ;
    buf_clk cell_973 ( .C ( clk ), .D ( signal_7454 ), .Q ( signal_7455 ) ) ;
    buf_clk cell_975 ( .C ( clk ), .D ( signal_7456 ), .Q ( signal_7457 ) ) ;
    buf_clk cell_977 ( .C ( clk ), .D ( signal_7458 ), .Q ( signal_7459 ) ) ;
    buf_clk cell_979 ( .C ( clk ), .D ( signal_7460 ), .Q ( signal_7461 ) ) ;
    buf_clk cell_981 ( .C ( clk ), .D ( signal_7462 ), .Q ( signal_7463 ) ) ;
    buf_clk cell_983 ( .C ( clk ), .D ( signal_7464 ), .Q ( signal_7465 ) ) ;
    buf_clk cell_985 ( .C ( clk ), .D ( signal_7466 ), .Q ( signal_7467 ) ) ;
    buf_clk cell_987 ( .C ( clk ), .D ( signal_7468 ), .Q ( signal_7469 ) ) ;
    buf_clk cell_989 ( .C ( clk ), .D ( signal_7470 ), .Q ( signal_7471 ) ) ;
    buf_clk cell_991 ( .C ( clk ), .D ( signal_7472 ), .Q ( signal_7473 ) ) ;
    buf_clk cell_993 ( .C ( clk ), .D ( signal_7474 ), .Q ( signal_7475 ) ) ;
    buf_clk cell_995 ( .C ( clk ), .D ( signal_7476 ), .Q ( signal_7477 ) ) ;
    buf_clk cell_997 ( .C ( clk ), .D ( signal_7478 ), .Q ( signal_7479 ) ) ;
    buf_clk cell_999 ( .C ( clk ), .D ( signal_7480 ), .Q ( signal_7481 ) ) ;
    buf_clk cell_1001 ( .C ( clk ), .D ( signal_7482 ), .Q ( signal_7483 ) ) ;
    buf_clk cell_1003 ( .C ( clk ), .D ( signal_7484 ), .Q ( signal_7485 ) ) ;
    buf_clk cell_1005 ( .C ( clk ), .D ( signal_7486 ), .Q ( signal_7487 ) ) ;
    buf_clk cell_1007 ( .C ( clk ), .D ( signal_7488 ), .Q ( signal_7489 ) ) ;
    buf_clk cell_1009 ( .C ( clk ), .D ( signal_7490 ), .Q ( signal_7491 ) ) ;
    buf_clk cell_1011 ( .C ( clk ), .D ( signal_7492 ), .Q ( signal_7493 ) ) ;
    buf_clk cell_1013 ( .C ( clk ), .D ( signal_7494 ), .Q ( signal_7495 ) ) ;
    buf_clk cell_1015 ( .C ( clk ), .D ( signal_7496 ), .Q ( signal_7497 ) ) ;
    buf_clk cell_1017 ( .C ( clk ), .D ( signal_7498 ), .Q ( signal_7499 ) ) ;
    buf_clk cell_1019 ( .C ( clk ), .D ( signal_7500 ), .Q ( signal_7501 ) ) ;
    buf_clk cell_1021 ( .C ( clk ), .D ( signal_7502 ), .Q ( signal_7503 ) ) ;
    buf_clk cell_1023 ( .C ( clk ), .D ( signal_7504 ), .Q ( signal_7505 ) ) ;
    buf_clk cell_1025 ( .C ( clk ), .D ( signal_7506 ), .Q ( signal_7507 ) ) ;
    buf_clk cell_1027 ( .C ( clk ), .D ( signal_7508 ), .Q ( signal_7509 ) ) ;
    buf_clk cell_1029 ( .C ( clk ), .D ( signal_7510 ), .Q ( signal_7511 ) ) ;
    buf_clk cell_1031 ( .C ( clk ), .D ( signal_7512 ), .Q ( signal_7513 ) ) ;
    buf_clk cell_1033 ( .C ( clk ), .D ( signal_7514 ), .Q ( signal_7515 ) ) ;
    buf_clk cell_1035 ( .C ( clk ), .D ( signal_7516 ), .Q ( signal_7517 ) ) ;
    buf_clk cell_1037 ( .C ( clk ), .D ( signal_7518 ), .Q ( signal_7519 ) ) ;
    buf_clk cell_1039 ( .C ( clk ), .D ( signal_7520 ), .Q ( signal_7521 ) ) ;
    buf_clk cell_1041 ( .C ( clk ), .D ( signal_7522 ), .Q ( signal_7523 ) ) ;
    buf_clk cell_1043 ( .C ( clk ), .D ( signal_7524 ), .Q ( signal_7525 ) ) ;
    buf_clk cell_1045 ( .C ( clk ), .D ( signal_7526 ), .Q ( signal_7527 ) ) ;
    buf_clk cell_1047 ( .C ( clk ), .D ( signal_7528 ), .Q ( signal_7529 ) ) ;
    buf_clk cell_1049 ( .C ( clk ), .D ( signal_7530 ), .Q ( signal_7531 ) ) ;
    buf_clk cell_1051 ( .C ( clk ), .D ( signal_7532 ), .Q ( signal_7533 ) ) ;
    buf_clk cell_1053 ( .C ( clk ), .D ( signal_7534 ), .Q ( signal_7535 ) ) ;
    buf_clk cell_1055 ( .C ( clk ), .D ( signal_7536 ), .Q ( signal_7537 ) ) ;
    buf_clk cell_1057 ( .C ( clk ), .D ( signal_7538 ), .Q ( signal_7539 ) ) ;
    buf_clk cell_1059 ( .C ( clk ), .D ( signal_7540 ), .Q ( signal_7541 ) ) ;
    buf_clk cell_1061 ( .C ( clk ), .D ( signal_7542 ), .Q ( signal_7543 ) ) ;
    buf_clk cell_1063 ( .C ( clk ), .D ( signal_7544 ), .Q ( signal_7545 ) ) ;
    buf_clk cell_1065 ( .C ( clk ), .D ( signal_7546 ), .Q ( signal_7547 ) ) ;
    buf_clk cell_1067 ( .C ( clk ), .D ( signal_7548 ), .Q ( signal_7549 ) ) ;
    buf_clk cell_1069 ( .C ( clk ), .D ( signal_7550 ), .Q ( signal_7551 ) ) ;
    buf_clk cell_1071 ( .C ( clk ), .D ( signal_7552 ), .Q ( signal_7553 ) ) ;
    buf_clk cell_1073 ( .C ( clk ), .D ( signal_7554 ), .Q ( signal_7555 ) ) ;
    buf_clk cell_1075 ( .C ( clk ), .D ( signal_7556 ), .Q ( signal_7557 ) ) ;
    buf_clk cell_1077 ( .C ( clk ), .D ( signal_7558 ), .Q ( signal_7559 ) ) ;
    buf_clk cell_1079 ( .C ( clk ), .D ( signal_7560 ), .Q ( signal_7561 ) ) ;
    buf_clk cell_1081 ( .C ( clk ), .D ( signal_7562 ), .Q ( signal_7563 ) ) ;
    buf_clk cell_1083 ( .C ( clk ), .D ( signal_7564 ), .Q ( signal_7565 ) ) ;
    buf_clk cell_1087 ( .C ( clk ), .D ( signal_7568 ), .Q ( signal_7569 ) ) ;
    buf_clk cell_1093 ( .C ( clk ), .D ( signal_7574 ), .Q ( signal_7575 ) ) ;
    buf_clk cell_1099 ( .C ( clk ), .D ( signal_7580 ), .Q ( signal_7581 ) ) ;
    buf_clk cell_1105 ( .C ( clk ), .D ( signal_7586 ), .Q ( signal_7587 ) ) ;
    buf_clk cell_1127 ( .C ( clk ), .D ( signal_7608 ), .Q ( signal_7609 ) ) ;
    buf_clk cell_1135 ( .C ( clk ), .D ( signal_7616 ), .Q ( signal_7617 ) ) ;
    buf_clk cell_1143 ( .C ( clk ), .D ( signal_7624 ), .Q ( signal_7625 ) ) ;
    buf_clk cell_1151 ( .C ( clk ), .D ( signal_7632 ), .Q ( signal_7633 ) ) ;
    buf_clk cell_1159 ( .C ( clk ), .D ( signal_7640 ), .Q ( signal_7641 ) ) ;
    buf_clk cell_1169 ( .C ( clk ), .D ( signal_7650 ), .Q ( signal_7651 ) ) ;
    buf_clk cell_1179 ( .C ( clk ), .D ( signal_7660 ), .Q ( signal_7661 ) ) ;
    buf_clk cell_1189 ( .C ( clk ), .D ( signal_7670 ), .Q ( signal_7671 ) ) ;
    buf_clk cell_1199 ( .C ( clk ), .D ( signal_7680 ), .Q ( signal_7681 ) ) ;
    buf_clk cell_1211 ( .C ( clk ), .D ( signal_7692 ), .Q ( signal_7693 ) ) ;
    buf_clk cell_1223 ( .C ( clk ), .D ( signal_7704 ), .Q ( signal_7705 ) ) ;
    buf_clk cell_1235 ( .C ( clk ), .D ( signal_7716 ), .Q ( signal_7717 ) ) ;
    buf_clk cell_1247 ( .C ( clk ), .D ( signal_7728 ), .Q ( signal_7729 ) ) ;
    buf_clk cell_1261 ( .C ( clk ), .D ( signal_7742 ), .Q ( signal_7743 ) ) ;
    buf_clk cell_1275 ( .C ( clk ), .D ( signal_7756 ), .Q ( signal_7757 ) ) ;
    buf_clk cell_1289 ( .C ( clk ), .D ( signal_7770 ), .Q ( signal_7771 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_1088 ( .C ( clk ), .D ( signal_7569 ), .Q ( signal_7570 ) ) ;
    buf_clk cell_1094 ( .C ( clk ), .D ( signal_7575 ), .Q ( signal_7576 ) ) ;
    buf_clk cell_1100 ( .C ( clk ), .D ( signal_7581 ), .Q ( signal_7582 ) ) ;
    buf_clk cell_1106 ( .C ( clk ), .D ( signal_7587 ), .Q ( signal_7588 ) ) ;
    buf_clk cell_1108 ( .C ( clk ), .D ( signal_334 ), .Q ( signal_7590 ) ) ;
    buf_clk cell_1110 ( .C ( clk ), .D ( signal_1329 ), .Q ( signal_7592 ) ) ;
    buf_clk cell_1112 ( .C ( clk ), .D ( signal_1330 ), .Q ( signal_7594 ) ) ;
    buf_clk cell_1114 ( .C ( clk ), .D ( signal_1331 ), .Q ( signal_7596 ) ) ;
    buf_clk cell_1116 ( .C ( clk ), .D ( signal_404 ), .Q ( signal_7598 ) ) ;
    buf_clk cell_1118 ( .C ( clk ), .D ( signal_1539 ), .Q ( signal_7600 ) ) ;
    buf_clk cell_1120 ( .C ( clk ), .D ( signal_1540 ), .Q ( signal_7602 ) ) ;
    buf_clk cell_1122 ( .C ( clk ), .D ( signal_1541 ), .Q ( signal_7604 ) ) ;
    buf_clk cell_1128 ( .C ( clk ), .D ( signal_7609 ), .Q ( signal_7610 ) ) ;
    buf_clk cell_1136 ( .C ( clk ), .D ( signal_7617 ), .Q ( signal_7618 ) ) ;
    buf_clk cell_1144 ( .C ( clk ), .D ( signal_7625 ), .Q ( signal_7626 ) ) ;
    buf_clk cell_1152 ( .C ( clk ), .D ( signal_7633 ), .Q ( signal_7634 ) ) ;
    buf_clk cell_1160 ( .C ( clk ), .D ( signal_7641 ), .Q ( signal_7642 ) ) ;
    buf_clk cell_1170 ( .C ( clk ), .D ( signal_7651 ), .Q ( signal_7652 ) ) ;
    buf_clk cell_1180 ( .C ( clk ), .D ( signal_7661 ), .Q ( signal_7662 ) ) ;
    buf_clk cell_1190 ( .C ( clk ), .D ( signal_7671 ), .Q ( signal_7672 ) ) ;
    buf_clk cell_1200 ( .C ( clk ), .D ( signal_7681 ), .Q ( signal_7682 ) ) ;
    buf_clk cell_1212 ( .C ( clk ), .D ( signal_7693 ), .Q ( signal_7694 ) ) ;
    buf_clk cell_1224 ( .C ( clk ), .D ( signal_7705 ), .Q ( signal_7706 ) ) ;
    buf_clk cell_1236 ( .C ( clk ), .D ( signal_7717 ), .Q ( signal_7718 ) ) ;
    buf_clk cell_1248 ( .C ( clk ), .D ( signal_7729 ), .Q ( signal_7730 ) ) ;
    buf_clk cell_1262 ( .C ( clk ), .D ( signal_7743 ), .Q ( signal_7744 ) ) ;
    buf_clk cell_1276 ( .C ( clk ), .D ( signal_7757 ), .Q ( signal_7758 ) ) ;
    buf_clk cell_1290 ( .C ( clk ), .D ( signal_7771 ), .Q ( signal_7772 ) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_264 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_962, signal_961, signal_960, signal_212}), .a ({signal_7409, signal_7407, signal_7405, signal_7403}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({signal_1169, signal_1168, signal_1167, signal_280}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_322 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_977, signal_976, signal_975, signal_217}), .a ({signal_962, signal_961, signal_960, signal_212}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({signal_1343, signal_1342, signal_1341, signal_338}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_325 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_971, signal_970, signal_969, signal_215}), .a ({signal_7417, signal_7415, signal_7413, signal_7411}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_1352, signal_1351, signal_1350, signal_341}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_329 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_947, signal_946, signal_945, signal_207}), .a ({signal_7425, signal_7423, signal_7421, signal_7419}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({signal_1364, signal_1363, signal_1362, signal_345}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_395 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1010, signal_1009, signal_1008, signal_228}), .a ({signal_7433, signal_7431, signal_7429, signal_7427}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({signal_1562, signal_1561, signal_1560, signal_411}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_396 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1025, signal_1024, signal_1023, signal_233}), .a ({signal_1022, signal_1021, signal_1020, signal_232}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({signal_1565, signal_1564, signal_1563, signal_412}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_397 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1031, signal_1030, signal_1029, signal_235}), .a ({signal_1028, signal_1027, signal_1026, signal_234}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({signal_1568, signal_1567, signal_1566, signal_413}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_398 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1034, signal_1033, signal_1032, signal_236}), .a ({signal_7441, signal_7439, signal_7437, signal_7435}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_1571, signal_1570, signal_1569, signal_414}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_399 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1040, signal_1039, signal_1038, signal_238}), .a ({signal_1037, signal_1036, signal_1035, signal_237}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({signal_1574, signal_1573, signal_1572, signal_415}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_400 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1025, signal_1024, signal_1023, signal_233}), .a ({signal_1043, signal_1042, signal_1041, signal_239}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({signal_1577, signal_1576, signal_1575, signal_416}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_401 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1049, signal_1048, signal_1047, signal_241}), .a ({signal_1046, signal_1045, signal_1044, signal_240}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({signal_1580, signal_1579, signal_1578, signal_417}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_402 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1055, signal_1054, signal_1053, signal_243}), .a ({signal_1052, signal_1051, signal_1050, signal_242}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({signal_1583, signal_1582, signal_1581, signal_418}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_403 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1022, signal_1021, signal_1020, signal_232}), .a ({signal_1058, signal_1057, signal_1056, signal_244}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_1586, signal_1585, signal_1584, signal_419}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_404 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1061, signal_1060, signal_1059, signal_245}), .a ({signal_1028, signal_1027, signal_1026, signal_234}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({signal_1589, signal_1588, signal_1587, signal_420}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_405 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1067, signal_1066, signal_1065, signal_247}), .a ({signal_1064, signal_1063, signal_1062, signal_246}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({signal_1592, signal_1591, signal_1590, signal_421}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_406 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1070, signal_1069, signal_1068, signal_248}), .a ({signal_947, signal_946, signal_945, signal_207}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({signal_1595, signal_1594, signal_1593, signal_422}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_407 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1076, signal_1075, signal_1074, signal_250}), .a ({signal_1073, signal_1072, signal_1071, signal_249}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({signal_1598, signal_1597, signal_1596, signal_423}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_408 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1082, signal_1081, signal_1080, signal_252}), .a ({signal_1079, signal_1078, signal_1077, signal_251}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_1601, signal_1600, signal_1599, signal_424}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_409 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1085, signal_1084, signal_1083, signal_253}), .a ({1'b0, 1'b0, 1'b0, signal_7443}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({signal_1604, signal_1603, signal_1602, signal_425}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_410 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7451, signal_7449, signal_7447, signal_7445}), .a ({signal_1088, signal_1087, signal_1086, signal_254}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({signal_1607, signal_1606, signal_1605, signal_426}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_411 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1094, signal_1093, signal_1092, signal_256}), .a ({signal_1091, signal_1090, signal_1089, signal_255}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({signal_1610, signal_1609, signal_1608, signal_427}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_412 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1097, signal_1096, signal_1095, signal_257}), .a ({signal_1043, signal_1042, signal_1041, signal_239}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({signal_1613, signal_1612, signal_1611, signal_428}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_413 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_947, signal_946, signal_945, signal_207}), .a ({signal_1100, signal_1099, signal_1098, signal_258}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_1616, signal_1615, signal_1614, signal_429}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_414 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1106, signal_1105, signal_1104, signal_260}), .a ({signal_1103, signal_1102, signal_1101, signal_259}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({signal_1619, signal_1618, signal_1617, signal_430}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_415 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1112, signal_1111, signal_1110, signal_262}), .a ({signal_1109, signal_1108, signal_1107, signal_261}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({signal_1622, signal_1621, signal_1620, signal_431}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_416 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7459, signal_7457, signal_7455, signal_7453}), .a ({signal_1115, signal_1114, signal_1113, signal_263}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({signal_1625, signal_1624, signal_1623, signal_432}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_417 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1121, signal_1120, signal_1119, signal_265}), .a ({signal_1118, signal_1117, signal_1116, signal_264}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({signal_1628, signal_1627, signal_1626, signal_433}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_418 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7467, signal_7465, signal_7463, signal_7461}), .a ({signal_1124, signal_1123, signal_1122, signal_266}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_1631, signal_1630, signal_1629, signal_434}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_419 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7475, signal_7473, signal_7471, signal_7469}), .a ({signal_1127, signal_1126, signal_1125, signal_267}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({signal_1634, signal_1633, signal_1632, signal_435}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_420 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1133, signal_1132, signal_1131, signal_269}), .a ({signal_1130, signal_1129, signal_1128, signal_268}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({signal_1637, signal_1636, signal_1635, signal_436}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_421 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1139, signal_1138, signal_1137, signal_271}), .a ({signal_1136, signal_1135, signal_1134, signal_270}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({signal_1640, signal_1639, signal_1638, signal_437}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_422 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1145, signal_1144, signal_1143, signal_273}), .a ({signal_1142, signal_1141, signal_1140, signal_272}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({signal_1643, signal_1642, signal_1641, signal_438}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_423 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1151, signal_1150, signal_1149, signal_275}), .a ({signal_1148, signal_1147, signal_1146, signal_274}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_1646, signal_1645, signal_1644, signal_439}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_424 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1154, signal_1153, signal_1152, signal_276}), .a ({signal_7483, signal_7481, signal_7479, signal_7477}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({signal_1649, signal_1648, signal_1647, signal_440}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_425 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1079, signal_1078, signal_1077, signal_251}), .a ({signal_1157, signal_1156, signal_1155, signal_277}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({signal_1652, signal_1651, signal_1650, signal_441}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_426 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1160, signal_1159, signal_1158, signal_278}), .a ({signal_1157, signal_1156, signal_1155, signal_277}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({signal_1655, signal_1654, signal_1653, signal_442}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_427 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1163, signal_1162, signal_1161, signal_279}), .a ({signal_1139, signal_1138, signal_1137, signal_271}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({signal_1658, signal_1657, signal_1656, signal_443}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_428 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1076, signal_1075, signal_1074, signal_250}), .a ({signal_1172, signal_1171, signal_1170, signal_281}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_1661, signal_1660, signal_1659, signal_444}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_429 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1178, signal_1177, signal_1176, signal_283}), .a ({signal_1175, signal_1174, signal_1173, signal_282}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({signal_1664, signal_1663, signal_1662, signal_445}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_430 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1184, signal_1183, signal_1182, signal_285}), .a ({signal_1181, signal_1180, signal_1179, signal_284}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({signal_1667, signal_1666, signal_1665, signal_446}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_431 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1187, signal_1186, signal_1185, signal_286}), .a ({signal_965, signal_964, signal_963, signal_213}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({signal_1670, signal_1669, signal_1668, signal_447}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_432 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1112, signal_1111, signal_1110, signal_262}), .a ({signal_1139, signal_1138, signal_1137, signal_271}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({signal_1673, signal_1672, signal_1671, signal_448}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_433 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1193, signal_1192, signal_1191, signal_288}), .a ({signal_1190, signal_1189, signal_1188, signal_287}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_1676, signal_1675, signal_1674, signal_449}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_434 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_965, signal_964, signal_963, signal_213}), .a ({signal_1100, signal_1099, signal_1098, signal_258}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({signal_1679, signal_1678, signal_1677, signal_450}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_435 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1199, signal_1198, signal_1197, signal_290}), .a ({signal_1196, signal_1195, signal_1194, signal_289}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({signal_1682, signal_1681, signal_1680, signal_451}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_436 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1094, signal_1093, signal_1092, signal_256}), .a ({signal_1181, signal_1180, signal_1179, signal_284}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({signal_1685, signal_1684, signal_1683, signal_452}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_437 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1130, signal_1129, signal_1128, signal_268}), .a ({signal_1202, signal_1201, signal_1200, signal_291}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({signal_1688, signal_1687, signal_1686, signal_453}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_438 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1160, signal_1159, signal_1158, signal_278}), .a ({signal_1205, signal_1204, signal_1203, signal_292}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_1691, signal_1690, signal_1689, signal_454}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_439 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1208, signal_1207, signal_1206, signal_293}), .a ({signal_7425, signal_7423, signal_7421, signal_7419}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({signal_1694, signal_1693, signal_1692, signal_455}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_440 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1214, signal_1213, signal_1212, signal_295}), .a ({signal_1211, signal_1210, signal_1209, signal_294}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({signal_1697, signal_1696, signal_1695, signal_456}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_441 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1157, signal_1156, signal_1155, signal_277}), .a ({signal_1217, signal_1216, signal_1215, signal_296}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({signal_1700, signal_1699, signal_1698, signal_457}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_442 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1220, signal_1219, signal_1218, signal_297}), .a ({signal_971, signal_970, signal_969, signal_215}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({signal_1703, signal_1702, signal_1701, signal_458}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_443 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1223, signal_1222, signal_1221, signal_298}), .a ({signal_974, signal_973, signal_972, signal_216}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_1706, signal_1705, signal_1704, signal_459}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_444 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1226, signal_1225, signal_1224, signal_299}), .a ({signal_1073, signal_1072, signal_1071, signal_249}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({signal_1709, signal_1708, signal_1707, signal_460}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_445 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1232, signal_1231, signal_1230, signal_301}), .a ({signal_1229, signal_1228, signal_1227, signal_300}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({signal_1712, signal_1711, signal_1710, signal_461}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_446 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1139, signal_1138, signal_1137, signal_271}), .a ({signal_1235, signal_1234, signal_1233, signal_302}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({signal_1715, signal_1714, signal_1713, signal_462}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_447 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1241, signal_1240, signal_1239, signal_304}), .a ({signal_1238, signal_1237, signal_1236, signal_303}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({signal_1718, signal_1717, signal_1716, signal_463}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_448 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1127, signal_1126, signal_1125, signal_267}), .a ({signal_962, signal_961, signal_960, signal_212}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_1721, signal_1720, signal_1719, signal_464}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_449 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({1'b0, 1'b0, 1'b0, signal_7485}), .a ({signal_1148, signal_1147, signal_1146, signal_274}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({signal_1724, signal_1723, signal_1722, signal_465}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_450 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7451, signal_7449, signal_7447, signal_7445}), .a ({signal_1052, signal_1051, signal_1050, signal_242}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({signal_1727, signal_1726, signal_1725, signal_466}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_451 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1244, signal_1243, signal_1242, signal_305}), .a ({signal_1151, signal_1150, signal_1149, signal_275}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({signal_1730, signal_1729, signal_1728, signal_467}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_452 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1250, signal_1249, signal_1248, signal_307}), .a ({signal_1247, signal_1246, signal_1245, signal_306}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({signal_1733, signal_1732, signal_1731, signal_468}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_453 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1253, signal_1252, signal_1251, signal_308}), .a ({1'b0, 1'b0, 1'b0, signal_7443}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_1736, signal_1735, signal_1734, signal_469}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_454 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1163, signal_1162, signal_1161, signal_279}), .a ({signal_977, signal_976, signal_975, signal_217}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({signal_1739, signal_1738, signal_1737, signal_470}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_455 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1079, signal_1078, signal_1077, signal_251}), .a ({signal_1229, signal_1228, signal_1227, signal_300}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({signal_1742, signal_1741, signal_1740, signal_471}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_456 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1256, signal_1255, signal_1254, signal_309}), .a ({signal_7493, signal_7491, signal_7489, signal_7487}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({signal_1745, signal_1744, signal_1743, signal_472}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_457 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1262, signal_1261, signal_1260, signal_311}), .a ({signal_1259, signal_1258, signal_1257, signal_310}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({signal_1748, signal_1747, signal_1746, signal_473}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_458 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1265, signal_1264, signal_1263, signal_312}), .a ({signal_1151, signal_1150, signal_1149, signal_275}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_1751, signal_1750, signal_1749, signal_474}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_459 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1271, signal_1270, signal_1269, signal_314}), .a ({signal_1268, signal_1267, signal_1266, signal_313}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({signal_1754, signal_1753, signal_1752, signal_475}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_460 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1277, signal_1276, signal_1275, signal_316}), .a ({signal_1274, signal_1273, signal_1272, signal_315}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({signal_1757, signal_1756, signal_1755, signal_476}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_461 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1280, signal_1279, signal_1278, signal_317}), .a ({signal_1121, signal_1120, signal_1119, signal_265}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({signal_1760, signal_1759, signal_1758, signal_477}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_462 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1286, signal_1285, signal_1284, signal_319}), .a ({signal_1283, signal_1282, signal_1281, signal_318}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({signal_1763, signal_1762, signal_1761, signal_478}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_463 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1043, signal_1042, signal_1041, signal_239}), .a ({signal_1289, signal_1288, signal_1287, signal_320}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_1766, signal_1765, signal_1764, signal_479}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_464 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1139, signal_1138, signal_1137, signal_271}), .a ({signal_1292, signal_1291, signal_1290, signal_321}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({signal_1769, signal_1768, signal_1767, signal_480}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_465 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1298, signal_1297, signal_1296, signal_323}), .a ({signal_1295, signal_1294, signal_1293, signal_322}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({signal_1772, signal_1771, signal_1770, signal_481}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_466 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7433, signal_7431, signal_7429, signal_7427}), .a ({signal_1301, signal_1300, signal_1299, signal_324}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({signal_1775, signal_1774, signal_1773, signal_482}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_467 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1304, signal_1303, signal_1302, signal_325}), .a ({signal_7501, signal_7499, signal_7497, signal_7495}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({signal_1778, signal_1777, signal_1776, signal_483}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_468 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1310, signal_1309, signal_1308, signal_327}), .a ({signal_1307, signal_1306, signal_1305, signal_326}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_1781, signal_1780, signal_1779, signal_484}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_469 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1022, signal_1021, signal_1020, signal_232}), .a ({signal_1196, signal_1195, signal_1194, signal_289}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({signal_1784, signal_1783, signal_1782, signal_485}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_470 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1313, signal_1312, signal_1311, signal_328}), .a ({signal_1160, signal_1159, signal_1158, signal_278}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({signal_1787, signal_1786, signal_1785, signal_486}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_471 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1064, signal_1063, signal_1062, signal_246}), .a ({signal_7509, signal_7507, signal_7505, signal_7503}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({signal_1790, signal_1789, signal_1788, signal_487}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_472 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1118, signal_1117, signal_1116, signal_264}), .a ({1'b0, 1'b0, 1'b0, signal_7443}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({signal_1793, signal_1792, signal_1791, signal_488}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_473 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1319, signal_1318, signal_1317, signal_330}), .a ({signal_1316, signal_1315, signal_1314, signal_329}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_1796, signal_1795, signal_1794, signal_489}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_474 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1121, signal_1120, signal_1119, signal_265}), .a ({signal_1322, signal_1321, signal_1320, signal_331}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({signal_1799, signal_1798, signal_1797, signal_490}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_475 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1316, signal_1315, signal_1314, signal_329}), .a ({signal_1205, signal_1204, signal_1203, signal_292}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({signal_1802, signal_1801, signal_1800, signal_491}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_476 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1325, signal_1324, signal_1323, signal_332}), .a ({signal_1100, signal_1099, signal_1098, signal_258}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({signal_1805, signal_1804, signal_1803, signal_492}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_477 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1328, signal_1327, signal_1326, signal_333}), .a ({signal_1148, signal_1147, signal_1146, signal_274}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({signal_1808, signal_1807, signal_1806, signal_493}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_478 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1205, signal_1204, signal_1203, signal_292}), .a ({signal_1331, signal_1330, signal_1329, signal_334}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_1811, signal_1810, signal_1809, signal_494}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_479 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1334, signal_1333, signal_1332, signal_335}), .a ({signal_7441, signal_7439, signal_7437, signal_7435}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({signal_1814, signal_1813, signal_1812, signal_495}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_480 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1337, signal_1336, signal_1335, signal_336}), .a ({signal_1070, signal_1069, signal_1068, signal_248}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({signal_1817, signal_1816, signal_1815, signal_496}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_481 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1334, signal_1333, signal_1332, signal_335}), .a ({signal_1118, signal_1117, signal_1116, signal_264}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({signal_1820, signal_1819, signal_1818, signal_497}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_482 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1187, signal_1186, signal_1185, signal_286}), .a ({signal_1340, signal_1339, signal_1338, signal_337}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({signal_1823, signal_1822, signal_1821, signal_498}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_483 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_986, signal_985, signal_984, signal_220}), .a ({signal_1055, signal_1054, signal_1053, signal_243}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_1826, signal_1825, signal_1824, signal_499}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_484 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1256, signal_1255, signal_1254, signal_309}), .a ({signal_1196, signal_1195, signal_1194, signal_289}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({signal_1829, signal_1828, signal_1827, signal_500}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_485 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1349, signal_1348, signal_1347, signal_340}), .a ({signal_1346, signal_1345, signal_1344, signal_339}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({signal_1832, signal_1831, signal_1830, signal_501}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_486 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1337, signal_1336, signal_1335, signal_336}), .a ({signal_1049, signal_1048, signal_1047, signal_241}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({signal_1835, signal_1834, signal_1833, signal_502}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_487 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1214, signal_1213, signal_1212, signal_295}), .a ({signal_1064, signal_1063, signal_1062, signal_246}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({signal_1838, signal_1837, signal_1836, signal_503}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_488 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1280, signal_1279, signal_1278, signal_317}), .a ({signal_1079, signal_1078, signal_1077, signal_251}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_1841, signal_1840, signal_1839, signal_504}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_489 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_989, signal_988, signal_987, signal_221}), .a ({signal_1187, signal_1186, signal_1185, signal_286}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({signal_1844, signal_1843, signal_1842, signal_505}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_490 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1163, signal_1162, signal_1161, signal_279}), .a ({signal_1238, signal_1237, signal_1236, signal_303}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({signal_1847, signal_1846, signal_1845, signal_506}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_491 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1130, signal_1129, signal_1128, signal_268}), .a ({signal_1142, signal_1141, signal_1140, signal_272}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({signal_1850, signal_1849, signal_1848, signal_507}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_492 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1148, signal_1147, signal_1146, signal_274}), .a ({signal_1124, signal_1123, signal_1122, signal_266}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({signal_1853, signal_1852, signal_1851, signal_508}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_493 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1358, signal_1357, signal_1356, signal_343}), .a ({signal_1355, signal_1354, signal_1353, signal_342}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_1856, signal_1855, signal_1854, signal_509}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_494 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1361, signal_1360, signal_1359, signal_344}), .a ({signal_1277, signal_1276, signal_1275, signal_316}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({signal_1859, signal_1858, signal_1857, signal_510}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_495 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1244, signal_1243, signal_1242, signal_305}), .a ({signal_986, signal_985, signal_984, signal_220}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({signal_1862, signal_1861, signal_1860, signal_511}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_496 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1328, signal_1327, signal_1326, signal_333}), .a ({signal_1367, signal_1366, signal_1365, signal_346}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({signal_1865, signal_1864, signal_1863, signal_512}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_497 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1268, signal_1267, signal_1266, signal_313}), .a ({signal_1142, signal_1141, signal_1140, signal_272}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({signal_1868, signal_1867, signal_1866, signal_513}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_498 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1214, signal_1213, signal_1212, signal_295}), .a ({signal_1097, signal_1096, signal_1095, signal_257}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_1871, signal_1870, signal_1869, signal_514}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_499 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1271, signal_1270, signal_1269, signal_314}), .a ({signal_1328, signal_1327, signal_1326, signal_333}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({signal_1874, signal_1873, signal_1872, signal_515}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_500 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1223, signal_1222, signal_1221, signal_298}), .a ({signal_1319, signal_1318, signal_1317, signal_330}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({signal_1877, signal_1876, signal_1875, signal_516}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_501 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1373, signal_1372, signal_1371, signal_348}), .a ({signal_1370, signal_1369, signal_1368, signal_347}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({signal_1880, signal_1879, signal_1878, signal_517}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_502 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7517, signal_7515, signal_7513, signal_7511}), .a ({signal_1085, signal_1084, signal_1083, signal_253}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({signal_1883, signal_1882, signal_1881, signal_518}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_503 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1376, signal_1375, signal_1374, signal_349}), .a ({signal_992, signal_991, signal_990, signal_222}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_1886, signal_1885, signal_1884, signal_519}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_504 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1379, signal_1378, signal_1377, signal_350}), .a ({signal_1361, signal_1360, signal_1359, signal_344}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({signal_1889, signal_1888, signal_1887, signal_520}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_505 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1325, signal_1324, signal_1323, signal_332}), .a ({signal_1382, signal_1381, signal_1380, signal_351}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({signal_1892, signal_1891, signal_1890, signal_521}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_506 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1112, signal_1111, signal_1110, signal_262}), .a ({signal_1385, signal_1384, signal_1383, signal_352}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({signal_1895, signal_1894, signal_1893, signal_522}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_507 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1388, signal_1387, signal_1386, signal_353}), .a ({signal_1046, signal_1045, signal_1044, signal_240}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({signal_1898, signal_1897, signal_1896, signal_523}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_508 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1391, signal_1390, signal_1389, signal_354}), .a ({signal_1301, signal_1300, signal_1299, signal_324}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_1901, signal_1900, signal_1899, signal_524}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_509 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1394, signal_1393, signal_1392, signal_355}), .a ({signal_7441, signal_7439, signal_7437, signal_7435}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({signal_1904, signal_1903, signal_1902, signal_525}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_510 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1361, signal_1360, signal_1359, signal_344}), .a ({signal_1397, signal_1396, signal_1395, signal_356}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({signal_1907, signal_1906, signal_1905, signal_526}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_511 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1400, signal_1399, signal_1398, signal_357}), .a ({signal_1178, signal_1177, signal_1176, signal_283}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({signal_1910, signal_1909, signal_1908, signal_527}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_512 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7525, signal_7523, signal_7521, signal_7519}), .a ({signal_1403, signal_1402, signal_1401, signal_358}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({signal_1913, signal_1912, signal_1911, signal_528}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_513 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7533, signal_7531, signal_7529, signal_7527}), .a ({signal_1175, signal_1174, signal_1173, signal_282}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_1916, signal_1915, signal_1914, signal_529}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_514 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1076, signal_1075, signal_1074, signal_250}), .a ({signal_1406, signal_1405, signal_1404, signal_359}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({signal_1919, signal_1918, signal_1917, signal_530}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_515 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_998, signal_997, signal_996, signal_224}), .a ({signal_1247, signal_1246, signal_1245, signal_306}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({signal_1922, signal_1921, signal_1920, signal_531}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_516 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1412, signal_1411, signal_1410, signal_361}), .a ({signal_1409, signal_1408, signal_1407, signal_360}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({signal_1925, signal_1924, signal_1923, signal_532}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_517 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1265, signal_1264, signal_1263, signal_312}), .a ({signal_1415, signal_1414, signal_1413, signal_362}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({signal_1928, signal_1927, signal_1926, signal_533}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_518 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1421, signal_1420, signal_1419, signal_364}), .a ({signal_1418, signal_1417, signal_1416, signal_363}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_1931, signal_1930, signal_1929, signal_534}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_519 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1100, signal_1099, signal_1098, signal_258}), .a ({signal_1280, signal_1279, signal_1278, signal_317}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({signal_1934, signal_1933, signal_1932, signal_535}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_520 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1424, signal_1423, signal_1422, signal_365}), .a ({signal_1346, signal_1345, signal_1344, signal_339}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({signal_1937, signal_1936, signal_1935, signal_536}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_521 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1253, signal_1252, signal_1251, signal_308}), .a ({signal_1427, signal_1426, signal_1425, signal_366}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({signal_1940, signal_1939, signal_1938, signal_537}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_522 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7541, signal_7539, signal_7537, signal_7535}), .a ({signal_1100, signal_1099, signal_1098, signal_258}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({signal_1943, signal_1942, signal_1941, signal_538}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_523 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1139, signal_1138, signal_1137, signal_271}), .a ({signal_1226, signal_1225, signal_1224, signal_299}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_1946, signal_1945, signal_1944, signal_539}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_524 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1145, signal_1144, signal_1143, signal_273}), .a ({signal_1283, signal_1282, signal_1281, signal_318}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({signal_1949, signal_1948, signal_1947, signal_540}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_525 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1178, signal_1177, signal_1176, signal_283}), .a ({signal_1181, signal_1180, signal_1179, signal_284}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({signal_1952, signal_1951, signal_1950, signal_541}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_526 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1433, signal_1432, signal_1431, signal_368}), .a ({signal_1430, signal_1429, signal_1428, signal_367}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({signal_1955, signal_1954, signal_1953, signal_542}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_527 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1436, signal_1435, signal_1434, signal_369}), .a ({signal_1418, signal_1417, signal_1416, signal_363}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({signal_1958, signal_1957, signal_1956, signal_543}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_528 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1043, signal_1042, signal_1041, signal_239}), .a ({signal_1295, signal_1294, signal_1293, signal_322}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_1961, signal_1960, signal_1959, signal_544}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_529 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1004, signal_1003, signal_1002, signal_226}), .a ({signal_1439, signal_1438, signal_1437, signal_370}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({signal_1964, signal_1963, signal_1962, signal_545}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_530 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_998, signal_997, signal_996, signal_224}), .a ({signal_1442, signal_1441, signal_1440, signal_371}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({signal_1967, signal_1966, signal_1965, signal_546}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_531 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1445, signal_1444, signal_1443, signal_372}), .a ({signal_1337, signal_1336, signal_1335, signal_336}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({signal_1970, signal_1969, signal_1968, signal_547}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_532 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1079, signal_1078, signal_1077, signal_251}), .a ({signal_1244, signal_1243, signal_1242, signal_305}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({signal_1973, signal_1972, signal_1971, signal_548}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_533 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1394, signal_1393, signal_1392, signal_355}), .a ({signal_1007, signal_1006, signal_1005, signal_227}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_1976, signal_1975, signal_1974, signal_549}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_534 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7433, signal_7431, signal_7429, signal_7427}), .a ({signal_1448, signal_1447, signal_1446, signal_373}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({signal_1979, signal_1978, signal_1977, signal_550}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_535 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1004, signal_1003, signal_1002, signal_226}), .a ({signal_1064, signal_1063, signal_1062, signal_246}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({signal_1982, signal_1981, signal_1980, signal_551}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_536 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1010, signal_1009, signal_1008, signal_228}), .a ({signal_1451, signal_1450, signal_1449, signal_374}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({signal_1985, signal_1984, signal_1983, signal_552}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_537 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1454, signal_1453, signal_1452, signal_375}), .a ({signal_1451, signal_1450, signal_1449, signal_374}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({signal_1988, signal_1987, signal_1986, signal_553}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_538 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7451, signal_7449, signal_7447, signal_7445}), .a ({signal_1124, signal_1123, signal_1122, signal_266}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_1991, signal_1990, signal_1989, signal_554}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_539 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1175, signal_1174, signal_1173, signal_282}), .a ({signal_1103, signal_1102, signal_1101, signal_259}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({signal_1994, signal_1993, signal_1992, signal_555}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_540 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1457, signal_1456, signal_1455, signal_376}), .a ({signal_1007, signal_1006, signal_1005, signal_227}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({signal_1997, signal_1996, signal_1995, signal_556}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_541 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1256, signal_1255, signal_1254, signal_309}), .a ({signal_1460, signal_1459, signal_1458, signal_377}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({signal_2000, signal_1999, signal_1998, signal_557}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_542 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7549, signal_7547, signal_7545, signal_7543}), .a ({signal_1202, signal_1201, signal_1200, signal_291}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({signal_2003, signal_2002, signal_2001, signal_558}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_543 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1115, signal_1114, signal_1113, signal_263}), .a ({signal_1235, signal_1234, signal_1233, signal_302}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_2006, signal_2005, signal_2004, signal_559}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_544 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1070, signal_1069, signal_1068, signal_248}), .a ({signal_1271, signal_1270, signal_1269, signal_314}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({signal_2009, signal_2008, signal_2007, signal_560}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_545 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1463, signal_1462, signal_1461, signal_378}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({signal_2012, signal_2011, signal_2010, signal_561}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_546 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1154, signal_1153, signal_1152, signal_276}), .a ({signal_1451, signal_1450, signal_1449, signal_374}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({signal_2015, signal_2014, signal_2013, signal_562}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_547 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1172, signal_1171, signal_1170, signal_281}), .a ({signal_1304, signal_1303, signal_1302, signal_325}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({signal_2018, signal_2017, signal_2016, signal_563}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_548 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1469, signal_1468, signal_1467, signal_380}), .a ({signal_1466, signal_1465, signal_1464, signal_379}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_2021, signal_2020, signal_2019, signal_564}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_549 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1394, signal_1393, signal_1392, signal_355}), .a ({signal_1349, signal_1348, signal_1347, signal_340}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({signal_2024, signal_2023, signal_2022, signal_565}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_550 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1472, signal_1471, signal_1470, signal_381}), .a ({signal_1442, signal_1441, signal_1440, signal_371}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({signal_2027, signal_2026, signal_2025, signal_566}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_551 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1478, signal_1477, signal_1476, signal_383}), .a ({signal_1475, signal_1474, signal_1473, signal_382}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({signal_2030, signal_2029, signal_2028, signal_567}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_552 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1022, signal_1021, signal_1020, signal_232}), .a ({signal_7501, signal_7499, signal_7497, signal_7495}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({signal_2033, signal_2032, signal_2031, signal_568}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_553 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1406, signal_1405, signal_1404, signal_359}), .a ({signal_971, signal_970, signal_969, signal_215}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_2036, signal_2035, signal_2034, signal_569}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_554 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1325, signal_1324, signal_1323, signal_332}), .a ({signal_1481, signal_1480, signal_1479, signal_384}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({signal_2039, signal_2038, signal_2037, signal_570}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_555 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1415, signal_1414, signal_1413, signal_362}), .a ({signal_1073, signal_1072, signal_1071, signal_249}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({signal_2042, signal_2041, signal_2040, signal_571}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_556 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1244, signal_1243, signal_1242, signal_305}), .a ({signal_1286, signal_1285, signal_1284, signal_319}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({signal_2045, signal_2044, signal_2043, signal_572}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_557 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1319, signal_1318, signal_1317, signal_330}), .a ({signal_1136, signal_1135, signal_1134, signal_270}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({signal_2048, signal_2047, signal_2046, signal_573}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_558 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1397, signal_1396, signal_1395, signal_356}), .a ({signal_1484, signal_1483, signal_1482, signal_385}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_2051, signal_2050, signal_2049, signal_574}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_559 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7425, signal_7423, signal_7421, signal_7419}), .a ({signal_1280, signal_1279, signal_1278, signal_317}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({signal_2054, signal_2053, signal_2052, signal_575}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_560 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1067, signal_1066, signal_1065, signal_247}), .a ({signal_1052, signal_1051, signal_1050, signal_242}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({signal_2057, signal_2056, signal_2055, signal_576}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_561 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1265, signal_1264, signal_1263, signal_312}), .a ({signal_1217, signal_1216, signal_1215, signal_296}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({signal_2060, signal_2059, signal_2058, signal_577}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_562 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1118, signal_1117, signal_1116, signal_264}), .a ({signal_1283, signal_1282, signal_1281, signal_318}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({signal_2063, signal_2062, signal_2061, signal_578}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_563 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1487, signal_1486, signal_1485, signal_386}), .a ({signal_1136, signal_1135, signal_1134, signal_270}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_2066, signal_2065, signal_2064, signal_579}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_564 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1157, signal_1156, signal_1155, signal_277}), .a ({signal_7525, signal_7523, signal_7521, signal_7519}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({signal_2069, signal_2068, signal_2067, signal_580}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_565 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1409, signal_1408, signal_1407, signal_360}), .a ({signal_1415, signal_1414, signal_1413, signal_362}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({signal_2072, signal_2071, signal_2070, signal_581}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_566 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_989, signal_988, signal_987, signal_221}), .a ({signal_1490, signal_1489, signal_1488, signal_387}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({signal_2075, signal_2074, signal_2073, signal_582}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_567 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1337, signal_1336, signal_1335, signal_336}), .a ({signal_7525, signal_7523, signal_7521, signal_7519}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({signal_2078, signal_2077, signal_2076, signal_583}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_568 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1493, signal_1492, signal_1491, signal_388}), .a ({signal_1280, signal_1279, signal_1278, signal_317}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_2081, signal_2080, signal_2079, signal_584}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_569 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_998, signal_997, signal_996, signal_224}), .a ({signal_1373, signal_1372, signal_1371, signal_348}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({signal_2084, signal_2083, signal_2082, signal_585}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_570 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1496, signal_1495, signal_1494, signal_389}), .a ({signal_1313, signal_1312, signal_1311, signal_328}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({signal_2087, signal_2086, signal_2085, signal_586}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_571 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1499, signal_1498, signal_1497, signal_390}), .a ({signal_977, signal_976, signal_975, signal_217}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({signal_2090, signal_2089, signal_2088, signal_587}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_572 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1370, signal_1369, signal_1368, signal_347}), .a ({signal_1178, signal_1177, signal_1176, signal_283}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({signal_2093, signal_2092, signal_2091, signal_588}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_573 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1334, signal_1333, signal_1332, signal_335}), .a ({signal_1370, signal_1369, signal_1368, signal_347}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_2096, signal_2095, signal_2094, signal_589}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_574 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1394, signal_1393, signal_1392, signal_355}), .a ({signal_1346, signal_1345, signal_1344, signal_339}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({signal_2099, signal_2098, signal_2097, signal_590}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_575 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1049, signal_1048, signal_1047, signal_241}), .a ({signal_1202, signal_1201, signal_1200, signal_291}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({signal_2102, signal_2101, signal_2100, signal_591}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_576 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1391, signal_1390, signal_1389, signal_354}), .a ({signal_1466, signal_1465, signal_1464, signal_379}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({signal_2105, signal_2104, signal_2103, signal_592}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_577 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1463, signal_1462, signal_1461, signal_378}), .a ({signal_1241, signal_1240, signal_1239, signal_304}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({signal_2108, signal_2107, signal_2106, signal_593}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_578 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1013, signal_1012, signal_1011, signal_229}), .a ({signal_1196, signal_1195, signal_1194, signal_289}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_2111, signal_2110, signal_2109, signal_594}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_579 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1115, signal_1114, signal_1113, signal_263}), .a ({signal_1502, signal_1501, signal_1500, signal_391}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({signal_2114, signal_2113, signal_2112, signal_595}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_580 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1265, signal_1264, signal_1263, signal_312}), .a ({signal_1163, signal_1162, signal_1161, signal_279}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({signal_2117, signal_2116, signal_2115, signal_596}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_581 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1109, signal_1108, signal_1107, signal_261}), .a ({signal_1172, signal_1171, signal_1170, signal_281}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({signal_2120, signal_2119, signal_2118, signal_597}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_582 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1475, signal_1474, signal_1473, signal_382}), .a ({signal_1340, signal_1339, signal_1338, signal_337}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({signal_2123, signal_2122, signal_2121, signal_598}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_583 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1286, signal_1285, signal_1284, signal_319}), .a ({signal_1388, signal_1387, signal_1386, signal_353}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_2126, signal_2125, signal_2124, signal_599}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_584 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1499, signal_1498, signal_1497, signal_390}), .a ({signal_1463, signal_1462, signal_1461, signal_378}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({signal_2129, signal_2128, signal_2127, signal_600}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_585 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1256, signal_1255, signal_1254, signal_309}), .a ({signal_1037, signal_1036, signal_1035, signal_237}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({signal_2132, signal_2131, signal_2130, signal_601}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_586 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1379, signal_1378, signal_1377, signal_350}), .a ({signal_1406, signal_1405, signal_1404, signal_359}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({signal_2135, signal_2134, signal_2133, signal_602}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_587 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1508, signal_1507, signal_1506, signal_393}), .a ({signal_1505, signal_1504, signal_1503, signal_392}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({signal_2138, signal_2137, signal_2136, signal_603}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_588 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1304, signal_1303, signal_1302, signal_325}), .a ({signal_1511, signal_1510, signal_1509, signal_394}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_2141, signal_2140, signal_2139, signal_604}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_589 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_998, signal_997, signal_996, signal_224}), .a ({signal_1514, signal_1513, signal_1512, signal_395}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({signal_2144, signal_2143, signal_2142, signal_605}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_590 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1259, signal_1258, signal_1257, signal_310}), .a ({signal_7509, signal_7507, signal_7505, signal_7503}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({signal_2147, signal_2146, signal_2145, signal_606}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_591 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_971, signal_970, signal_969, signal_215}), .a ({signal_1382, signal_1381, signal_1380, signal_351}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({signal_2150, signal_2149, signal_2148, signal_607}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_592 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1349, signal_1348, signal_1347, signal_340}), .a ({signal_7409, signal_7407, signal_7405, signal_7403}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({signal_2153, signal_2152, signal_2151, signal_608}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_593 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1475, signal_1474, signal_1473, signal_382}), .a ({signal_1154, signal_1153, signal_1152, signal_276}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_2156, signal_2155, signal_2154, signal_609}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_594 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1436, signal_1435, signal_1434, signal_369}), .a ({signal_1442, signal_1441, signal_1440, signal_371}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({signal_2159, signal_2158, signal_2157, signal_610}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_595 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1142, signal_1141, signal_1140, signal_272}), .a ({signal_1313, signal_1312, signal_1311, signal_328}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({signal_2162, signal_2161, signal_2160, signal_611}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_596 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1094, signal_1093, signal_1092, signal_256}), .a ({signal_1517, signal_1516, signal_1515, signal_396}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({signal_2165, signal_2164, signal_2163, signal_612}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_597 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1520, signal_1519, signal_1518, signal_397}), .a ({signal_7493, signal_7491, signal_7489, signal_7487}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({signal_2168, signal_2167, signal_2166, signal_613}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_598 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1220, signal_1219, signal_1218, signal_297}), .a ({signal_1088, signal_1087, signal_1086, signal_254}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_2171, signal_2170, signal_2169, signal_614}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_599 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1397, signal_1396, signal_1395, signal_356}), .a ({signal_1337, signal_1336, signal_1335, signal_336}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({signal_2174, signal_2173, signal_2172, signal_615}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_600 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1244, signal_1243, signal_1242, signal_305}), .a ({signal_1523, signal_1522, signal_1521, signal_398}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({signal_2177, signal_2176, signal_2175, signal_616}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_601 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1526, signal_1525, signal_1524, signal_399}), .a ({signal_1037, signal_1036, signal_1035, signal_237}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({signal_2180, signal_2179, signal_2178, signal_617}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_602 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1529, signal_1528, signal_1527, signal_400}), .a ({1'b0, 1'b0, 1'b0, signal_7485}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({signal_2183, signal_2182, signal_2181, signal_618}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_603 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1130, signal_1129, signal_1128, signal_268}), .a ({signal_1199, signal_1198, signal_1197, signal_290}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_2186, signal_2185, signal_2184, signal_619}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_604 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1532, signal_1531, signal_1530, signal_401}), .a ({signal_1070, signal_1069, signal_1068, signal_248}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({signal_2189, signal_2188, signal_2187, signal_620}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_605 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({1'b0, 1'b0, 1'b0, signal_7443}), .a ({signal_1535, signal_1534, signal_1533, signal_402}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({signal_2192, signal_2191, signal_2190, signal_621}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_606 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1016, signal_1015, signal_1014, signal_230}), .a ({signal_1538, signal_1537, signal_1536, signal_403}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({signal_2195, signal_2194, signal_2193, signal_622}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_607 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1247, signal_1246, signal_1245, signal_306}), .a ({signal_1061, signal_1060, signal_1059, signal_245}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({signal_2198, signal_2197, signal_2196, signal_623}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_608 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1070, signal_1069, signal_1068, signal_248}), .a ({signal_1373, signal_1372, signal_1371, signal_348}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_2201, signal_2200, signal_2199, signal_624}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_609 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1361, signal_1360, signal_1359, signal_344}), .a ({signal_7557, signal_7555, signal_7553, signal_7551}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({signal_2204, signal_2203, signal_2202, signal_625}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_610 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1544, signal_1543, signal_1542, signal_405}), .a ({signal_1109, signal_1108, signal_1107, signal_261}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({signal_2207, signal_2206, signal_2205, signal_626}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_611 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1136, signal_1135, signal_1134, signal_270}), .a ({signal_1442, signal_1441, signal_1440, signal_371}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({signal_2210, signal_2209, signal_2208, signal_627}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_612 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1319, signal_1318, signal_1317, signal_330}), .a ({1'b0, 1'b0, 1'b0, signal_7485}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({signal_2213, signal_2212, signal_2211, signal_628}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_613 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1469, signal_1468, signal_1467, signal_380}), .a ({signal_7565, signal_7563, signal_7561, signal_7559}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_2216, signal_2215, signal_2214, signal_629}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_614 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1547, signal_1546, signal_1545, signal_406}), .a ({signal_1208, signal_1207, signal_1206, signal_293}), .clk ( clk ), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({signal_2219, signal_2218, signal_2217, signal_630}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_615 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1310, signal_1309, signal_1308, signal_327}), .a ({signal_1538, signal_1537, signal_1536, signal_403}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({signal_2222, signal_2221, signal_2220, signal_631}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_616 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1124, signal_1123, signal_1122, signal_266}), .a ({signal_1460, signal_1459, signal_1458, signal_377}), .clk ( clk ), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({signal_2225, signal_2224, signal_2223, signal_632}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_617 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1550, signal_1549, signal_1548, signal_407}), .a ({signal_1130, signal_1129, signal_1128, signal_268}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({signal_2228, signal_2227, signal_2226, signal_633}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_618 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1481, signal_1480, signal_1479, signal_384}), .a ({signal_1136, signal_1135, signal_1134, signal_270}), .clk ( clk ), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_2231, signal_2230, signal_2229, signal_634}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_619 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1211, signal_1210, signal_1209, signal_294}), .a ({signal_1388, signal_1387, signal_1386, signal_353}), .clk ( clk ), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({signal_2234, signal_2233, signal_2232, signal_635}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_620 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1553, signal_1552, signal_1551, signal_408}), .a ({signal_1160, signal_1159, signal_1158, signal_278}), .clk ( clk ), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({signal_2237, signal_2236, signal_2235, signal_636}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_621 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7557, signal_7555, signal_7553, signal_7551}), .a ({signal_1229, signal_1228, signal_1227, signal_300}), .clk ( clk ), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({signal_2240, signal_2239, signal_2238, signal_637}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_622 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1211, signal_1210, signal_1209, signal_294}), .a ({signal_1091, signal_1090, signal_1089, signal_255}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({signal_2243, signal_2242, signal_2241, signal_638}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_623 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1151, signal_1150, signal_1149, signal_275}), .a ({signal_1556, signal_1555, signal_1554, signal_409}), .clk ( clk ), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_2246, signal_2245, signal_2244, signal_639}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_624 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1028, signal_1027, signal_1026, signal_234}), .a ({signal_7483, signal_7481, signal_7479, signal_7477}), .clk ( clk ), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({signal_2249, signal_2248, signal_2247, signal_640}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_625 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1043, signal_1042, signal_1041, signal_239}), .a ({signal_1154, signal_1153, signal_1152, signal_276}), .clk ( clk ), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({signal_2252, signal_2251, signal_2250, signal_641}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_626 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1331, signal_1330, signal_1329, signal_334}), .a ({signal_1457, signal_1456, signal_1455, signal_376}), .clk ( clk ), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({signal_2255, signal_2254, signal_2253, signal_642}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_627 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7509, signal_7507, signal_7505, signal_7503}), .a ({signal_1559, signal_1558, signal_1557, signal_410}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({signal_2258, signal_2257, signal_2256, signal_643}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_628 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1412, signal_1411, signal_1410, signal_361}), .a ({signal_1361, signal_1360, signal_1359, signal_344}), .clk ( clk ), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_2261, signal_2260, signal_2259, signal_644}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_629 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_977, signal_976, signal_975, signal_217}), .a ({signal_1139, signal_1138, signal_1137, signal_271}), .clk ( clk ), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({signal_2264, signal_2263, signal_2262, signal_645}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_630 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1055, signal_1054, signal_1053, signal_243}), .a ({signal_1376, signal_1375, signal_1374, signal_349}), .clk ( clk ), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({signal_2267, signal_2266, signal_2265, signal_646}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_631 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1070, signal_1069, signal_1068, signal_248}), .a ({signal_7433, signal_7431, signal_7429, signal_7427}), .clk ( clk ), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({signal_2270, signal_2269, signal_2268, signal_647}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_632 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1322, signal_1321, signal_1320, signal_331}), .a ({signal_1115, signal_1114, signal_1113, signal_263}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({signal_2273, signal_2272, signal_2271, signal_648}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_633 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1085, signal_1084, signal_1083, signal_253}), .a ({signal_1097, signal_1096, signal_1095, signal_257}), .clk ( clk ), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_2276, signal_2275, signal_2274, signal_649}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_634 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_7467, signal_7465, signal_7463, signal_7461}), .a ({signal_1157, signal_1156, signal_1155, signal_277}), .clk ( clk ), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({signal_2279, signal_2278, signal_2277, signal_650}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_635 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1457, signal_1456, signal_1455, signal_376}), .a ({signal_1226, signal_1225, signal_1224, signal_299}), .clk ( clk ), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({signal_2282, signal_2281, signal_2280, signal_651}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_636 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1439, signal_1438, signal_1437, signal_370}), .a ({signal_1394, signal_1393, signal_1392, signal_355}), .clk ( clk ), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({signal_2285, signal_2284, signal_2283, signal_652}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_637 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1271, signal_1270, signal_1269, signal_314}), .a ({signal_1379, signal_1378, signal_1377, signal_350}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({signal_2288, signal_2287, signal_2286, signal_653}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_638 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1112, signal_1111, signal_1110, signal_262}), .a ({signal_7459, signal_7457, signal_7455, signal_7453}), .clk ( clk ), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_2291, signal_2290, signal_2289, signal_654}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_639 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1160, signal_1159, signal_1158, signal_278}), .a ({signal_1439, signal_1438, signal_1437, signal_370}), .clk ( clk ), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({signal_2294, signal_2293, signal_2292, signal_655}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_640 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1451, signal_1450, signal_1449, signal_374}), .a ({signal_1130, signal_1129, signal_1128, signal_268}), .clk ( clk ), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({signal_2297, signal_2296, signal_2295, signal_656}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_641 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1487, signal_1486, signal_1485, signal_386}), .a ({signal_1277, signal_1276, signal_1275, signal_316}), .clk ( clk ), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({signal_2300, signal_2299, signal_2298, signal_657}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_642 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1202, signal_1201, signal_1200, signal_291}), .a ({signal_1172, signal_1171, signal_1170, signal_281}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({signal_2303, signal_2302, signal_2301, signal_658}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_643 ( .s ({signal_7401, signal_7399, signal_7397, signal_7395}), .b ({signal_1286, signal_1285, signal_1284, signal_319}), .a ({signal_1154, signal_1153, signal_1152, signal_276}), .clk ( clk ), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_2306, signal_2305, signal_2304, signal_659}) ) ;
    buf_clk cell_1089 ( .C ( clk ), .D ( signal_7570 ), .Q ( signal_7571 ) ) ;
    buf_clk cell_1095 ( .C ( clk ), .D ( signal_7576 ), .Q ( signal_7577 ) ) ;
    buf_clk cell_1101 ( .C ( clk ), .D ( signal_7582 ), .Q ( signal_7583 ) ) ;
    buf_clk cell_1107 ( .C ( clk ), .D ( signal_7588 ), .Q ( signal_7589 ) ) ;
    buf_clk cell_1109 ( .C ( clk ), .D ( signal_7590 ), .Q ( signal_7591 ) ) ;
    buf_clk cell_1111 ( .C ( clk ), .D ( signal_7592 ), .Q ( signal_7593 ) ) ;
    buf_clk cell_1113 ( .C ( clk ), .D ( signal_7594 ), .Q ( signal_7595 ) ) ;
    buf_clk cell_1115 ( .C ( clk ), .D ( signal_7596 ), .Q ( signal_7597 ) ) ;
    buf_clk cell_1117 ( .C ( clk ), .D ( signal_7598 ), .Q ( signal_7599 ) ) ;
    buf_clk cell_1119 ( .C ( clk ), .D ( signal_7600 ), .Q ( signal_7601 ) ) ;
    buf_clk cell_1121 ( .C ( clk ), .D ( signal_7602 ), .Q ( signal_7603 ) ) ;
    buf_clk cell_1123 ( .C ( clk ), .D ( signal_7604 ), .Q ( signal_7605 ) ) ;
    buf_clk cell_1129 ( .C ( clk ), .D ( signal_7610 ), .Q ( signal_7611 ) ) ;
    buf_clk cell_1137 ( .C ( clk ), .D ( signal_7618 ), .Q ( signal_7619 ) ) ;
    buf_clk cell_1145 ( .C ( clk ), .D ( signal_7626 ), .Q ( signal_7627 ) ) ;
    buf_clk cell_1153 ( .C ( clk ), .D ( signal_7634 ), .Q ( signal_7635 ) ) ;
    buf_clk cell_1161 ( .C ( clk ), .D ( signal_7642 ), .Q ( signal_7643 ) ) ;
    buf_clk cell_1171 ( .C ( clk ), .D ( signal_7652 ), .Q ( signal_7653 ) ) ;
    buf_clk cell_1181 ( .C ( clk ), .D ( signal_7662 ), .Q ( signal_7663 ) ) ;
    buf_clk cell_1191 ( .C ( clk ), .D ( signal_7672 ), .Q ( signal_7673 ) ) ;
    buf_clk cell_1201 ( .C ( clk ), .D ( signal_7682 ), .Q ( signal_7683 ) ) ;
    buf_clk cell_1213 ( .C ( clk ), .D ( signal_7694 ), .Q ( signal_7695 ) ) ;
    buf_clk cell_1225 ( .C ( clk ), .D ( signal_7706 ), .Q ( signal_7707 ) ) ;
    buf_clk cell_1237 ( .C ( clk ), .D ( signal_7718 ), .Q ( signal_7719 ) ) ;
    buf_clk cell_1249 ( .C ( clk ), .D ( signal_7730 ), .Q ( signal_7731 ) ) ;
    buf_clk cell_1263 ( .C ( clk ), .D ( signal_7744 ), .Q ( signal_7745 ) ) ;
    buf_clk cell_1277 ( .C ( clk ), .D ( signal_7758 ), .Q ( signal_7759 ) ) ;
    buf_clk cell_1291 ( .C ( clk ), .D ( signal_7772 ), .Q ( signal_7773 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_1130 ( .C ( clk ), .D ( signal_7611 ), .Q ( signal_7612 ) ) ;
    buf_clk cell_1138 ( .C ( clk ), .D ( signal_7619 ), .Q ( signal_7620 ) ) ;
    buf_clk cell_1146 ( .C ( clk ), .D ( signal_7627 ), .Q ( signal_7628 ) ) ;
    buf_clk cell_1154 ( .C ( clk ), .D ( signal_7635 ), .Q ( signal_7636 ) ) ;
    buf_clk cell_1162 ( .C ( clk ), .D ( signal_7643 ), .Q ( signal_7644 ) ) ;
    buf_clk cell_1172 ( .C ( clk ), .D ( signal_7653 ), .Q ( signal_7654 ) ) ;
    buf_clk cell_1182 ( .C ( clk ), .D ( signal_7663 ), .Q ( signal_7664 ) ) ;
    buf_clk cell_1192 ( .C ( clk ), .D ( signal_7673 ), .Q ( signal_7674 ) ) ;
    buf_clk cell_1202 ( .C ( clk ), .D ( signal_7683 ), .Q ( signal_7684 ) ) ;
    buf_clk cell_1214 ( .C ( clk ), .D ( signal_7695 ), .Q ( signal_7696 ) ) ;
    buf_clk cell_1226 ( .C ( clk ), .D ( signal_7707 ), .Q ( signal_7708 ) ) ;
    buf_clk cell_1238 ( .C ( clk ), .D ( signal_7719 ), .Q ( signal_7720 ) ) ;
    buf_clk cell_1250 ( .C ( clk ), .D ( signal_7731 ), .Q ( signal_7732 ) ) ;
    buf_clk cell_1264 ( .C ( clk ), .D ( signal_7745 ), .Q ( signal_7746 ) ) ;
    buf_clk cell_1278 ( .C ( clk ), .D ( signal_7759 ), .Q ( signal_7760 ) ) ;
    buf_clk cell_1292 ( .C ( clk ), .D ( signal_7773 ), .Q ( signal_7774 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_644 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1568, signal_1567, signal_1566, signal_413}), .a ({signal_1565, signal_1564, signal_1563, signal_412}), .clk ( clk ), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({signal_2312, signal_2311, signal_2310, signal_660}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_645 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1574, signal_1573, signal_1572, signal_415}), .a ({signal_1571, signal_1570, signal_1569, signal_414}), .clk ( clk ), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({signal_2315, signal_2314, signal_2313, signal_661}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_646 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1580, signal_1579, signal_1578, signal_417}), .a ({signal_1577, signal_1576, signal_1575, signal_416}), .clk ( clk ), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({signal_2318, signal_2317, signal_2316, signal_662}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_647 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1586, signal_1585, signal_1584, signal_419}), .a ({signal_1583, signal_1582, signal_1581, signal_418}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({signal_2321, signal_2320, signal_2319, signal_663}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_648 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1592, signal_1591, signal_1590, signal_421}), .a ({signal_1589, signal_1588, signal_1587, signal_420}), .clk ( clk ), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_2324, signal_2323, signal_2322, signal_664}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_649 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1598, signal_1597, signal_1596, signal_423}), .a ({signal_1595, signal_1594, signal_1593, signal_422}), .clk ( clk ), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({signal_2327, signal_2326, signal_2325, signal_665}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_650 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1604, signal_1603, signal_1602, signal_425}), .a ({signal_1601, signal_1600, signal_1599, signal_424}), .clk ( clk ), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({signal_2330, signal_2329, signal_2328, signal_666}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_651 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1610, signal_1609, signal_1608, signal_427}), .a ({signal_1607, signal_1606, signal_1605, signal_426}), .clk ( clk ), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({signal_2333, signal_2332, signal_2331, signal_667}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_652 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1616, signal_1615, signal_1614, signal_429}), .a ({signal_1613, signal_1612, signal_1611, signal_428}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({signal_2336, signal_2335, signal_2334, signal_668}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_653 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1622, signal_1621, signal_1620, signal_431}), .a ({signal_1619, signal_1618, signal_1617, signal_430}), .clk ( clk ), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_2339, signal_2338, signal_2337, signal_669}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_654 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1628, signal_1627, signal_1626, signal_433}), .a ({signal_1625, signal_1624, signal_1623, signal_432}), .clk ( clk ), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({signal_2342, signal_2341, signal_2340, signal_670}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_655 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1634, signal_1633, signal_1632, signal_435}), .a ({signal_1631, signal_1630, signal_1629, signal_434}), .clk ( clk ), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({signal_2345, signal_2344, signal_2343, signal_671}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_656 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1640, signal_1639, signal_1638, signal_437}), .a ({signal_1637, signal_1636, signal_1635, signal_436}), .clk ( clk ), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({signal_2348, signal_2347, signal_2346, signal_672}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_657 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1646, signal_1645, signal_1644, signal_439}), .a ({signal_1643, signal_1642, signal_1641, signal_438}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({signal_2351, signal_2350, signal_2349, signal_673}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_658 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1652, signal_1651, signal_1650, signal_441}), .a ({signal_1649, signal_1648, signal_1647, signal_440}), .clk ( clk ), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_2354, signal_2353, signal_2352, signal_674}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_659 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1658, signal_1657, signal_1656, signal_443}), .a ({signal_1655, signal_1654, signal_1653, signal_442}), .clk ( clk ), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({signal_2357, signal_2356, signal_2355, signal_675}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_660 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1661, signal_1660, signal_1659, signal_444}), .a ({signal_1169, signal_1168, signal_1167, signal_280}), .clk ( clk ), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({signal_2360, signal_2359, signal_2358, signal_676}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_661 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1667, signal_1666, signal_1665, signal_446}), .a ({signal_1664, signal_1663, signal_1662, signal_445}), .clk ( clk ), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({signal_2363, signal_2362, signal_2361, signal_677}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_662 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1673, signal_1672, signal_1671, signal_448}), .a ({signal_1670, signal_1669, signal_1668, signal_447}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({signal_2366, signal_2365, signal_2364, signal_678}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_663 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1679, signal_1678, signal_1677, signal_450}), .a ({signal_1676, signal_1675, signal_1674, signal_449}), .clk ( clk ), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_2369, signal_2368, signal_2367, signal_679}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_664 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1685, signal_1684, signal_1683, signal_452}), .a ({signal_1682, signal_1681, signal_1680, signal_451}), .clk ( clk ), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({signal_2372, signal_2371, signal_2370, signal_680}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_665 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1691, signal_1690, signal_1689, signal_454}), .a ({signal_1688, signal_1687, signal_1686, signal_453}), .clk ( clk ), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({signal_2375, signal_2374, signal_2373, signal_681}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_666 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1697, signal_1696, signal_1695, signal_456}), .a ({signal_1694, signal_1693, signal_1692, signal_455}), .clk ( clk ), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({signal_2378, signal_2377, signal_2376, signal_682}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_667 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1703, signal_1702, signal_1701, signal_458}), .a ({signal_1700, signal_1699, signal_1698, signal_457}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({signal_2381, signal_2380, signal_2379, signal_683}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_668 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1709, signal_1708, signal_1707, signal_460}), .a ({signal_1706, signal_1705, signal_1704, signal_459}), .clk ( clk ), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_2384, signal_2383, signal_2382, signal_684}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_669 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1715, signal_1714, signal_1713, signal_462}), .a ({signal_1712, signal_1711, signal_1710, signal_461}), .clk ( clk ), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({signal_2387, signal_2386, signal_2385, signal_685}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_670 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1721, signal_1720, signal_1719, signal_464}), .a ({signal_1718, signal_1717, signal_1716, signal_463}), .clk ( clk ), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({signal_2390, signal_2389, signal_2388, signal_686}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_671 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1727, signal_1726, signal_1725, signal_466}), .a ({signal_1724, signal_1723, signal_1722, signal_465}), .clk ( clk ), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({signal_2393, signal_2392, signal_2391, signal_687}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_672 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1733, signal_1732, signal_1731, signal_468}), .a ({signal_1730, signal_1729, signal_1728, signal_467}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({signal_2396, signal_2395, signal_2394, signal_688}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_673 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1739, signal_1738, signal_1737, signal_470}), .a ({signal_1736, signal_1735, signal_1734, signal_469}), .clk ( clk ), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_2399, signal_2398, signal_2397, signal_689}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_674 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1745, signal_1744, signal_1743, signal_472}), .a ({signal_1742, signal_1741, signal_1740, signal_471}), .clk ( clk ), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({signal_2402, signal_2401, signal_2400, signal_690}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_675 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1751, signal_1750, signal_1749, signal_474}), .a ({signal_1748, signal_1747, signal_1746, signal_473}), .clk ( clk ), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({signal_2405, signal_2404, signal_2403, signal_691}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_676 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1757, signal_1756, signal_1755, signal_476}), .a ({signal_1754, signal_1753, signal_1752, signal_475}), .clk ( clk ), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({signal_2408, signal_2407, signal_2406, signal_692}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_677 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1763, signal_1762, signal_1761, signal_478}), .a ({signal_1760, signal_1759, signal_1758, signal_477}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({signal_2411, signal_2410, signal_2409, signal_693}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_678 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1769, signal_1768, signal_1767, signal_480}), .a ({signal_1766, signal_1765, signal_1764, signal_479}), .clk ( clk ), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_2414, signal_2413, signal_2412, signal_694}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_679 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1775, signal_1774, signal_1773, signal_482}), .a ({signal_1772, signal_1771, signal_1770, signal_481}), .clk ( clk ), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({signal_2417, signal_2416, signal_2415, signal_695}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_680 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1781, signal_1780, signal_1779, signal_484}), .a ({signal_1778, signal_1777, signal_1776, signal_483}), .clk ( clk ), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({signal_2420, signal_2419, signal_2418, signal_696}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_681 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1787, signal_1786, signal_1785, signal_486}), .a ({signal_1784, signal_1783, signal_1782, signal_485}), .clk ( clk ), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({signal_2423, signal_2422, signal_2421, signal_697}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_682 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1793, signal_1792, signal_1791, signal_488}), .a ({signal_1790, signal_1789, signal_1788, signal_487}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({signal_2426, signal_2425, signal_2424, signal_698}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_683 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1799, signal_1798, signal_1797, signal_490}), .a ({signal_1796, signal_1795, signal_1794, signal_489}), .clk ( clk ), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_2429, signal_2428, signal_2427, signal_699}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_684 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1805, signal_1804, signal_1803, signal_492}), .a ({signal_1802, signal_1801, signal_1800, signal_491}), .clk ( clk ), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({signal_2432, signal_2431, signal_2430, signal_700}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_685 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1811, signal_1810, signal_1809, signal_494}), .a ({signal_1808, signal_1807, signal_1806, signal_493}), .clk ( clk ), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({signal_2435, signal_2434, signal_2433, signal_701}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_686 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1817, signal_1816, signal_1815, signal_496}), .a ({signal_1814, signal_1813, signal_1812, signal_495}), .clk ( clk ), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({signal_2438, signal_2437, signal_2436, signal_702}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_687 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1823, signal_1822, signal_1821, signal_498}), .a ({signal_1820, signal_1819, signal_1818, signal_497}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({signal_2441, signal_2440, signal_2439, signal_703}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_688 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1829, signal_1828, signal_1827, signal_500}), .a ({signal_1826, signal_1825, signal_1824, signal_499}), .clk ( clk ), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_2444, signal_2443, signal_2442, signal_704}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_689 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1832, signal_1831, signal_1830, signal_501}), .a ({signal_1343, signal_1342, signal_1341, signal_338}), .clk ( clk ), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({signal_2447, signal_2446, signal_2445, signal_705}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_690 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1835, signal_1834, signal_1833, signal_502}), .a ({signal_1352, signal_1351, signal_1350, signal_341}), .clk ( clk ), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({signal_2450, signal_2449, signal_2448, signal_706}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_691 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1841, signal_1840, signal_1839, signal_504}), .a ({signal_1838, signal_1837, signal_1836, signal_503}), .clk ( clk ), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({signal_2453, signal_2452, signal_2451, signal_707}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_692 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1847, signal_1846, signal_1845, signal_506}), .a ({signal_1844, signal_1843, signal_1842, signal_505}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({signal_2456, signal_2455, signal_2454, signal_708}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_693 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1853, signal_1852, signal_1851, signal_508}), .a ({signal_1850, signal_1849, signal_1848, signal_507}), .clk ( clk ), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_2459, signal_2458, signal_2457, signal_709}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_694 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1859, signal_1858, signal_1857, signal_510}), .a ({signal_1856, signal_1855, signal_1854, signal_509}), .clk ( clk ), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({signal_2462, signal_2461, signal_2460, signal_710}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_695 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1862, signal_1861, signal_1860, signal_511}), .a ({signal_1364, signal_1363, signal_1362, signal_345}), .clk ( clk ), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({signal_2465, signal_2464, signal_2463, signal_711}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_696 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1868, signal_1867, signal_1866, signal_513}), .a ({signal_1865, signal_1864, signal_1863, signal_512}), .clk ( clk ), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({signal_2468, signal_2467, signal_2466, signal_712}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_697 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1874, signal_1873, signal_1872, signal_515}), .a ({signal_1871, signal_1870, signal_1869, signal_514}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({signal_2471, signal_2470, signal_2469, signal_713}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_698 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1880, signal_1879, signal_1878, signal_517}), .a ({signal_1877, signal_1876, signal_1875, signal_516}), .clk ( clk ), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_2474, signal_2473, signal_2472, signal_714}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_699 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1886, signal_1885, signal_1884, signal_519}), .a ({signal_1883, signal_1882, signal_1881, signal_518}), .clk ( clk ), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({signal_2477, signal_2476, signal_2475, signal_715}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_700 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1892, signal_1891, signal_1890, signal_521}), .a ({signal_1889, signal_1888, signal_1887, signal_520}), .clk ( clk ), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({signal_2480, signal_2479, signal_2478, signal_716}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_701 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1898, signal_1897, signal_1896, signal_523}), .a ({signal_1895, signal_1894, signal_1893, signal_522}), .clk ( clk ), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({signal_2483, signal_2482, signal_2481, signal_717}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_702 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1904, signal_1903, signal_1902, signal_525}), .a ({signal_1901, signal_1900, signal_1899, signal_524}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({signal_2486, signal_2485, signal_2484, signal_718}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_703 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1910, signal_1909, signal_1908, signal_527}), .a ({signal_1907, signal_1906, signal_1905, signal_526}), .clk ( clk ), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_2489, signal_2488, signal_2487, signal_719}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_704 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1916, signal_1915, signal_1914, signal_529}), .a ({signal_1913, signal_1912, signal_1911, signal_528}), .clk ( clk ), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({signal_2492, signal_2491, signal_2490, signal_720}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_705 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1922, signal_1921, signal_1920, signal_531}), .a ({signal_1919, signal_1918, signal_1917, signal_530}), .clk ( clk ), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({signal_2495, signal_2494, signal_2493, signal_721}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_706 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1928, signal_1927, signal_1926, signal_533}), .a ({signal_1925, signal_1924, signal_1923, signal_532}), .clk ( clk ), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({signal_2498, signal_2497, signal_2496, signal_722}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_707 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1934, signal_1933, signal_1932, signal_535}), .a ({signal_1931, signal_1930, signal_1929, signal_534}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({signal_2501, signal_2500, signal_2499, signal_723}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_708 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1940, signal_1939, signal_1938, signal_537}), .a ({signal_1937, signal_1936, signal_1935, signal_536}), .clk ( clk ), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_2504, signal_2503, signal_2502, signal_724}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_709 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1946, signal_1945, signal_1944, signal_539}), .a ({signal_1943, signal_1942, signal_1941, signal_538}), .clk ( clk ), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({signal_2507, signal_2506, signal_2505, signal_725}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_710 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1952, signal_1951, signal_1950, signal_541}), .a ({signal_1949, signal_1948, signal_1947, signal_540}), .clk ( clk ), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({signal_2510, signal_2509, signal_2508, signal_726}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_711 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1958, signal_1957, signal_1956, signal_543}), .a ({signal_1955, signal_1954, signal_1953, signal_542}), .clk ( clk ), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({signal_2513, signal_2512, signal_2511, signal_727}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_712 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1964, signal_1963, signal_1962, signal_545}), .a ({signal_1961, signal_1960, signal_1959, signal_544}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({signal_2516, signal_2515, signal_2514, signal_728}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_713 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1970, signal_1969, signal_1968, signal_547}), .a ({signal_1967, signal_1966, signal_1965, signal_546}), .clk ( clk ), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_2519, signal_2518, signal_2517, signal_729}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_714 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1976, signal_1975, signal_1974, signal_549}), .a ({signal_1973, signal_1972, signal_1971, signal_548}), .clk ( clk ), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({signal_2522, signal_2521, signal_2520, signal_730}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_715 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1982, signal_1981, signal_1980, signal_551}), .a ({signal_1979, signal_1978, signal_1977, signal_550}), .clk ( clk ), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({signal_2525, signal_2524, signal_2523, signal_731}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_716 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1988, signal_1987, signal_1986, signal_553}), .a ({signal_1985, signal_1984, signal_1983, signal_552}), .clk ( clk ), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({signal_2528, signal_2527, signal_2526, signal_732}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_717 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1994, signal_1993, signal_1992, signal_555}), .a ({signal_1991, signal_1990, signal_1989, signal_554}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({signal_2531, signal_2530, signal_2529, signal_733}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_718 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2000, signal_1999, signal_1998, signal_557}), .a ({signal_1997, signal_1996, signal_1995, signal_556}), .clk ( clk ), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_2534, signal_2533, signal_2532, signal_734}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_719 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2006, signal_2005, signal_2004, signal_559}), .a ({signal_2003, signal_2002, signal_2001, signal_558}), .clk ( clk ), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({signal_2537, signal_2536, signal_2535, signal_735}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_720 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2012, signal_2011, signal_2010, signal_561}), .a ({signal_2009, signal_2008, signal_2007, signal_560}), .clk ( clk ), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({signal_2540, signal_2539, signal_2538, signal_736}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_721 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2018, signal_2017, signal_2016, signal_563}), .a ({signal_2015, signal_2014, signal_2013, signal_562}), .clk ( clk ), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({signal_2543, signal_2542, signal_2541, signal_737}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_722 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2024, signal_2023, signal_2022, signal_565}), .a ({signal_2021, signal_2020, signal_2019, signal_564}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({signal_2546, signal_2545, signal_2544, signal_738}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_723 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2030, signal_2029, signal_2028, signal_567}), .a ({signal_2027, signal_2026, signal_2025, signal_566}), .clk ( clk ), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_2549, signal_2548, signal_2547, signal_739}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_724 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2036, signal_2035, signal_2034, signal_569}), .a ({signal_2033, signal_2032, signal_2031, signal_568}), .clk ( clk ), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({signal_2552, signal_2551, signal_2550, signal_740}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_725 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2042, signal_2041, signal_2040, signal_571}), .a ({signal_2039, signal_2038, signal_2037, signal_570}), .clk ( clk ), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({signal_2555, signal_2554, signal_2553, signal_741}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_726 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2048, signal_2047, signal_2046, signal_573}), .a ({signal_2045, signal_2044, signal_2043, signal_572}), .clk ( clk ), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({signal_2558, signal_2557, signal_2556, signal_742}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_727 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2054, signal_2053, signal_2052, signal_575}), .a ({signal_2051, signal_2050, signal_2049, signal_574}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({signal_2561, signal_2560, signal_2559, signal_743}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_728 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2060, signal_2059, signal_2058, signal_577}), .a ({signal_2057, signal_2056, signal_2055, signal_576}), .clk ( clk ), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_2564, signal_2563, signal_2562, signal_744}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_729 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2066, signal_2065, signal_2064, signal_579}), .a ({signal_2063, signal_2062, signal_2061, signal_578}), .clk ( clk ), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({signal_2567, signal_2566, signal_2565, signal_745}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_730 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2072, signal_2071, signal_2070, signal_581}), .a ({signal_2069, signal_2068, signal_2067, signal_580}), .clk ( clk ), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({signal_2570, signal_2569, signal_2568, signal_746}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_731 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2078, signal_2077, signal_2076, signal_583}), .a ({signal_2075, signal_2074, signal_2073, signal_582}), .clk ( clk ), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({signal_2573, signal_2572, signal_2571, signal_747}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_732 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2084, signal_2083, signal_2082, signal_585}), .a ({signal_2081, signal_2080, signal_2079, signal_584}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({signal_2576, signal_2575, signal_2574, signal_748}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_733 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1640, signal_1639, signal_1638, signal_437}), .a ({signal_7597, signal_7595, signal_7593, signal_7591}), .clk ( clk ), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_2579, signal_2578, signal_2577, signal_749}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_734 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2090, signal_2089, signal_2088, signal_587}), .a ({signal_2087, signal_2086, signal_2085, signal_586}), .clk ( clk ), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({signal_2582, signal_2581, signal_2580, signal_750}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_735 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2096, signal_2095, signal_2094, signal_589}), .a ({signal_2093, signal_2092, signal_2091, signal_588}), .clk ( clk ), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({signal_2585, signal_2584, signal_2583, signal_751}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_736 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2102, signal_2101, signal_2100, signal_591}), .a ({signal_2099, signal_2098, signal_2097, signal_590}), .clk ( clk ), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({signal_2588, signal_2587, signal_2586, signal_752}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_737 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2108, signal_2107, signal_2106, signal_593}), .a ({signal_2105, signal_2104, signal_2103, signal_592}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({signal_2591, signal_2590, signal_2589, signal_753}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_738 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2114, signal_2113, signal_2112, signal_595}), .a ({signal_2111, signal_2110, signal_2109, signal_594}), .clk ( clk ), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_2594, signal_2593, signal_2592, signal_754}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_739 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2120, signal_2119, signal_2118, signal_597}), .a ({signal_2117, signal_2116, signal_2115, signal_596}), .clk ( clk ), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({signal_2597, signal_2596, signal_2595, signal_755}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_740 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2126, signal_2125, signal_2124, signal_599}), .a ({signal_2123, signal_2122, signal_2121, signal_598}), .clk ( clk ), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({signal_2600, signal_2599, signal_2598, signal_756}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_741 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2132, signal_2131, signal_2130, signal_601}), .a ({signal_2129, signal_2128, signal_2127, signal_600}), .clk ( clk ), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({signal_2603, signal_2602, signal_2601, signal_757}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_742 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2138, signal_2137, signal_2136, signal_603}), .a ({signal_2135, signal_2134, signal_2133, signal_602}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({signal_2606, signal_2605, signal_2604, signal_758}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_743 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2144, signal_2143, signal_2142, signal_605}), .a ({signal_2141, signal_2140, signal_2139, signal_604}), .clk ( clk ), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_2609, signal_2608, signal_2607, signal_759}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_744 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2150, signal_2149, signal_2148, signal_607}), .a ({signal_2147, signal_2146, signal_2145, signal_606}), .clk ( clk ), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({signal_2612, signal_2611, signal_2610, signal_760}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_745 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2156, signal_2155, signal_2154, signal_609}), .a ({signal_2153, signal_2152, signal_2151, signal_608}), .clk ( clk ), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({signal_2615, signal_2614, signal_2613, signal_761}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_746 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2162, signal_2161, signal_2160, signal_611}), .a ({signal_2159, signal_2158, signal_2157, signal_610}), .clk ( clk ), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({signal_2618, signal_2617, signal_2616, signal_762}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_747 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2168, signal_2167, signal_2166, signal_613}), .a ({signal_2165, signal_2164, signal_2163, signal_612}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({signal_2621, signal_2620, signal_2619, signal_763}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_748 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2174, signal_2173, signal_2172, signal_615}), .a ({signal_2171, signal_2170, signal_2169, signal_614}), .clk ( clk ), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_2624, signal_2623, signal_2622, signal_764}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_749 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2180, signal_2179, signal_2178, signal_617}), .a ({signal_2177, signal_2176, signal_2175, signal_616}), .clk ( clk ), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({signal_2627, signal_2626, signal_2625, signal_765}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_750 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2186, signal_2185, signal_2184, signal_619}), .a ({signal_2183, signal_2182, signal_2181, signal_618}), .clk ( clk ), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({signal_2630, signal_2629, signal_2628, signal_766}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_751 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2192, signal_2191, signal_2190, signal_621}), .a ({signal_2189, signal_2188, signal_2187, signal_620}), .clk ( clk ), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({signal_2633, signal_2632, signal_2631, signal_767}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_752 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2198, signal_2197, signal_2196, signal_623}), .a ({signal_2195, signal_2194, signal_2193, signal_622}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({signal_2636, signal_2635, signal_2634, signal_768}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_753 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2201, signal_2200, signal_2199, signal_624}), .a ({signal_7605, signal_7603, signal_7601, signal_7599}), .clk ( clk ), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_2639, signal_2638, signal_2637, signal_769}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_754 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2207, signal_2206, signal_2205, signal_626}), .a ({signal_2204, signal_2203, signal_2202, signal_625}), .clk ( clk ), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({signal_2642, signal_2641, signal_2640, signal_770}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_755 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2213, signal_2212, signal_2211, signal_628}), .a ({signal_2210, signal_2209, signal_2208, signal_627}), .clk ( clk ), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({signal_2645, signal_2644, signal_2643, signal_771}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_756 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2219, signal_2218, signal_2217, signal_630}), .a ({signal_2216, signal_2215, signal_2214, signal_629}), .clk ( clk ), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({signal_2648, signal_2647, signal_2646, signal_772}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_757 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2225, signal_2224, signal_2223, signal_632}), .a ({signal_2222, signal_2221, signal_2220, signal_631}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({signal_2651, signal_2650, signal_2649, signal_773}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_758 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2231, signal_2230, signal_2229, signal_634}), .a ({signal_2228, signal_2227, signal_2226, signal_633}), .clk ( clk ), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_2654, signal_2653, signal_2652, signal_774}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_759 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2237, signal_2236, signal_2235, signal_636}), .a ({signal_2234, signal_2233, signal_2232, signal_635}), .clk ( clk ), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({signal_2657, signal_2656, signal_2655, signal_775}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_760 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2243, signal_2242, signal_2241, signal_638}), .a ({signal_2240, signal_2239, signal_2238, signal_637}), .clk ( clk ), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({signal_2660, signal_2659, signal_2658, signal_776}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_761 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2249, signal_2248, signal_2247, signal_640}), .a ({signal_2246, signal_2245, signal_2244, signal_639}), .clk ( clk ), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({signal_2663, signal_2662, signal_2661, signal_777}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_762 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2255, signal_2254, signal_2253, signal_642}), .a ({signal_2252, signal_2251, signal_2250, signal_641}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({signal_2666, signal_2665, signal_2664, signal_778}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_763 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2261, signal_2260, signal_2259, signal_644}), .a ({signal_2258, signal_2257, signal_2256, signal_643}), .clk ( clk ), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_2669, signal_2668, signal_2667, signal_779}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_764 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2267, signal_2266, signal_2265, signal_646}), .a ({signal_2264, signal_2263, signal_2262, signal_645}), .clk ( clk ), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({signal_2672, signal_2671, signal_2670, signal_780}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_765 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2273, signal_2272, signal_2271, signal_648}), .a ({signal_2270, signal_2269, signal_2268, signal_647}), .clk ( clk ), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({signal_2675, signal_2674, signal_2673, signal_781}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_766 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2279, signal_2278, signal_2277, signal_650}), .a ({signal_2276, signal_2275, signal_2274, signal_649}), .clk ( clk ), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({signal_2678, signal_2677, signal_2676, signal_782}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_767 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2285, signal_2284, signal_2283, signal_652}), .a ({signal_2282, signal_2281, signal_2280, signal_651}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({signal_2681, signal_2680, signal_2679, signal_783}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_768 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2291, signal_2290, signal_2289, signal_654}), .a ({signal_2288, signal_2287, signal_2286, signal_653}), .clk ( clk ), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_2684, signal_2683, signal_2682, signal_784}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_769 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_1562, signal_1561, signal_1560, signal_411}), .a ({signal_2294, signal_2293, signal_2292, signal_655}), .clk ( clk ), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({signal_2687, signal_2686, signal_2685, signal_785}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_770 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2300, signal_2299, signal_2298, signal_657}), .a ({signal_2297, signal_2296, signal_2295, signal_656}), .clk ( clk ), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({signal_2690, signal_2689, signal_2688, signal_786}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_771 ( .s ({signal_7589, signal_7583, signal_7577, signal_7571}), .b ({signal_2306, signal_2305, signal_2304, signal_659}), .a ({signal_2303, signal_2302, signal_2301, signal_658}), .clk ( clk ), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({signal_2693, signal_2692, signal_2691, signal_787}) ) ;
    buf_clk cell_1131 ( .C ( clk ), .D ( signal_7612 ), .Q ( signal_7613 ) ) ;
    buf_clk cell_1139 ( .C ( clk ), .D ( signal_7620 ), .Q ( signal_7621 ) ) ;
    buf_clk cell_1147 ( .C ( clk ), .D ( signal_7628 ), .Q ( signal_7629 ) ) ;
    buf_clk cell_1155 ( .C ( clk ), .D ( signal_7636 ), .Q ( signal_7637 ) ) ;
    buf_clk cell_1163 ( .C ( clk ), .D ( signal_7644 ), .Q ( signal_7645 ) ) ;
    buf_clk cell_1173 ( .C ( clk ), .D ( signal_7654 ), .Q ( signal_7655 ) ) ;
    buf_clk cell_1183 ( .C ( clk ), .D ( signal_7664 ), .Q ( signal_7665 ) ) ;
    buf_clk cell_1193 ( .C ( clk ), .D ( signal_7674 ), .Q ( signal_7675 ) ) ;
    buf_clk cell_1203 ( .C ( clk ), .D ( signal_7684 ), .Q ( signal_7685 ) ) ;
    buf_clk cell_1215 ( .C ( clk ), .D ( signal_7696 ), .Q ( signal_7697 ) ) ;
    buf_clk cell_1227 ( .C ( clk ), .D ( signal_7708 ), .Q ( signal_7709 ) ) ;
    buf_clk cell_1239 ( .C ( clk ), .D ( signal_7720 ), .Q ( signal_7721 ) ) ;
    buf_clk cell_1251 ( .C ( clk ), .D ( signal_7732 ), .Q ( signal_7733 ) ) ;
    buf_clk cell_1265 ( .C ( clk ), .D ( signal_7746 ), .Q ( signal_7747 ) ) ;
    buf_clk cell_1279 ( .C ( clk ), .D ( signal_7760 ), .Q ( signal_7761 ) ) ;
    buf_clk cell_1293 ( .C ( clk ), .D ( signal_7774 ), .Q ( signal_7775 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_1164 ( .C ( clk ), .D ( signal_7645 ), .Q ( signal_7646 ) ) ;
    buf_clk cell_1174 ( .C ( clk ), .D ( signal_7655 ), .Q ( signal_7656 ) ) ;
    buf_clk cell_1184 ( .C ( clk ), .D ( signal_7665 ), .Q ( signal_7666 ) ) ;
    buf_clk cell_1194 ( .C ( clk ), .D ( signal_7675 ), .Q ( signal_7676 ) ) ;
    buf_clk cell_1204 ( .C ( clk ), .D ( signal_7685 ), .Q ( signal_7686 ) ) ;
    buf_clk cell_1216 ( .C ( clk ), .D ( signal_7697 ), .Q ( signal_7698 ) ) ;
    buf_clk cell_1228 ( .C ( clk ), .D ( signal_7709 ), .Q ( signal_7710 ) ) ;
    buf_clk cell_1240 ( .C ( clk ), .D ( signal_7721 ), .Q ( signal_7722 ) ) ;
    buf_clk cell_1252 ( .C ( clk ), .D ( signal_7733 ), .Q ( signal_7734 ) ) ;
    buf_clk cell_1266 ( .C ( clk ), .D ( signal_7747 ), .Q ( signal_7748 ) ) ;
    buf_clk cell_1280 ( .C ( clk ), .D ( signal_7761 ), .Q ( signal_7762 ) ) ;
    buf_clk cell_1294 ( .C ( clk ), .D ( signal_7775 ), .Q ( signal_7776 ) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_772 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2315, signal_2314, signal_2313, signal_661}), .a ({signal_2312, signal_2311, signal_2310, signal_660}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({signal_2699, signal_2698, signal_2697, signal_788}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_773 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2321, signal_2320, signal_2319, signal_663}), .a ({signal_2318, signal_2317, signal_2316, signal_662}), .clk ( clk ), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_2702, signal_2701, signal_2700, signal_789}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_774 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2327, signal_2326, signal_2325, signal_665}), .a ({signal_2324, signal_2323, signal_2322, signal_664}), .clk ( clk ), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({signal_2705, signal_2704, signal_2703, signal_790}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_775 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2333, signal_2332, signal_2331, signal_667}), .a ({signal_2330, signal_2329, signal_2328, signal_666}), .clk ( clk ), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({signal_2708, signal_2707, signal_2706, signal_791}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_776 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2339, signal_2338, signal_2337, signal_669}), .a ({signal_2336, signal_2335, signal_2334, signal_668}), .clk ( clk ), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({signal_2711, signal_2710, signal_2709, signal_792}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_777 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2345, signal_2344, signal_2343, signal_671}), .a ({signal_2342, signal_2341, signal_2340, signal_670}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({signal_2714, signal_2713, signal_2712, signal_793}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_778 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2351, signal_2350, signal_2349, signal_673}), .a ({signal_2348, signal_2347, signal_2346, signal_672}), .clk ( clk ), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_2717, signal_2716, signal_2715, signal_794}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_779 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2357, signal_2356, signal_2355, signal_675}), .a ({signal_2354, signal_2353, signal_2352, signal_674}), .clk ( clk ), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({signal_2720, signal_2719, signal_2718, signal_795}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_780 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2363, signal_2362, signal_2361, signal_677}), .a ({signal_2360, signal_2359, signal_2358, signal_676}), .clk ( clk ), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({signal_2723, signal_2722, signal_2721, signal_796}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_781 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2369, signal_2368, signal_2367, signal_679}), .a ({signal_2366, signal_2365, signal_2364, signal_678}), .clk ( clk ), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({signal_2726, signal_2725, signal_2724, signal_797}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_782 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2375, signal_2374, signal_2373, signal_681}), .a ({signal_2372, signal_2371, signal_2370, signal_680}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({signal_2729, signal_2728, signal_2727, signal_798}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_783 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2381, signal_2380, signal_2379, signal_683}), .a ({signal_2378, signal_2377, signal_2376, signal_682}), .clk ( clk ), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_2732, signal_2731, signal_2730, signal_799}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_784 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2387, signal_2386, signal_2385, signal_685}), .a ({signal_2384, signal_2383, signal_2382, signal_684}), .clk ( clk ), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({signal_2735, signal_2734, signal_2733, signal_800}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_785 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2393, signal_2392, signal_2391, signal_687}), .a ({signal_2390, signal_2389, signal_2388, signal_686}), .clk ( clk ), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({signal_2738, signal_2737, signal_2736, signal_801}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_786 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2399, signal_2398, signal_2397, signal_689}), .a ({signal_2396, signal_2395, signal_2394, signal_688}), .clk ( clk ), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({signal_2741, signal_2740, signal_2739, signal_802}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_787 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2405, signal_2404, signal_2403, signal_691}), .a ({signal_2402, signal_2401, signal_2400, signal_690}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({signal_2744, signal_2743, signal_2742, signal_803}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_788 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2411, signal_2410, signal_2409, signal_693}), .a ({signal_2408, signal_2407, signal_2406, signal_692}), .clk ( clk ), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_2747, signal_2746, signal_2745, signal_804}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_789 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2417, signal_2416, signal_2415, signal_695}), .a ({signal_2414, signal_2413, signal_2412, signal_694}), .clk ( clk ), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({signal_2750, signal_2749, signal_2748, signal_805}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_790 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2423, signal_2422, signal_2421, signal_697}), .a ({signal_2420, signal_2419, signal_2418, signal_696}), .clk ( clk ), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({signal_2753, signal_2752, signal_2751, signal_806}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_791 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2429, signal_2428, signal_2427, signal_699}), .a ({signal_2426, signal_2425, signal_2424, signal_698}), .clk ( clk ), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({signal_2756, signal_2755, signal_2754, signal_807}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_792 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2435, signal_2434, signal_2433, signal_701}), .a ({signal_2432, signal_2431, signal_2430, signal_700}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({signal_2759, signal_2758, signal_2757, signal_808}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_793 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2441, signal_2440, signal_2439, signal_703}), .a ({signal_2438, signal_2437, signal_2436, signal_702}), .clk ( clk ), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_2762, signal_2761, signal_2760, signal_809}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_794 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2447, signal_2446, signal_2445, signal_705}), .a ({signal_2444, signal_2443, signal_2442, signal_704}), .clk ( clk ), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({signal_2765, signal_2764, signal_2763, signal_810}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_795 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2453, signal_2452, signal_2451, signal_707}), .a ({signal_2450, signal_2449, signal_2448, signal_706}), .clk ( clk ), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({signal_2768, signal_2767, signal_2766, signal_811}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_796 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2459, signal_2458, signal_2457, signal_709}), .a ({signal_2456, signal_2455, signal_2454, signal_708}), .clk ( clk ), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({signal_2771, signal_2770, signal_2769, signal_812}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_797 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2465, signal_2464, signal_2463, signal_711}), .a ({signal_2462, signal_2461, signal_2460, signal_710}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({signal_2774, signal_2773, signal_2772, signal_813}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_798 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2471, signal_2470, signal_2469, signal_713}), .a ({signal_2468, signal_2467, signal_2466, signal_712}), .clk ( clk ), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_2777, signal_2776, signal_2775, signal_814}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_799 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2477, signal_2476, signal_2475, signal_715}), .a ({signal_2474, signal_2473, signal_2472, signal_714}), .clk ( clk ), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({signal_2780, signal_2779, signal_2778, signal_815}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_800 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2483, signal_2482, signal_2481, signal_717}), .a ({signal_2480, signal_2479, signal_2478, signal_716}), .clk ( clk ), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({signal_2783, signal_2782, signal_2781, signal_816}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_801 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2489, signal_2488, signal_2487, signal_719}), .a ({signal_2486, signal_2485, signal_2484, signal_718}), .clk ( clk ), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({signal_2786, signal_2785, signal_2784, signal_817}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_802 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2495, signal_2494, signal_2493, signal_721}), .a ({signal_2492, signal_2491, signal_2490, signal_720}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({signal_2789, signal_2788, signal_2787, signal_818}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_803 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2501, signal_2500, signal_2499, signal_723}), .a ({signal_2498, signal_2497, signal_2496, signal_722}), .clk ( clk ), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_2792, signal_2791, signal_2790, signal_819}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_804 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2507, signal_2506, signal_2505, signal_725}), .a ({signal_2504, signal_2503, signal_2502, signal_724}), .clk ( clk ), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({signal_2795, signal_2794, signal_2793, signal_820}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_805 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2513, signal_2512, signal_2511, signal_727}), .a ({signal_2510, signal_2509, signal_2508, signal_726}), .clk ( clk ), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({signal_2798, signal_2797, signal_2796, signal_821}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_806 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2519, signal_2518, signal_2517, signal_729}), .a ({signal_2516, signal_2515, signal_2514, signal_728}), .clk ( clk ), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({signal_2801, signal_2800, signal_2799, signal_822}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_807 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2525, signal_2524, signal_2523, signal_731}), .a ({signal_2522, signal_2521, signal_2520, signal_730}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({signal_2804, signal_2803, signal_2802, signal_823}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_808 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2531, signal_2530, signal_2529, signal_733}), .a ({signal_2528, signal_2527, signal_2526, signal_732}), .clk ( clk ), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_2807, signal_2806, signal_2805, signal_824}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_809 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2537, signal_2536, signal_2535, signal_735}), .a ({signal_2534, signal_2533, signal_2532, signal_734}), .clk ( clk ), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({signal_2810, signal_2809, signal_2808, signal_825}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_810 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2543, signal_2542, signal_2541, signal_737}), .a ({signal_2540, signal_2539, signal_2538, signal_736}), .clk ( clk ), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({signal_2813, signal_2812, signal_2811, signal_826}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_811 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2549, signal_2548, signal_2547, signal_739}), .a ({signal_2546, signal_2545, signal_2544, signal_738}), .clk ( clk ), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({signal_2816, signal_2815, signal_2814, signal_827}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_812 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2555, signal_2554, signal_2553, signal_741}), .a ({signal_2552, signal_2551, signal_2550, signal_740}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({signal_2819, signal_2818, signal_2817, signal_828}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_813 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2561, signal_2560, signal_2559, signal_743}), .a ({signal_2558, signal_2557, signal_2556, signal_742}), .clk ( clk ), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_2822, signal_2821, signal_2820, signal_829}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_814 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2567, signal_2566, signal_2565, signal_745}), .a ({signal_2564, signal_2563, signal_2562, signal_744}), .clk ( clk ), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({signal_2825, signal_2824, signal_2823, signal_830}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_815 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2573, signal_2572, signal_2571, signal_747}), .a ({signal_2570, signal_2569, signal_2568, signal_746}), .clk ( clk ), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({signal_2828, signal_2827, signal_2826, signal_831}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_816 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2579, signal_2578, signal_2577, signal_749}), .a ({signal_2576, signal_2575, signal_2574, signal_748}), .clk ( clk ), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({signal_2831, signal_2830, signal_2829, signal_832}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_817 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2585, signal_2584, signal_2583, signal_751}), .a ({signal_2582, signal_2581, signal_2580, signal_750}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({signal_2834, signal_2833, signal_2832, signal_833}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_818 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2591, signal_2590, signal_2589, signal_753}), .a ({signal_2588, signal_2587, signal_2586, signal_752}), .clk ( clk ), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_2837, signal_2836, signal_2835, signal_834}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_819 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2597, signal_2596, signal_2595, signal_755}), .a ({signal_2594, signal_2593, signal_2592, signal_754}), .clk ( clk ), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({signal_2840, signal_2839, signal_2838, signal_835}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_820 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2603, signal_2602, signal_2601, signal_757}), .a ({signal_2600, signal_2599, signal_2598, signal_756}), .clk ( clk ), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({signal_2843, signal_2842, signal_2841, signal_836}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_821 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2609, signal_2608, signal_2607, signal_759}), .a ({signal_2606, signal_2605, signal_2604, signal_758}), .clk ( clk ), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({signal_2846, signal_2845, signal_2844, signal_837}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_822 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2615, signal_2614, signal_2613, signal_761}), .a ({signal_2612, signal_2611, signal_2610, signal_760}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({signal_2849, signal_2848, signal_2847, signal_838}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_823 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2621, signal_2620, signal_2619, signal_763}), .a ({signal_2618, signal_2617, signal_2616, signal_762}), .clk ( clk ), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_2852, signal_2851, signal_2850, signal_839}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_824 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2627, signal_2626, signal_2625, signal_765}), .a ({signal_2624, signal_2623, signal_2622, signal_764}), .clk ( clk ), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({signal_2855, signal_2854, signal_2853, signal_840}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_825 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2633, signal_2632, signal_2631, signal_767}), .a ({signal_2630, signal_2629, signal_2628, signal_766}), .clk ( clk ), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({signal_2858, signal_2857, signal_2856, signal_841}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_826 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2639, signal_2638, signal_2637, signal_769}), .a ({signal_2636, signal_2635, signal_2634, signal_768}), .clk ( clk ), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({signal_2861, signal_2860, signal_2859, signal_842}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_827 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2645, signal_2644, signal_2643, signal_771}), .a ({signal_2642, signal_2641, signal_2640, signal_770}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({signal_2864, signal_2863, signal_2862, signal_843}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_828 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2651, signal_2650, signal_2649, signal_773}), .a ({signal_2648, signal_2647, signal_2646, signal_772}), .clk ( clk ), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_2867, signal_2866, signal_2865, signal_844}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_829 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2657, signal_2656, signal_2655, signal_775}), .a ({signal_2654, signal_2653, signal_2652, signal_774}), .clk ( clk ), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({signal_2870, signal_2869, signal_2868, signal_845}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_830 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2663, signal_2662, signal_2661, signal_777}), .a ({signal_2660, signal_2659, signal_2658, signal_776}), .clk ( clk ), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({signal_2873, signal_2872, signal_2871, signal_846}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_831 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2669, signal_2668, signal_2667, signal_779}), .a ({signal_2666, signal_2665, signal_2664, signal_778}), .clk ( clk ), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({signal_2876, signal_2875, signal_2874, signal_847}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_832 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2675, signal_2674, signal_2673, signal_781}), .a ({signal_2672, signal_2671, signal_2670, signal_780}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({signal_2879, signal_2878, signal_2877, signal_848}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_833 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2681, signal_2680, signal_2679, signal_783}), .a ({signal_2678, signal_2677, signal_2676, signal_782}), .clk ( clk ), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_2882, signal_2881, signal_2880, signal_849}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_834 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2687, signal_2686, signal_2685, signal_785}), .a ({signal_2684, signal_2683, signal_2682, signal_784}), .clk ( clk ), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({signal_2885, signal_2884, signal_2883, signal_850}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_835 ( .s ({signal_7637, signal_7629, signal_7621, signal_7613}), .b ({signal_2693, signal_2692, signal_2691, signal_787}), .a ({signal_2690, signal_2689, signal_2688, signal_786}), .clk ( clk ), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({signal_2888, signal_2887, signal_2886, signal_851}) ) ;
    buf_clk cell_1165 ( .C ( clk ), .D ( signal_7646 ), .Q ( signal_7647 ) ) ;
    buf_clk cell_1175 ( .C ( clk ), .D ( signal_7656 ), .Q ( signal_7657 ) ) ;
    buf_clk cell_1185 ( .C ( clk ), .D ( signal_7666 ), .Q ( signal_7667 ) ) ;
    buf_clk cell_1195 ( .C ( clk ), .D ( signal_7676 ), .Q ( signal_7677 ) ) ;
    buf_clk cell_1205 ( .C ( clk ), .D ( signal_7686 ), .Q ( signal_7687 ) ) ;
    buf_clk cell_1217 ( .C ( clk ), .D ( signal_7698 ), .Q ( signal_7699 ) ) ;
    buf_clk cell_1229 ( .C ( clk ), .D ( signal_7710 ), .Q ( signal_7711 ) ) ;
    buf_clk cell_1241 ( .C ( clk ), .D ( signal_7722 ), .Q ( signal_7723 ) ) ;
    buf_clk cell_1253 ( .C ( clk ), .D ( signal_7734 ), .Q ( signal_7735 ) ) ;
    buf_clk cell_1267 ( .C ( clk ), .D ( signal_7748 ), .Q ( signal_7749 ) ) ;
    buf_clk cell_1281 ( .C ( clk ), .D ( signal_7762 ), .Q ( signal_7763 ) ) ;
    buf_clk cell_1295 ( .C ( clk ), .D ( signal_7776 ), .Q ( signal_7777 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_1206 ( .C ( clk ), .D ( signal_7687 ), .Q ( signal_7688 ) ) ;
    buf_clk cell_1218 ( .C ( clk ), .D ( signal_7699 ), .Q ( signal_7700 ) ) ;
    buf_clk cell_1230 ( .C ( clk ), .D ( signal_7711 ), .Q ( signal_7712 ) ) ;
    buf_clk cell_1242 ( .C ( clk ), .D ( signal_7723 ), .Q ( signal_7724 ) ) ;
    buf_clk cell_1254 ( .C ( clk ), .D ( signal_7735 ), .Q ( signal_7736 ) ) ;
    buf_clk cell_1268 ( .C ( clk ), .D ( signal_7749 ), .Q ( signal_7750 ) ) ;
    buf_clk cell_1282 ( .C ( clk ), .D ( signal_7763 ), .Q ( signal_7764 ) ) ;
    buf_clk cell_1296 ( .C ( clk ), .D ( signal_7777 ), .Q ( signal_7778 ) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_836 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2702, signal_2701, signal_2700, signal_789}), .a ({signal_2699, signal_2698, signal_2697, signal_788}), .clk ( clk ), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({signal_2894, signal_2893, signal_2892, signal_852}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_837 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2708, signal_2707, signal_2706, signal_791}), .a ({signal_2705, signal_2704, signal_2703, signal_790}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({signal_2897, signal_2896, signal_2895, signal_853}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_838 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2714, signal_2713, signal_2712, signal_793}), .a ({signal_2711, signal_2710, signal_2709, signal_792}), .clk ( clk ), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_2900, signal_2899, signal_2898, signal_854}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_839 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2720, signal_2719, signal_2718, signal_795}), .a ({signal_2717, signal_2716, signal_2715, signal_794}), .clk ( clk ), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({signal_2903, signal_2902, signal_2901, signal_855}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_840 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2726, signal_2725, signal_2724, signal_797}), .a ({signal_2723, signal_2722, signal_2721, signal_796}), .clk ( clk ), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({signal_2906, signal_2905, signal_2904, signal_856}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_841 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2732, signal_2731, signal_2730, signal_799}), .a ({signal_2729, signal_2728, signal_2727, signal_798}), .clk ( clk ), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({signal_2909, signal_2908, signal_2907, signal_857}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_842 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2738, signal_2737, signal_2736, signal_801}), .a ({signal_2735, signal_2734, signal_2733, signal_800}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({signal_2912, signal_2911, signal_2910, signal_858}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_843 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2744, signal_2743, signal_2742, signal_803}), .a ({signal_2741, signal_2740, signal_2739, signal_802}), .clk ( clk ), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_2915, signal_2914, signal_2913, signal_859}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_844 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2750, signal_2749, signal_2748, signal_805}), .a ({signal_2747, signal_2746, signal_2745, signal_804}), .clk ( clk ), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({signal_2918, signal_2917, signal_2916, signal_860}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_845 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2756, signal_2755, signal_2754, signal_807}), .a ({signal_2753, signal_2752, signal_2751, signal_806}), .clk ( clk ), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({signal_2921, signal_2920, signal_2919, signal_861}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_846 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2762, signal_2761, signal_2760, signal_809}), .a ({signal_2759, signal_2758, signal_2757, signal_808}), .clk ( clk ), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({signal_2924, signal_2923, signal_2922, signal_862}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_847 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2768, signal_2767, signal_2766, signal_811}), .a ({signal_2765, signal_2764, signal_2763, signal_810}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({signal_2927, signal_2926, signal_2925, signal_863}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_848 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2774, signal_2773, signal_2772, signal_813}), .a ({signal_2771, signal_2770, signal_2769, signal_812}), .clk ( clk ), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_2930, signal_2929, signal_2928, signal_864}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_849 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2780, signal_2779, signal_2778, signal_815}), .a ({signal_2777, signal_2776, signal_2775, signal_814}), .clk ( clk ), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({signal_2933, signal_2932, signal_2931, signal_865}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_850 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2786, signal_2785, signal_2784, signal_817}), .a ({signal_2783, signal_2782, signal_2781, signal_816}), .clk ( clk ), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({signal_2936, signal_2935, signal_2934, signal_866}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_851 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2792, signal_2791, signal_2790, signal_819}), .a ({signal_2789, signal_2788, signal_2787, signal_818}), .clk ( clk ), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({signal_2939, signal_2938, signal_2937, signal_867}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_852 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2798, signal_2797, signal_2796, signal_821}), .a ({signal_2795, signal_2794, signal_2793, signal_820}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({signal_2942, signal_2941, signal_2940, signal_868}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_853 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2804, signal_2803, signal_2802, signal_823}), .a ({signal_2801, signal_2800, signal_2799, signal_822}), .clk ( clk ), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_2945, signal_2944, signal_2943, signal_869}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_854 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2810, signal_2809, signal_2808, signal_825}), .a ({signal_2807, signal_2806, signal_2805, signal_824}), .clk ( clk ), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({signal_2948, signal_2947, signal_2946, signal_870}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_855 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2816, signal_2815, signal_2814, signal_827}), .a ({signal_2813, signal_2812, signal_2811, signal_826}), .clk ( clk ), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({signal_2951, signal_2950, signal_2949, signal_871}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_856 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2822, signal_2821, signal_2820, signal_829}), .a ({signal_2819, signal_2818, signal_2817, signal_828}), .clk ( clk ), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({signal_2954, signal_2953, signal_2952, signal_872}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_857 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2828, signal_2827, signal_2826, signal_831}), .a ({signal_2825, signal_2824, signal_2823, signal_830}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({signal_2957, signal_2956, signal_2955, signal_873}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_858 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2834, signal_2833, signal_2832, signal_833}), .a ({signal_2831, signal_2830, signal_2829, signal_832}), .clk ( clk ), .r ({Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_2960, signal_2959, signal_2958, signal_874}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_859 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2840, signal_2839, signal_2838, signal_835}), .a ({signal_2837, signal_2836, signal_2835, signal_834}), .clk ( clk ), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086]}), .c ({signal_2963, signal_2962, signal_2961, signal_875}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_860 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2846, signal_2845, signal_2844, signal_837}), .a ({signal_2843, signal_2842, signal_2841, signal_836}), .clk ( clk ), .r ({Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({signal_2966, signal_2965, signal_2964, signal_876}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_861 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2852, signal_2851, signal_2850, signal_839}), .a ({signal_2849, signal_2848, signal_2847, signal_838}), .clk ( clk ), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098]}), .c ({signal_2969, signal_2968, signal_2967, signal_877}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_862 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2858, signal_2857, signal_2856, signal_841}), .a ({signal_2855, signal_2854, signal_2853, signal_840}), .clk ( clk ), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({signal_2972, signal_2971, signal_2970, signal_878}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_863 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2864, signal_2863, signal_2862, signal_843}), .a ({signal_2861, signal_2860, signal_2859, signal_842}), .clk ( clk ), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({signal_2975, signal_2974, signal_2973, signal_879}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_864 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2870, signal_2869, signal_2868, signal_845}), .a ({signal_2867, signal_2866, signal_2865, signal_844}), .clk ( clk ), .r ({Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({signal_2978, signal_2977, signal_2976, signal_880}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_865 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2876, signal_2875, signal_2874, signal_847}), .a ({signal_2873, signal_2872, signal_2871, signal_846}), .clk ( clk ), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122]}), .c ({signal_2981, signal_2980, signal_2979, signal_881}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_866 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2882, signal_2881, signal_2880, signal_849}), .a ({signal_2879, signal_2878, signal_2877, signal_848}), .clk ( clk ), .r ({Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({signal_2984, signal_2983, signal_2982, signal_882}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_867 ( .s ({signal_7677, signal_7667, signal_7657, signal_7647}), .b ({signal_2888, signal_2887, signal_2886, signal_851}), .a ({signal_2885, signal_2884, signal_2883, signal_850}), .clk ( clk ), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134]}), .c ({signal_2987, signal_2986, signal_2985, signal_883}) ) ;
    buf_clk cell_1207 ( .C ( clk ), .D ( signal_7688 ), .Q ( signal_7689 ) ) ;
    buf_clk cell_1219 ( .C ( clk ), .D ( signal_7700 ), .Q ( signal_7701 ) ) ;
    buf_clk cell_1231 ( .C ( clk ), .D ( signal_7712 ), .Q ( signal_7713 ) ) ;
    buf_clk cell_1243 ( .C ( clk ), .D ( signal_7724 ), .Q ( signal_7725 ) ) ;
    buf_clk cell_1255 ( .C ( clk ), .D ( signal_7736 ), .Q ( signal_7737 ) ) ;
    buf_clk cell_1269 ( .C ( clk ), .D ( signal_7750 ), .Q ( signal_7751 ) ) ;
    buf_clk cell_1283 ( .C ( clk ), .D ( signal_7764 ), .Q ( signal_7765 ) ) ;
    buf_clk cell_1297 ( .C ( clk ), .D ( signal_7778 ), .Q ( signal_7779 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_1256 ( .C ( clk ), .D ( signal_7737 ), .Q ( signal_7738 ) ) ;
    buf_clk cell_1270 ( .C ( clk ), .D ( signal_7751 ), .Q ( signal_7752 ) ) ;
    buf_clk cell_1284 ( .C ( clk ), .D ( signal_7765 ), .Q ( signal_7766 ) ) ;
    buf_clk cell_1298 ( .C ( clk ), .D ( signal_7779 ), .Q ( signal_7780 ) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_868 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2897, signal_2896, signal_2895, signal_853}), .a ({signal_2894, signal_2893, signal_2892, signal_852}), .clk ( clk ), .r ({Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({signal_2993, signal_2992, signal_2991, signal_884}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_869 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2903, signal_2902, signal_2901, signal_855}), .a ({signal_2900, signal_2899, signal_2898, signal_854}), .clk ( clk ), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146]}), .c ({signal_2996, signal_2995, signal_2994, signal_885}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_870 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2909, signal_2908, signal_2907, signal_857}), .a ({signal_2906, signal_2905, signal_2904, signal_856}), .clk ( clk ), .r ({Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({signal_2999, signal_2998, signal_2997, signal_886}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_871 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2915, signal_2914, signal_2913, signal_859}), .a ({signal_2912, signal_2911, signal_2910, signal_858}), .clk ( clk ), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158]}), .c ({signal_3002, signal_3001, signal_3000, signal_887}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_872 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2921, signal_2920, signal_2919, signal_861}), .a ({signal_2918, signal_2917, signal_2916, signal_860}), .clk ( clk ), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({signal_3005, signal_3004, signal_3003, signal_888}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_873 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2927, signal_2926, signal_2925, signal_863}), .a ({signal_2924, signal_2923, signal_2922, signal_862}), .clk ( clk ), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({signal_3008, signal_3007, signal_3006, signal_889}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_874 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2933, signal_2932, signal_2931, signal_865}), .a ({signal_2930, signal_2929, signal_2928, signal_864}), .clk ( clk ), .r ({Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({signal_3011, signal_3010, signal_3009, signal_890}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_875 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2939, signal_2938, signal_2937, signal_867}), .a ({signal_2936, signal_2935, signal_2934, signal_866}), .clk ( clk ), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182]}), .c ({signal_3014, signal_3013, signal_3012, signal_891}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_876 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2945, signal_2944, signal_2943, signal_869}), .a ({signal_2942, signal_2941, signal_2940, signal_868}), .clk ( clk ), .r ({Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({signal_3017, signal_3016, signal_3015, signal_892}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_877 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2951, signal_2950, signal_2949, signal_871}), .a ({signal_2948, signal_2947, signal_2946, signal_870}), .clk ( clk ), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194]}), .c ({signal_3020, signal_3019, signal_3018, signal_893}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_878 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2957, signal_2956, signal_2955, signal_873}), .a ({signal_2954, signal_2953, signal_2952, signal_872}), .clk ( clk ), .r ({Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({signal_3023, signal_3022, signal_3021, signal_894}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_879 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2963, signal_2962, signal_2961, signal_875}), .a ({signal_2960, signal_2959, signal_2958, signal_874}), .clk ( clk ), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206]}), .c ({signal_3026, signal_3025, signal_3024, signal_895}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_880 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2969, signal_2968, signal_2967, signal_877}), .a ({signal_2966, signal_2965, signal_2964, signal_876}), .clk ( clk ), .r ({Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({signal_3029, signal_3028, signal_3027, signal_896}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_881 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2975, signal_2974, signal_2973, signal_879}), .a ({signal_2972, signal_2971, signal_2970, signal_878}), .clk ( clk ), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218]}), .c ({signal_3032, signal_3031, signal_3030, signal_897}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_882 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2981, signal_2980, signal_2979, signal_881}), .a ({signal_2978, signal_2977, signal_2976, signal_880}), .clk ( clk ), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({signal_3035, signal_3034, signal_3033, signal_898}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_883 ( .s ({signal_7725, signal_7713, signal_7701, signal_7689}), .b ({signal_2987, signal_2986, signal_2985, signal_883}), .a ({signal_2984, signal_2983, signal_2982, signal_882}), .clk ( clk ), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({signal_3038, signal_3037, signal_3036, signal_899}) ) ;
    buf_clk cell_1257 ( .C ( clk ), .D ( signal_7738 ), .Q ( signal_7739 ) ) ;
    buf_clk cell_1271 ( .C ( clk ), .D ( signal_7752 ), .Q ( signal_7753 ) ) ;
    buf_clk cell_1285 ( .C ( clk ), .D ( signal_7766 ), .Q ( signal_7767 ) ) ;
    buf_clk cell_1299 ( .C ( clk ), .D ( signal_7780 ), .Q ( signal_7781 ) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_884 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_2996, signal_2995, signal_2994, signal_885}), .a ({signal_2993, signal_2992, signal_2991, signal_884}), .clk ( clk ), .r ({Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({signal_3044, signal_3043, signal_3042, signal_167}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_885 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3002, signal_3001, signal_3000, signal_887}), .a ({signal_2999, signal_2998, signal_2997, signal_886}), .clk ( clk ), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242]}), .c ({signal_3047, signal_3046, signal_3045, signal_166}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_886 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3008, signal_3007, signal_3006, signal_889}), .a ({signal_3005, signal_3004, signal_3003, signal_888}), .clk ( clk ), .r ({Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({signal_3050, signal_3049, signal_3048, signal_165}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_887 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3014, signal_3013, signal_3012, signal_891}), .a ({signal_3011, signal_3010, signal_3009, signal_890}), .clk ( clk ), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254]}), .c ({signal_3053, signal_3052, signal_3051, signal_164}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_888 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3020, signal_3019, signal_3018, signal_893}), .a ({signal_3017, signal_3016, signal_3015, signal_892}), .clk ( clk ), .r ({Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({signal_3056, signal_3055, signal_3054, signal_163}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_889 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3026, signal_3025, signal_3024, signal_895}), .a ({signal_3023, signal_3022, signal_3021, signal_894}), .clk ( clk ), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266]}), .c ({signal_3059, signal_3058, signal_3057, signal_162}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_890 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3032, signal_3031, signal_3030, signal_897}), .a ({signal_3029, signal_3028, signal_3027, signal_896}), .clk ( clk ), .r ({Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({signal_3062, signal_3061, signal_3060, signal_161}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_891 ( .s ({signal_7781, signal_7767, signal_7753, signal_7739}), .b ({signal_3038, signal_3037, signal_3036, signal_899}), .a ({signal_3035, signal_3034, signal_3033, signal_898}), .clk ( clk ), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278]}), .c ({signal_3065, signal_3064, signal_3063, signal_160}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_3065, signal_3064, signal_3063, signal_160}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_3062, signal_3061, signal_3060, signal_161}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_3059, signal_3058, signal_3057, signal_162}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_3056, signal_3055, signal_3054, signal_163}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_3053, signal_3052, signal_3051, signal_164}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_3050, signal_3049, signal_3048, signal_165}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_3047, signal_3046, signal_3045, signal_166}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_3044, signal_3043, signal_3042, signal_167}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
