////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_round-based/AGEMA/AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d3 (plaintext_s0, key_s0, clk, reset, key_s1, key_s2, key_s3, plaintext_s1, plaintext_s2, plaintext_s3, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, ciphertext_s3);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] plaintext_s3 ;
    input [8159:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output [127:0] ciphertext_s3 ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16253 ;
    wire new_AGEMA_signal_16254 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16264 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16270 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16276 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16282 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16288 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16294 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16300 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16307 ;
    wire new_AGEMA_signal_16308 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16313 ;
    wire new_AGEMA_signal_16314 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16319 ;
    wire new_AGEMA_signal_16320 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16325 ;
    wire new_AGEMA_signal_16326 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16331 ;
    wire new_AGEMA_signal_16332 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16337 ;
    wire new_AGEMA_signal_16338 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16343 ;
    wire new_AGEMA_signal_16344 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16349 ;
    wire new_AGEMA_signal_16350 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16421 ;
    wire new_AGEMA_signal_16422 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16427 ;
    wire new_AGEMA_signal_16428 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16433 ;
    wire new_AGEMA_signal_16434 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16440 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16445 ;
    wire new_AGEMA_signal_16446 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16451 ;
    wire new_AGEMA_signal_16452 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16457 ;
    wire new_AGEMA_signal_16458 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire new_AGEMA_signal_25165 ;
    wire new_AGEMA_signal_25166 ;
    wire new_AGEMA_signal_25167 ;
    wire new_AGEMA_signal_25168 ;
    wire new_AGEMA_signal_25169 ;
    wire new_AGEMA_signal_25170 ;
    wire new_AGEMA_signal_25171 ;
    wire new_AGEMA_signal_25172 ;
    wire new_AGEMA_signal_25173 ;
    wire new_AGEMA_signal_25174 ;
    wire new_AGEMA_signal_25175 ;
    wire new_AGEMA_signal_25176 ;
    wire new_AGEMA_signal_25177 ;
    wire new_AGEMA_signal_25178 ;
    wire new_AGEMA_signal_25179 ;
    wire new_AGEMA_signal_25180 ;
    wire new_AGEMA_signal_25181 ;
    wire new_AGEMA_signal_25182 ;
    wire new_AGEMA_signal_25183 ;
    wire new_AGEMA_signal_25184 ;
    wire new_AGEMA_signal_25185 ;
    wire new_AGEMA_signal_25186 ;
    wire new_AGEMA_signal_25187 ;
    wire new_AGEMA_signal_25188 ;
    wire new_AGEMA_signal_25189 ;
    wire new_AGEMA_signal_25190 ;
    wire new_AGEMA_signal_25191 ;
    wire new_AGEMA_signal_25192 ;
    wire new_AGEMA_signal_25193 ;
    wire new_AGEMA_signal_25194 ;
    wire new_AGEMA_signal_25195 ;
    wire new_AGEMA_signal_25196 ;
    wire new_AGEMA_signal_25197 ;
    wire new_AGEMA_signal_25198 ;
    wire new_AGEMA_signal_25199 ;
    wire new_AGEMA_signal_25200 ;
    wire new_AGEMA_signal_25201 ;
    wire new_AGEMA_signal_25202 ;
    wire new_AGEMA_signal_25203 ;
    wire new_AGEMA_signal_25204 ;
    wire new_AGEMA_signal_25205 ;
    wire new_AGEMA_signal_25206 ;
    wire new_AGEMA_signal_25207 ;
    wire new_AGEMA_signal_25208 ;
    wire new_AGEMA_signal_25209 ;
    wire new_AGEMA_signal_25210 ;
    wire new_AGEMA_signal_25211 ;
    wire new_AGEMA_signal_25212 ;
    wire new_AGEMA_signal_25213 ;
    wire new_AGEMA_signal_25214 ;
    wire new_AGEMA_signal_25215 ;
    wire new_AGEMA_signal_25216 ;
    wire new_AGEMA_signal_25217 ;
    wire new_AGEMA_signal_25218 ;
    wire new_AGEMA_signal_25219 ;
    wire new_AGEMA_signal_25220 ;
    wire new_AGEMA_signal_25221 ;
    wire new_AGEMA_signal_25222 ;
    wire new_AGEMA_signal_25223 ;
    wire new_AGEMA_signal_25224 ;
    wire new_AGEMA_signal_25225 ;
    wire new_AGEMA_signal_25226 ;
    wire new_AGEMA_signal_25227 ;
    wire new_AGEMA_signal_25228 ;
    wire new_AGEMA_signal_25229 ;
    wire new_AGEMA_signal_25230 ;
    wire new_AGEMA_signal_25231 ;
    wire new_AGEMA_signal_25232 ;
    wire new_AGEMA_signal_25233 ;
    wire new_AGEMA_signal_25234 ;
    wire new_AGEMA_signal_25235 ;
    wire new_AGEMA_signal_25236 ;
    wire new_AGEMA_signal_25237 ;
    wire new_AGEMA_signal_25238 ;
    wire new_AGEMA_signal_25239 ;
    wire new_AGEMA_signal_25240 ;
    wire new_AGEMA_signal_25241 ;
    wire new_AGEMA_signal_25242 ;
    wire new_AGEMA_signal_25243 ;
    wire new_AGEMA_signal_25244 ;
    wire new_AGEMA_signal_25245 ;
    wire new_AGEMA_signal_25246 ;
    wire new_AGEMA_signal_25247 ;
    wire new_AGEMA_signal_25248 ;
    wire new_AGEMA_signal_25249 ;
    wire new_AGEMA_signal_25250 ;
    wire new_AGEMA_signal_25251 ;
    wire new_AGEMA_signal_25252 ;
    wire new_AGEMA_signal_25253 ;
    wire new_AGEMA_signal_25254 ;
    wire new_AGEMA_signal_25255 ;
    wire new_AGEMA_signal_25256 ;
    wire new_AGEMA_signal_25257 ;
    wire new_AGEMA_signal_25258 ;
    wire new_AGEMA_signal_25259 ;
    wire new_AGEMA_signal_25260 ;
    wire new_AGEMA_signal_25261 ;
    wire new_AGEMA_signal_25262 ;
    wire new_AGEMA_signal_25263 ;
    wire new_AGEMA_signal_25264 ;
    wire new_AGEMA_signal_25265 ;
    wire new_AGEMA_signal_25266 ;
    wire new_AGEMA_signal_25267 ;
    wire new_AGEMA_signal_25268 ;
    wire new_AGEMA_signal_25269 ;
    wire new_AGEMA_signal_25270 ;
    wire new_AGEMA_signal_25271 ;
    wire new_AGEMA_signal_25272 ;
    wire new_AGEMA_signal_25273 ;
    wire new_AGEMA_signal_25274 ;
    wire new_AGEMA_signal_25275 ;
    wire new_AGEMA_signal_25276 ;
    wire new_AGEMA_signal_25277 ;
    wire new_AGEMA_signal_25278 ;
    wire new_AGEMA_signal_25279 ;
    wire new_AGEMA_signal_25280 ;
    wire new_AGEMA_signal_25281 ;
    wire new_AGEMA_signal_25282 ;
    wire new_AGEMA_signal_25283 ;
    wire new_AGEMA_signal_25284 ;
    wire new_AGEMA_signal_25285 ;
    wire new_AGEMA_signal_25286 ;
    wire new_AGEMA_signal_25287 ;
    wire new_AGEMA_signal_25288 ;
    wire new_AGEMA_signal_25289 ;
    wire new_AGEMA_signal_25290 ;
    wire new_AGEMA_signal_25291 ;
    wire new_AGEMA_signal_25292 ;
    wire new_AGEMA_signal_25293 ;
    wire new_AGEMA_signal_25294 ;
    wire new_AGEMA_signal_25295 ;
    wire new_AGEMA_signal_25296 ;
    wire new_AGEMA_signal_25297 ;
    wire new_AGEMA_signal_25298 ;
    wire new_AGEMA_signal_25299 ;
    wire new_AGEMA_signal_25300 ;
    wire new_AGEMA_signal_25301 ;
    wire new_AGEMA_signal_25302 ;
    wire new_AGEMA_signal_25303 ;
    wire new_AGEMA_signal_25304 ;
    wire new_AGEMA_signal_25305 ;
    wire new_AGEMA_signal_25306 ;
    wire new_AGEMA_signal_25307 ;
    wire new_AGEMA_signal_25308 ;
    wire new_AGEMA_signal_25309 ;
    wire new_AGEMA_signal_25310 ;
    wire new_AGEMA_signal_25311 ;
    wire new_AGEMA_signal_25312 ;
    wire new_AGEMA_signal_25313 ;
    wire new_AGEMA_signal_25314 ;
    wire new_AGEMA_signal_25315 ;
    wire new_AGEMA_signal_25316 ;
    wire new_AGEMA_signal_25317 ;
    wire new_AGEMA_signal_25318 ;
    wire new_AGEMA_signal_25319 ;
    wire new_AGEMA_signal_25320 ;
    wire new_AGEMA_signal_25321 ;
    wire new_AGEMA_signal_25322 ;
    wire new_AGEMA_signal_25323 ;
    wire new_AGEMA_signal_25324 ;
    wire new_AGEMA_signal_25325 ;
    wire new_AGEMA_signal_25326 ;
    wire new_AGEMA_signal_25327 ;
    wire new_AGEMA_signal_25328 ;
    wire new_AGEMA_signal_25329 ;
    wire new_AGEMA_signal_25330 ;
    wire new_AGEMA_signal_25331 ;
    wire new_AGEMA_signal_25332 ;
    wire new_AGEMA_signal_25333 ;
    wire new_AGEMA_signal_25334 ;
    wire new_AGEMA_signal_25335 ;
    wire new_AGEMA_signal_25336 ;
    wire new_AGEMA_signal_25337 ;
    wire new_AGEMA_signal_25338 ;
    wire new_AGEMA_signal_25339 ;
    wire new_AGEMA_signal_25340 ;
    wire new_AGEMA_signal_25341 ;
    wire new_AGEMA_signal_25342 ;
    wire new_AGEMA_signal_25343 ;
    wire new_AGEMA_signal_25344 ;
    wire new_AGEMA_signal_25345 ;
    wire new_AGEMA_signal_25346 ;
    wire new_AGEMA_signal_25347 ;
    wire new_AGEMA_signal_25348 ;
    wire new_AGEMA_signal_25349 ;
    wire new_AGEMA_signal_25350 ;
    wire new_AGEMA_signal_25351 ;
    wire new_AGEMA_signal_25352 ;
    wire new_AGEMA_signal_25353 ;
    wire new_AGEMA_signal_25354 ;
    wire new_AGEMA_signal_25355 ;
    wire new_AGEMA_signal_25356 ;
    wire new_AGEMA_signal_25357 ;
    wire new_AGEMA_signal_25358 ;
    wire new_AGEMA_signal_25359 ;
    wire new_AGEMA_signal_25360 ;
    wire new_AGEMA_signal_25361 ;
    wire new_AGEMA_signal_25362 ;
    wire new_AGEMA_signal_25363 ;
    wire new_AGEMA_signal_25364 ;
    wire new_AGEMA_signal_25365 ;
    wire new_AGEMA_signal_25366 ;
    wire new_AGEMA_signal_25367 ;
    wire new_AGEMA_signal_25368 ;
    wire new_AGEMA_signal_25369 ;
    wire new_AGEMA_signal_25370 ;
    wire new_AGEMA_signal_25371 ;
    wire new_AGEMA_signal_25372 ;
    wire new_AGEMA_signal_25373 ;
    wire new_AGEMA_signal_25374 ;
    wire new_AGEMA_signal_25375 ;
    wire new_AGEMA_signal_25376 ;
    wire new_AGEMA_signal_25377 ;
    wire new_AGEMA_signal_25378 ;
    wire new_AGEMA_signal_25379 ;
    wire new_AGEMA_signal_25380 ;
    wire new_AGEMA_signal_25381 ;
    wire new_AGEMA_signal_25382 ;
    wire new_AGEMA_signal_25383 ;
    wire new_AGEMA_signal_25384 ;
    wire new_AGEMA_signal_25385 ;
    wire new_AGEMA_signal_25386 ;
    wire new_AGEMA_signal_25387 ;
    wire new_AGEMA_signal_25388 ;
    wire new_AGEMA_signal_25389 ;
    wire new_AGEMA_signal_25390 ;
    wire new_AGEMA_signal_25391 ;
    wire new_AGEMA_signal_25392 ;
    wire new_AGEMA_signal_25393 ;
    wire new_AGEMA_signal_25394 ;
    wire new_AGEMA_signal_25395 ;
    wire new_AGEMA_signal_25396 ;
    wire new_AGEMA_signal_25397 ;
    wire new_AGEMA_signal_25398 ;
    wire new_AGEMA_signal_25399 ;
    wire new_AGEMA_signal_25400 ;
    wire new_AGEMA_signal_25401 ;
    wire new_AGEMA_signal_25402 ;
    wire new_AGEMA_signal_25403 ;
    wire new_AGEMA_signal_25404 ;
    wire new_AGEMA_signal_25405 ;
    wire new_AGEMA_signal_25406 ;
    wire new_AGEMA_signal_25407 ;
    wire new_AGEMA_signal_25408 ;
    wire new_AGEMA_signal_25409 ;
    wire new_AGEMA_signal_25410 ;
    wire new_AGEMA_signal_25411 ;
    wire new_AGEMA_signal_25412 ;
    wire new_AGEMA_signal_25413 ;
    wire new_AGEMA_signal_25414 ;
    wire new_AGEMA_signal_25415 ;
    wire new_AGEMA_signal_25416 ;
    wire new_AGEMA_signal_25417 ;
    wire new_AGEMA_signal_25418 ;
    wire new_AGEMA_signal_25419 ;
    wire new_AGEMA_signal_25420 ;
    wire new_AGEMA_signal_25421 ;
    wire new_AGEMA_signal_25422 ;
    wire new_AGEMA_signal_25423 ;
    wire new_AGEMA_signal_25424 ;
    wire new_AGEMA_signal_25425 ;
    wire new_AGEMA_signal_25426 ;
    wire new_AGEMA_signal_25427 ;
    wire new_AGEMA_signal_25428 ;
    wire new_AGEMA_signal_25429 ;
    wire new_AGEMA_signal_25430 ;
    wire new_AGEMA_signal_25431 ;
    wire new_AGEMA_signal_25432 ;
    wire new_AGEMA_signal_25433 ;
    wire new_AGEMA_signal_25434 ;
    wire new_AGEMA_signal_25435 ;
    wire new_AGEMA_signal_25436 ;
    wire new_AGEMA_signal_25437 ;
    wire new_AGEMA_signal_25438 ;
    wire new_AGEMA_signal_25439 ;
    wire new_AGEMA_signal_25440 ;
    wire new_AGEMA_signal_25441 ;
    wire new_AGEMA_signal_25442 ;
    wire new_AGEMA_signal_25443 ;
    wire new_AGEMA_signal_25444 ;
    wire new_AGEMA_signal_25445 ;
    wire new_AGEMA_signal_25446 ;
    wire new_AGEMA_signal_25447 ;
    wire new_AGEMA_signal_25448 ;
    wire new_AGEMA_signal_25449 ;
    wire new_AGEMA_signal_25450 ;
    wire new_AGEMA_signal_25451 ;
    wire new_AGEMA_signal_25452 ;
    wire new_AGEMA_signal_25453 ;
    wire new_AGEMA_signal_25454 ;
    wire new_AGEMA_signal_25455 ;
    wire new_AGEMA_signal_25456 ;
    wire new_AGEMA_signal_25457 ;
    wire new_AGEMA_signal_25458 ;
    wire new_AGEMA_signal_25459 ;
    wire new_AGEMA_signal_25460 ;
    wire new_AGEMA_signal_25461 ;
    wire new_AGEMA_signal_25462 ;
    wire new_AGEMA_signal_25463 ;
    wire new_AGEMA_signal_25464 ;
    wire new_AGEMA_signal_25465 ;
    wire new_AGEMA_signal_25466 ;
    wire new_AGEMA_signal_25467 ;
    wire new_AGEMA_signal_25468 ;
    wire new_AGEMA_signal_25469 ;
    wire new_AGEMA_signal_25470 ;
    wire new_AGEMA_signal_25471 ;
    wire new_AGEMA_signal_25472 ;
    wire new_AGEMA_signal_25473 ;
    wire new_AGEMA_signal_25474 ;
    wire new_AGEMA_signal_25475 ;
    wire new_AGEMA_signal_25476 ;
    wire new_AGEMA_signal_25477 ;
    wire new_AGEMA_signal_25478 ;
    wire new_AGEMA_signal_25479 ;
    wire new_AGEMA_signal_25480 ;
    wire new_AGEMA_signal_25481 ;
    wire new_AGEMA_signal_25482 ;
    wire new_AGEMA_signal_25483 ;
    wire new_AGEMA_signal_25484 ;
    wire new_AGEMA_signal_25485 ;
    wire new_AGEMA_signal_25486 ;
    wire new_AGEMA_signal_25487 ;
    wire new_AGEMA_signal_25488 ;
    wire new_AGEMA_signal_25489 ;
    wire new_AGEMA_signal_25490 ;
    wire new_AGEMA_signal_25491 ;
    wire new_AGEMA_signal_25492 ;
    wire new_AGEMA_signal_25493 ;
    wire new_AGEMA_signal_25494 ;
    wire new_AGEMA_signal_25495 ;
    wire new_AGEMA_signal_25496 ;
    wire new_AGEMA_signal_25497 ;
    wire new_AGEMA_signal_25498 ;
    wire new_AGEMA_signal_25499 ;
    wire new_AGEMA_signal_25500 ;
    wire new_AGEMA_signal_25501 ;
    wire new_AGEMA_signal_25502 ;
    wire new_AGEMA_signal_25503 ;
    wire new_AGEMA_signal_25504 ;
    wire new_AGEMA_signal_25505 ;
    wire new_AGEMA_signal_25506 ;
    wire new_AGEMA_signal_25507 ;
    wire new_AGEMA_signal_25508 ;
    wire new_AGEMA_signal_25509 ;
    wire new_AGEMA_signal_25510 ;
    wire new_AGEMA_signal_25511 ;
    wire new_AGEMA_signal_25512 ;
    wire new_AGEMA_signal_25513 ;
    wire new_AGEMA_signal_25514 ;
    wire new_AGEMA_signal_25515 ;
    wire new_AGEMA_signal_25516 ;
    wire new_AGEMA_signal_25517 ;
    wire new_AGEMA_signal_25518 ;
    wire new_AGEMA_signal_25519 ;
    wire new_AGEMA_signal_25520 ;
    wire new_AGEMA_signal_25521 ;
    wire new_AGEMA_signal_25522 ;
    wire new_AGEMA_signal_25523 ;
    wire new_AGEMA_signal_25524 ;
    wire new_AGEMA_signal_25525 ;
    wire new_AGEMA_signal_25526 ;
    wire new_AGEMA_signal_25527 ;
    wire new_AGEMA_signal_25528 ;
    wire new_AGEMA_signal_25529 ;
    wire new_AGEMA_signal_25530 ;
    wire new_AGEMA_signal_25531 ;
    wire new_AGEMA_signal_25532 ;
    wire new_AGEMA_signal_25533 ;
    wire new_AGEMA_signal_25534 ;
    wire new_AGEMA_signal_25535 ;
    wire new_AGEMA_signal_25536 ;
    wire new_AGEMA_signal_25537 ;
    wire new_AGEMA_signal_25538 ;
    wire new_AGEMA_signal_25539 ;
    wire new_AGEMA_signal_25540 ;
    wire new_AGEMA_signal_25541 ;
    wire new_AGEMA_signal_25542 ;
    wire new_AGEMA_signal_25543 ;
    wire new_AGEMA_signal_25544 ;
    wire new_AGEMA_signal_25545 ;
    wire new_AGEMA_signal_25546 ;
    wire new_AGEMA_signal_25547 ;
    wire new_AGEMA_signal_25548 ;
    wire new_AGEMA_signal_25549 ;
    wire new_AGEMA_signal_25550 ;
    wire new_AGEMA_signal_25551 ;
    wire new_AGEMA_signal_25552 ;
    wire new_AGEMA_signal_25553 ;
    wire new_AGEMA_signal_25554 ;
    wire new_AGEMA_signal_25555 ;
    wire new_AGEMA_signal_25556 ;
    wire new_AGEMA_signal_25557 ;
    wire new_AGEMA_signal_25558 ;
    wire new_AGEMA_signal_25559 ;
    wire new_AGEMA_signal_25560 ;
    wire new_AGEMA_signal_25561 ;
    wire new_AGEMA_signal_25562 ;
    wire new_AGEMA_signal_25563 ;
    wire new_AGEMA_signal_25564 ;
    wire new_AGEMA_signal_25565 ;
    wire new_AGEMA_signal_25566 ;
    wire new_AGEMA_signal_25567 ;
    wire new_AGEMA_signal_25568 ;
    wire new_AGEMA_signal_25569 ;
    wire new_AGEMA_signal_25570 ;
    wire new_AGEMA_signal_25571 ;
    wire new_AGEMA_signal_25572 ;
    wire new_AGEMA_signal_25573 ;
    wire new_AGEMA_signal_25574 ;
    wire new_AGEMA_signal_25575 ;
    wire new_AGEMA_signal_25576 ;
    wire new_AGEMA_signal_25577 ;
    wire new_AGEMA_signal_25578 ;
    wire new_AGEMA_signal_25579 ;
    wire new_AGEMA_signal_25580 ;
    wire new_AGEMA_signal_25581 ;
    wire new_AGEMA_signal_25582 ;
    wire new_AGEMA_signal_25583 ;
    wire new_AGEMA_signal_25584 ;
    wire new_AGEMA_signal_25585 ;
    wire new_AGEMA_signal_25586 ;
    wire new_AGEMA_signal_25587 ;
    wire new_AGEMA_signal_25588 ;
    wire new_AGEMA_signal_25589 ;
    wire new_AGEMA_signal_25590 ;
    wire new_AGEMA_signal_25591 ;
    wire new_AGEMA_signal_25592 ;
    wire new_AGEMA_signal_25593 ;
    wire new_AGEMA_signal_25594 ;
    wire new_AGEMA_signal_25595 ;
    wire new_AGEMA_signal_25596 ;
    wire new_AGEMA_signal_25597 ;
    wire new_AGEMA_signal_25598 ;
    wire new_AGEMA_signal_25599 ;
    wire new_AGEMA_signal_25600 ;
    wire new_AGEMA_signal_25601 ;
    wire new_AGEMA_signal_25602 ;
    wire new_AGEMA_signal_25603 ;
    wire new_AGEMA_signal_25604 ;
    wire new_AGEMA_signal_25605 ;
    wire new_AGEMA_signal_25606 ;
    wire new_AGEMA_signal_25607 ;
    wire new_AGEMA_signal_25608 ;
    wire new_AGEMA_signal_25609 ;
    wire new_AGEMA_signal_25610 ;
    wire new_AGEMA_signal_25611 ;
    wire new_AGEMA_signal_25612 ;
    wire new_AGEMA_signal_25613 ;
    wire new_AGEMA_signal_25614 ;
    wire new_AGEMA_signal_25615 ;
    wire new_AGEMA_signal_25616 ;
    wire new_AGEMA_signal_25617 ;
    wire new_AGEMA_signal_25618 ;
    wire new_AGEMA_signal_25619 ;
    wire new_AGEMA_signal_25620 ;
    wire new_AGEMA_signal_25621 ;
    wire new_AGEMA_signal_25622 ;
    wire new_AGEMA_signal_25623 ;
    wire new_AGEMA_signal_25624 ;
    wire new_AGEMA_signal_25625 ;
    wire new_AGEMA_signal_25626 ;
    wire new_AGEMA_signal_25627 ;
    wire new_AGEMA_signal_25628 ;
    wire new_AGEMA_signal_25629 ;
    wire new_AGEMA_signal_25630 ;
    wire new_AGEMA_signal_25631 ;
    wire new_AGEMA_signal_25632 ;
    wire new_AGEMA_signal_25633 ;
    wire new_AGEMA_signal_25634 ;
    wire new_AGEMA_signal_25635 ;
    wire new_AGEMA_signal_25636 ;
    wire new_AGEMA_signal_25637 ;
    wire new_AGEMA_signal_25638 ;
    wire new_AGEMA_signal_25639 ;
    wire new_AGEMA_signal_25640 ;
    wire new_AGEMA_signal_25641 ;
    wire new_AGEMA_signal_25642 ;
    wire new_AGEMA_signal_25643 ;
    wire new_AGEMA_signal_25644 ;
    wire new_AGEMA_signal_25645 ;
    wire new_AGEMA_signal_25646 ;
    wire new_AGEMA_signal_25647 ;
    wire new_AGEMA_signal_25648 ;
    wire new_AGEMA_signal_25649 ;
    wire new_AGEMA_signal_25650 ;
    wire new_AGEMA_signal_25651 ;
    wire new_AGEMA_signal_25652 ;
    wire new_AGEMA_signal_25653 ;
    wire new_AGEMA_signal_25654 ;
    wire new_AGEMA_signal_25655 ;
    wire new_AGEMA_signal_25656 ;
    wire new_AGEMA_signal_25657 ;
    wire new_AGEMA_signal_25658 ;
    wire new_AGEMA_signal_25659 ;
    wire new_AGEMA_signal_25660 ;
    wire new_AGEMA_signal_25661 ;
    wire new_AGEMA_signal_25662 ;
    wire new_AGEMA_signal_25663 ;
    wire new_AGEMA_signal_25664 ;
    wire new_AGEMA_signal_25665 ;
    wire new_AGEMA_signal_25666 ;
    wire new_AGEMA_signal_25667 ;
    wire new_AGEMA_signal_25668 ;
    wire new_AGEMA_signal_25669 ;
    wire new_AGEMA_signal_25670 ;
    wire new_AGEMA_signal_25671 ;
    wire new_AGEMA_signal_25672 ;
    wire new_AGEMA_signal_25673 ;
    wire new_AGEMA_signal_25674 ;
    wire new_AGEMA_signal_25675 ;
    wire new_AGEMA_signal_25676 ;
    wire new_AGEMA_signal_25677 ;
    wire new_AGEMA_signal_25678 ;
    wire new_AGEMA_signal_25679 ;
    wire new_AGEMA_signal_25680 ;
    wire new_AGEMA_signal_25681 ;
    wire new_AGEMA_signal_25682 ;
    wire new_AGEMA_signal_25683 ;
    wire new_AGEMA_signal_25684 ;
    wire new_AGEMA_signal_25685 ;
    wire new_AGEMA_signal_25686 ;
    wire new_AGEMA_signal_25687 ;
    wire new_AGEMA_signal_25688 ;
    wire new_AGEMA_signal_25689 ;
    wire new_AGEMA_signal_25690 ;
    wire new_AGEMA_signal_25691 ;
    wire new_AGEMA_signal_25692 ;
    wire new_AGEMA_signal_25693 ;
    wire new_AGEMA_signal_25694 ;
    wire new_AGEMA_signal_25695 ;
    wire new_AGEMA_signal_25696 ;
    wire new_AGEMA_signal_25697 ;
    wire new_AGEMA_signal_25698 ;
    wire new_AGEMA_signal_25699 ;
    wire new_AGEMA_signal_25700 ;
    wire new_AGEMA_signal_25701 ;
    wire new_AGEMA_signal_25702 ;
    wire new_AGEMA_signal_25703 ;
    wire new_AGEMA_signal_25704 ;
    wire new_AGEMA_signal_25705 ;
    wire new_AGEMA_signal_25706 ;
    wire new_AGEMA_signal_25707 ;
    wire new_AGEMA_signal_25708 ;
    wire new_AGEMA_signal_25709 ;
    wire new_AGEMA_signal_25710 ;
    wire new_AGEMA_signal_25711 ;
    wire new_AGEMA_signal_25712 ;
    wire new_AGEMA_signal_25713 ;
    wire new_AGEMA_signal_25714 ;
    wire new_AGEMA_signal_25715 ;
    wire new_AGEMA_signal_25716 ;
    wire new_AGEMA_signal_25717 ;
    wire new_AGEMA_signal_25718 ;
    wire new_AGEMA_signal_25719 ;
    wire new_AGEMA_signal_25720 ;
    wire new_AGEMA_signal_25721 ;
    wire new_AGEMA_signal_25722 ;
    wire new_AGEMA_signal_25723 ;
    wire new_AGEMA_signal_25724 ;
    wire new_AGEMA_signal_25725 ;
    wire new_AGEMA_signal_25726 ;
    wire new_AGEMA_signal_25727 ;
    wire new_AGEMA_signal_25728 ;
    wire new_AGEMA_signal_25729 ;
    wire new_AGEMA_signal_25730 ;
    wire new_AGEMA_signal_25731 ;
    wire new_AGEMA_signal_25732 ;
    wire new_AGEMA_signal_25733 ;
    wire new_AGEMA_signal_25734 ;
    wire new_AGEMA_signal_25735 ;
    wire new_AGEMA_signal_25736 ;
    wire new_AGEMA_signal_25737 ;
    wire new_AGEMA_signal_25738 ;
    wire new_AGEMA_signal_25739 ;
    wire new_AGEMA_signal_25740 ;
    wire new_AGEMA_signal_25741 ;
    wire new_AGEMA_signal_25742 ;
    wire new_AGEMA_signal_25743 ;
    wire new_AGEMA_signal_25744 ;
    wire new_AGEMA_signal_25745 ;
    wire new_AGEMA_signal_25746 ;
    wire new_AGEMA_signal_25747 ;
    wire new_AGEMA_signal_25748 ;
    wire new_AGEMA_signal_25749 ;
    wire new_AGEMA_signal_25750 ;
    wire new_AGEMA_signal_25751 ;
    wire new_AGEMA_signal_25752 ;
    wire new_AGEMA_signal_25753 ;
    wire new_AGEMA_signal_25754 ;
    wire new_AGEMA_signal_25755 ;
    wire new_AGEMA_signal_25756 ;
    wire new_AGEMA_signal_25757 ;
    wire new_AGEMA_signal_25758 ;
    wire new_AGEMA_signal_25759 ;
    wire new_AGEMA_signal_25760 ;
    wire new_AGEMA_signal_25761 ;
    wire new_AGEMA_signal_25762 ;
    wire new_AGEMA_signal_25763 ;
    wire new_AGEMA_signal_25764 ;
    wire new_AGEMA_signal_25765 ;
    wire new_AGEMA_signal_25766 ;
    wire new_AGEMA_signal_25767 ;
    wire new_AGEMA_signal_25768 ;
    wire new_AGEMA_signal_25769 ;
    wire new_AGEMA_signal_25770 ;
    wire new_AGEMA_signal_25771 ;
    wire new_AGEMA_signal_25772 ;
    wire new_AGEMA_signal_25773 ;
    wire new_AGEMA_signal_25774 ;
    wire new_AGEMA_signal_25775 ;
    wire new_AGEMA_signal_25776 ;
    wire new_AGEMA_signal_25777 ;
    wire new_AGEMA_signal_25778 ;
    wire new_AGEMA_signal_25779 ;
    wire new_AGEMA_signal_25780 ;
    wire new_AGEMA_signal_25781 ;
    wire new_AGEMA_signal_25782 ;
    wire new_AGEMA_signal_25783 ;
    wire new_AGEMA_signal_25784 ;
    wire new_AGEMA_signal_25785 ;
    wire new_AGEMA_signal_25786 ;
    wire new_AGEMA_signal_25787 ;
    wire new_AGEMA_signal_25788 ;
    wire new_AGEMA_signal_25789 ;
    wire new_AGEMA_signal_25790 ;
    wire new_AGEMA_signal_25791 ;
    wire new_AGEMA_signal_25792 ;
    wire new_AGEMA_signal_25793 ;
    wire new_AGEMA_signal_25794 ;
    wire new_AGEMA_signal_25795 ;
    wire new_AGEMA_signal_25796 ;
    wire new_AGEMA_signal_25797 ;
    wire new_AGEMA_signal_25798 ;
    wire new_AGEMA_signal_25799 ;
    wire new_AGEMA_signal_25800 ;
    wire new_AGEMA_signal_25801 ;
    wire new_AGEMA_signal_25802 ;
    wire new_AGEMA_signal_25803 ;
    wire new_AGEMA_signal_25804 ;
    wire new_AGEMA_signal_25805 ;
    wire new_AGEMA_signal_25806 ;
    wire new_AGEMA_signal_25807 ;
    wire new_AGEMA_signal_25808 ;
    wire new_AGEMA_signal_25809 ;
    wire new_AGEMA_signal_25810 ;
    wire new_AGEMA_signal_25811 ;
    wire new_AGEMA_signal_25812 ;
    wire new_AGEMA_signal_25813 ;
    wire new_AGEMA_signal_25814 ;
    wire new_AGEMA_signal_25815 ;
    wire new_AGEMA_signal_25816 ;
    wire new_AGEMA_signal_25817 ;
    wire new_AGEMA_signal_25818 ;
    wire new_AGEMA_signal_25819 ;
    wire new_AGEMA_signal_25820 ;
    wire new_AGEMA_signal_25821 ;
    wire new_AGEMA_signal_25822 ;
    wire new_AGEMA_signal_25823 ;
    wire new_AGEMA_signal_25824 ;
    wire new_AGEMA_signal_25825 ;
    wire new_AGEMA_signal_25826 ;
    wire new_AGEMA_signal_25827 ;
    wire new_AGEMA_signal_25828 ;
    wire new_AGEMA_signal_25829 ;
    wire new_AGEMA_signal_25830 ;
    wire new_AGEMA_signal_25831 ;
    wire new_AGEMA_signal_25832 ;
    wire new_AGEMA_signal_25833 ;
    wire new_AGEMA_signal_25834 ;
    wire new_AGEMA_signal_25835 ;
    wire new_AGEMA_signal_25836 ;
    wire new_AGEMA_signal_25837 ;
    wire new_AGEMA_signal_25838 ;
    wire new_AGEMA_signal_25839 ;
    wire new_AGEMA_signal_25840 ;
    wire new_AGEMA_signal_25841 ;
    wire new_AGEMA_signal_25842 ;
    wire new_AGEMA_signal_25843 ;
    wire new_AGEMA_signal_25844 ;
    wire new_AGEMA_signal_25845 ;
    wire new_AGEMA_signal_25846 ;
    wire new_AGEMA_signal_25847 ;
    wire new_AGEMA_signal_25848 ;
    wire new_AGEMA_signal_25849 ;
    wire new_AGEMA_signal_25850 ;
    wire new_AGEMA_signal_25851 ;
    wire new_AGEMA_signal_25852 ;
    wire new_AGEMA_signal_25853 ;
    wire new_AGEMA_signal_25854 ;
    wire new_AGEMA_signal_25855 ;
    wire new_AGEMA_signal_25856 ;
    wire new_AGEMA_signal_25857 ;
    wire new_AGEMA_signal_25858 ;
    wire new_AGEMA_signal_25859 ;
    wire new_AGEMA_signal_25860 ;
    wire new_AGEMA_signal_25861 ;
    wire new_AGEMA_signal_25862 ;
    wire new_AGEMA_signal_25863 ;
    wire new_AGEMA_signal_25864 ;
    wire new_AGEMA_signal_25865 ;
    wire new_AGEMA_signal_25866 ;
    wire new_AGEMA_signal_25867 ;
    wire new_AGEMA_signal_25868 ;
    wire new_AGEMA_signal_25869 ;
    wire new_AGEMA_signal_25870 ;
    wire new_AGEMA_signal_25871 ;
    wire new_AGEMA_signal_25872 ;
    wire new_AGEMA_signal_25873 ;
    wire new_AGEMA_signal_25874 ;
    wire new_AGEMA_signal_25875 ;
    wire new_AGEMA_signal_25876 ;
    wire new_AGEMA_signal_25877 ;
    wire new_AGEMA_signal_25878 ;
    wire new_AGEMA_signal_25879 ;
    wire new_AGEMA_signal_25880 ;
    wire new_AGEMA_signal_25881 ;
    wire new_AGEMA_signal_25882 ;
    wire new_AGEMA_signal_25883 ;
    wire new_AGEMA_signal_25884 ;
    wire new_AGEMA_signal_25885 ;
    wire new_AGEMA_signal_25886 ;
    wire new_AGEMA_signal_25887 ;
    wire new_AGEMA_signal_25888 ;
    wire new_AGEMA_signal_25889 ;
    wire new_AGEMA_signal_25890 ;
    wire new_AGEMA_signal_25891 ;
    wire new_AGEMA_signal_25892 ;
    wire new_AGEMA_signal_25893 ;
    wire new_AGEMA_signal_25894 ;
    wire new_AGEMA_signal_25895 ;
    wire new_AGEMA_signal_25896 ;
    wire new_AGEMA_signal_25897 ;
    wire new_AGEMA_signal_25898 ;
    wire new_AGEMA_signal_25899 ;
    wire new_AGEMA_signal_25900 ;
    wire new_AGEMA_signal_25901 ;
    wire new_AGEMA_signal_25902 ;
    wire new_AGEMA_signal_25903 ;
    wire new_AGEMA_signal_25904 ;
    wire new_AGEMA_signal_25905 ;
    wire new_AGEMA_signal_25906 ;
    wire new_AGEMA_signal_25907 ;
    wire new_AGEMA_signal_25908 ;
    wire new_AGEMA_signal_25909 ;
    wire new_AGEMA_signal_25910 ;
    wire new_AGEMA_signal_25911 ;
    wire new_AGEMA_signal_25912 ;
    wire new_AGEMA_signal_25913 ;
    wire new_AGEMA_signal_25914 ;
    wire new_AGEMA_signal_25915 ;
    wire new_AGEMA_signal_25916 ;
    wire new_AGEMA_signal_25917 ;
    wire new_AGEMA_signal_25918 ;
    wire new_AGEMA_signal_25919 ;
    wire new_AGEMA_signal_25920 ;
    wire new_AGEMA_signal_25921 ;
    wire new_AGEMA_signal_25922 ;
    wire new_AGEMA_signal_25923 ;
    wire new_AGEMA_signal_25924 ;
    wire new_AGEMA_signal_25925 ;
    wire new_AGEMA_signal_25926 ;
    wire new_AGEMA_signal_25927 ;
    wire new_AGEMA_signal_25928 ;
    wire new_AGEMA_signal_25929 ;
    wire new_AGEMA_signal_25930 ;
    wire new_AGEMA_signal_25931 ;
    wire new_AGEMA_signal_25932 ;
    wire new_AGEMA_signal_25933 ;
    wire new_AGEMA_signal_25934 ;
    wire new_AGEMA_signal_25935 ;
    wire new_AGEMA_signal_25936 ;
    wire new_AGEMA_signal_25937 ;
    wire new_AGEMA_signal_25938 ;
    wire new_AGEMA_signal_25939 ;
    wire new_AGEMA_signal_25940 ;
    wire new_AGEMA_signal_25941 ;
    wire new_AGEMA_signal_25942 ;
    wire new_AGEMA_signal_25943 ;
    wire new_AGEMA_signal_25944 ;
    wire new_AGEMA_signal_25945 ;
    wire new_AGEMA_signal_25946 ;
    wire new_AGEMA_signal_25947 ;
    wire new_AGEMA_signal_25948 ;
    wire new_AGEMA_signal_25949 ;
    wire new_AGEMA_signal_25950 ;
    wire new_AGEMA_signal_25951 ;
    wire new_AGEMA_signal_25952 ;
    wire new_AGEMA_signal_25953 ;
    wire new_AGEMA_signal_25954 ;
    wire new_AGEMA_signal_25955 ;
    wire new_AGEMA_signal_25956 ;
    wire new_AGEMA_signal_25957 ;
    wire new_AGEMA_signal_25958 ;
    wire new_AGEMA_signal_25959 ;
    wire new_AGEMA_signal_25960 ;
    wire new_AGEMA_signal_25961 ;
    wire new_AGEMA_signal_25962 ;
    wire new_AGEMA_signal_25963 ;
    wire new_AGEMA_signal_25964 ;
    wire new_AGEMA_signal_25965 ;
    wire new_AGEMA_signal_25966 ;
    wire new_AGEMA_signal_25967 ;
    wire new_AGEMA_signal_25968 ;
    wire new_AGEMA_signal_25969 ;
    wire new_AGEMA_signal_25970 ;
    wire new_AGEMA_signal_25971 ;
    wire new_AGEMA_signal_25972 ;
    wire new_AGEMA_signal_25973 ;
    wire new_AGEMA_signal_25974 ;
    wire new_AGEMA_signal_25975 ;
    wire new_AGEMA_signal_25976 ;
    wire new_AGEMA_signal_25977 ;
    wire new_AGEMA_signal_25978 ;
    wire new_AGEMA_signal_25979 ;
    wire new_AGEMA_signal_25980 ;
    wire new_AGEMA_signal_25981 ;
    wire new_AGEMA_signal_25982 ;
    wire new_AGEMA_signal_25983 ;
    wire new_AGEMA_signal_25984 ;
    wire new_AGEMA_signal_25985 ;
    wire new_AGEMA_signal_25986 ;
    wire new_AGEMA_signal_25987 ;
    wire new_AGEMA_signal_25988 ;
    wire new_AGEMA_signal_25989 ;
    wire new_AGEMA_signal_25990 ;
    wire new_AGEMA_signal_25991 ;
    wire new_AGEMA_signal_25992 ;
    wire new_AGEMA_signal_25993 ;
    wire new_AGEMA_signal_25994 ;
    wire new_AGEMA_signal_25995 ;
    wire new_AGEMA_signal_25996 ;
    wire new_AGEMA_signal_25997 ;
    wire new_AGEMA_signal_25998 ;
    wire new_AGEMA_signal_25999 ;
    wire new_AGEMA_signal_26000 ;
    wire new_AGEMA_signal_26001 ;
    wire new_AGEMA_signal_26002 ;
    wire new_AGEMA_signal_26003 ;
    wire new_AGEMA_signal_26004 ;
    wire new_AGEMA_signal_26005 ;
    wire new_AGEMA_signal_26006 ;
    wire new_AGEMA_signal_26007 ;
    wire new_AGEMA_signal_26008 ;
    wire new_AGEMA_signal_26009 ;
    wire new_AGEMA_signal_26010 ;
    wire new_AGEMA_signal_26011 ;
    wire new_AGEMA_signal_26012 ;
    wire new_AGEMA_signal_26013 ;
    wire new_AGEMA_signal_26014 ;
    wire new_AGEMA_signal_26015 ;
    wire new_AGEMA_signal_26016 ;
    wire new_AGEMA_signal_26017 ;
    wire new_AGEMA_signal_26018 ;
    wire new_AGEMA_signal_26019 ;
    wire new_AGEMA_signal_26020 ;
    wire new_AGEMA_signal_26021 ;
    wire new_AGEMA_signal_26022 ;
    wire new_AGEMA_signal_26023 ;
    wire new_AGEMA_signal_26024 ;
    wire new_AGEMA_signal_26025 ;
    wire new_AGEMA_signal_26026 ;
    wire new_AGEMA_signal_26027 ;
    wire new_AGEMA_signal_26028 ;
    wire new_AGEMA_signal_26029 ;
    wire new_AGEMA_signal_26030 ;
    wire new_AGEMA_signal_26031 ;
    wire new_AGEMA_signal_26032 ;
    wire new_AGEMA_signal_26033 ;
    wire new_AGEMA_signal_26034 ;
    wire new_AGEMA_signal_26035 ;
    wire new_AGEMA_signal_26036 ;
    wire new_AGEMA_signal_26037 ;
    wire new_AGEMA_signal_26038 ;
    wire new_AGEMA_signal_26039 ;
    wire new_AGEMA_signal_26040 ;
    wire new_AGEMA_signal_26041 ;
    wire new_AGEMA_signal_26042 ;
    wire new_AGEMA_signal_26043 ;
    wire new_AGEMA_signal_26044 ;
    wire new_AGEMA_signal_26045 ;
    wire new_AGEMA_signal_26046 ;
    wire new_AGEMA_signal_26047 ;
    wire new_AGEMA_signal_26048 ;
    wire new_AGEMA_signal_26049 ;
    wire new_AGEMA_signal_26050 ;
    wire new_AGEMA_signal_26051 ;
    wire new_AGEMA_signal_26052 ;
    wire new_AGEMA_signal_26053 ;
    wire new_AGEMA_signal_26054 ;
    wire new_AGEMA_signal_26055 ;
    wire new_AGEMA_signal_26056 ;
    wire new_AGEMA_signal_26057 ;
    wire new_AGEMA_signal_26058 ;
    wire new_AGEMA_signal_26059 ;
    wire new_AGEMA_signal_26060 ;
    wire new_AGEMA_signal_26061 ;
    wire new_AGEMA_signal_26062 ;
    wire new_AGEMA_signal_26063 ;
    wire new_AGEMA_signal_26064 ;
    wire new_AGEMA_signal_26065 ;
    wire new_AGEMA_signal_26066 ;
    wire new_AGEMA_signal_26067 ;
    wire new_AGEMA_signal_26068 ;
    wire new_AGEMA_signal_26069 ;
    wire new_AGEMA_signal_26070 ;
    wire new_AGEMA_signal_26071 ;
    wire new_AGEMA_signal_26072 ;
    wire new_AGEMA_signal_26073 ;
    wire new_AGEMA_signal_26074 ;
    wire new_AGEMA_signal_26075 ;
    wire new_AGEMA_signal_26076 ;
    wire new_AGEMA_signal_26077 ;
    wire new_AGEMA_signal_26078 ;
    wire new_AGEMA_signal_26079 ;
    wire new_AGEMA_signal_26080 ;
    wire new_AGEMA_signal_26081 ;
    wire new_AGEMA_signal_26082 ;
    wire new_AGEMA_signal_26083 ;
    wire new_AGEMA_signal_26084 ;
    wire new_AGEMA_signal_26085 ;
    wire new_AGEMA_signal_26086 ;
    wire new_AGEMA_signal_26087 ;
    wire new_AGEMA_signal_26088 ;
    wire new_AGEMA_signal_26089 ;
    wire new_AGEMA_signal_26090 ;
    wire new_AGEMA_signal_26091 ;
    wire new_AGEMA_signal_26092 ;
    wire new_AGEMA_signal_26093 ;
    wire new_AGEMA_signal_26094 ;
    wire new_AGEMA_signal_26095 ;
    wire new_AGEMA_signal_26096 ;
    wire new_AGEMA_signal_26097 ;
    wire new_AGEMA_signal_26098 ;
    wire new_AGEMA_signal_26099 ;
    wire new_AGEMA_signal_26100 ;
    wire new_AGEMA_signal_26101 ;
    wire new_AGEMA_signal_26102 ;
    wire new_AGEMA_signal_26103 ;
    wire new_AGEMA_signal_26104 ;
    wire new_AGEMA_signal_26105 ;
    wire new_AGEMA_signal_26106 ;
    wire new_AGEMA_signal_26107 ;
    wire new_AGEMA_signal_26108 ;
    wire new_AGEMA_signal_26109 ;
    wire new_AGEMA_signal_26110 ;
    wire new_AGEMA_signal_26111 ;
    wire new_AGEMA_signal_26112 ;
    wire new_AGEMA_signal_26113 ;
    wire new_AGEMA_signal_26114 ;
    wire new_AGEMA_signal_26115 ;
    wire new_AGEMA_signal_26116 ;
    wire new_AGEMA_signal_26117 ;
    wire new_AGEMA_signal_26118 ;
    wire new_AGEMA_signal_26119 ;
    wire new_AGEMA_signal_26120 ;
    wire new_AGEMA_signal_26121 ;
    wire new_AGEMA_signal_26122 ;
    wire new_AGEMA_signal_26123 ;
    wire new_AGEMA_signal_26124 ;
    wire new_AGEMA_signal_26125 ;
    wire new_AGEMA_signal_26126 ;
    wire new_AGEMA_signal_26127 ;
    wire new_AGEMA_signal_26128 ;
    wire new_AGEMA_signal_26129 ;
    wire new_AGEMA_signal_26130 ;
    wire new_AGEMA_signal_26131 ;
    wire new_AGEMA_signal_26132 ;
    wire new_AGEMA_signal_26133 ;
    wire new_AGEMA_signal_26134 ;
    wire new_AGEMA_signal_26135 ;
    wire new_AGEMA_signal_26136 ;
    wire new_AGEMA_signal_26137 ;
    wire new_AGEMA_signal_26138 ;
    wire new_AGEMA_signal_26139 ;
    wire new_AGEMA_signal_26140 ;
    wire new_AGEMA_signal_26141 ;
    wire new_AGEMA_signal_26142 ;
    wire new_AGEMA_signal_26143 ;
    wire new_AGEMA_signal_26144 ;
    wire new_AGEMA_signal_26145 ;
    wire new_AGEMA_signal_26146 ;
    wire new_AGEMA_signal_26147 ;
    wire new_AGEMA_signal_26148 ;
    wire new_AGEMA_signal_26149 ;
    wire new_AGEMA_signal_26150 ;
    wire new_AGEMA_signal_26151 ;
    wire new_AGEMA_signal_26152 ;
    wire new_AGEMA_signal_26153 ;
    wire new_AGEMA_signal_26154 ;
    wire new_AGEMA_signal_26155 ;
    wire new_AGEMA_signal_26156 ;
    wire new_AGEMA_signal_26157 ;
    wire new_AGEMA_signal_26158 ;
    wire new_AGEMA_signal_26159 ;
    wire new_AGEMA_signal_26160 ;
    wire new_AGEMA_signal_26161 ;
    wire new_AGEMA_signal_26162 ;
    wire new_AGEMA_signal_26163 ;
    wire new_AGEMA_signal_26164 ;
    wire new_AGEMA_signal_26165 ;
    wire new_AGEMA_signal_26166 ;
    wire new_AGEMA_signal_26167 ;
    wire new_AGEMA_signal_26168 ;
    wire new_AGEMA_signal_26169 ;
    wire new_AGEMA_signal_26170 ;
    wire new_AGEMA_signal_26171 ;
    wire new_AGEMA_signal_26172 ;
    wire new_AGEMA_signal_26173 ;
    wire new_AGEMA_signal_26174 ;
    wire new_AGEMA_signal_26175 ;
    wire new_AGEMA_signal_26176 ;
    wire new_AGEMA_signal_26177 ;
    wire new_AGEMA_signal_26178 ;
    wire new_AGEMA_signal_26179 ;
    wire new_AGEMA_signal_26180 ;
    wire new_AGEMA_signal_26181 ;
    wire new_AGEMA_signal_26182 ;
    wire new_AGEMA_signal_26183 ;
    wire new_AGEMA_signal_26184 ;
    wire new_AGEMA_signal_26185 ;
    wire new_AGEMA_signal_26186 ;
    wire new_AGEMA_signal_26187 ;
    wire new_AGEMA_signal_26188 ;
    wire new_AGEMA_signal_26189 ;
    wire new_AGEMA_signal_26190 ;
    wire new_AGEMA_signal_26191 ;
    wire new_AGEMA_signal_26192 ;
    wire new_AGEMA_signal_26193 ;
    wire new_AGEMA_signal_26194 ;
    wire new_AGEMA_signal_26195 ;
    wire new_AGEMA_signal_26196 ;
    wire new_AGEMA_signal_26197 ;
    wire new_AGEMA_signal_26198 ;
    wire new_AGEMA_signal_26199 ;
    wire new_AGEMA_signal_26200 ;
    wire new_AGEMA_signal_26201 ;
    wire new_AGEMA_signal_26202 ;
    wire new_AGEMA_signal_26203 ;
    wire new_AGEMA_signal_26204 ;
    wire new_AGEMA_signal_26205 ;
    wire new_AGEMA_signal_26206 ;
    wire new_AGEMA_signal_26207 ;
    wire new_AGEMA_signal_26208 ;
    wire new_AGEMA_signal_26209 ;
    wire new_AGEMA_signal_26210 ;
    wire new_AGEMA_signal_26211 ;
    wire new_AGEMA_signal_26212 ;
    wire new_AGEMA_signal_26213 ;
    wire new_AGEMA_signal_26214 ;
    wire new_AGEMA_signal_26215 ;
    wire new_AGEMA_signal_26216 ;
    wire new_AGEMA_signal_26217 ;
    wire new_AGEMA_signal_26218 ;
    wire new_AGEMA_signal_26219 ;
    wire new_AGEMA_signal_26220 ;
    wire new_AGEMA_signal_26221 ;
    wire new_AGEMA_signal_26222 ;
    wire new_AGEMA_signal_26223 ;
    wire new_AGEMA_signal_26224 ;
    wire new_AGEMA_signal_26225 ;
    wire new_AGEMA_signal_26226 ;
    wire new_AGEMA_signal_26227 ;
    wire new_AGEMA_signal_26228 ;
    wire new_AGEMA_signal_26229 ;
    wire new_AGEMA_signal_26230 ;
    wire new_AGEMA_signal_26231 ;
    wire new_AGEMA_signal_26232 ;
    wire new_AGEMA_signal_26233 ;
    wire new_AGEMA_signal_26234 ;
    wire new_AGEMA_signal_26235 ;
    wire new_AGEMA_signal_26236 ;
    wire new_AGEMA_signal_26237 ;
    wire new_AGEMA_signal_26238 ;
    wire new_AGEMA_signal_26239 ;
    wire new_AGEMA_signal_26240 ;
    wire new_AGEMA_signal_26241 ;
    wire new_AGEMA_signal_26242 ;
    wire new_AGEMA_signal_26243 ;
    wire new_AGEMA_signal_26244 ;
    wire new_AGEMA_signal_26245 ;
    wire new_AGEMA_signal_26246 ;
    wire new_AGEMA_signal_26247 ;
    wire new_AGEMA_signal_26248 ;
    wire new_AGEMA_signal_26249 ;
    wire new_AGEMA_signal_26250 ;
    wire new_AGEMA_signal_26251 ;
    wire new_AGEMA_signal_26252 ;
    wire new_AGEMA_signal_26253 ;
    wire new_AGEMA_signal_26254 ;
    wire new_AGEMA_signal_26255 ;
    wire new_AGEMA_signal_26256 ;
    wire new_AGEMA_signal_26257 ;
    wire new_AGEMA_signal_26258 ;
    wire new_AGEMA_signal_26259 ;
    wire new_AGEMA_signal_26260 ;
    wire new_AGEMA_signal_26261 ;
    wire new_AGEMA_signal_26262 ;
    wire new_AGEMA_signal_26263 ;
    wire new_AGEMA_signal_26264 ;
    wire new_AGEMA_signal_26265 ;
    wire new_AGEMA_signal_26266 ;
    wire new_AGEMA_signal_26267 ;
    wire new_AGEMA_signal_26268 ;
    wire new_AGEMA_signal_26269 ;
    wire new_AGEMA_signal_26270 ;
    wire new_AGEMA_signal_26271 ;
    wire new_AGEMA_signal_26272 ;
    wire new_AGEMA_signal_26273 ;
    wire new_AGEMA_signal_26274 ;
    wire new_AGEMA_signal_26275 ;
    wire new_AGEMA_signal_26276 ;
    wire new_AGEMA_signal_26277 ;
    wire new_AGEMA_signal_26278 ;
    wire new_AGEMA_signal_26279 ;
    wire new_AGEMA_signal_26280 ;
    wire new_AGEMA_signal_26281 ;
    wire new_AGEMA_signal_26282 ;
    wire new_AGEMA_signal_26283 ;
    wire new_AGEMA_signal_26284 ;
    wire new_AGEMA_signal_26285 ;
    wire new_AGEMA_signal_26286 ;
    wire new_AGEMA_signal_26287 ;
    wire new_AGEMA_signal_26288 ;
    wire new_AGEMA_signal_26289 ;
    wire new_AGEMA_signal_26290 ;
    wire new_AGEMA_signal_26291 ;
    wire new_AGEMA_signal_26292 ;
    wire new_AGEMA_signal_26293 ;
    wire new_AGEMA_signal_26294 ;
    wire new_AGEMA_signal_26295 ;
    wire new_AGEMA_signal_26296 ;
    wire new_AGEMA_signal_26297 ;
    wire new_AGEMA_signal_26298 ;
    wire new_AGEMA_signal_26299 ;
    wire new_AGEMA_signal_26300 ;
    wire new_AGEMA_signal_26301 ;
    wire new_AGEMA_signal_26302 ;
    wire new_AGEMA_signal_26303 ;
    wire new_AGEMA_signal_26304 ;
    wire new_AGEMA_signal_26305 ;
    wire new_AGEMA_signal_26306 ;
    wire new_AGEMA_signal_26307 ;
    wire new_AGEMA_signal_26308 ;
    wire new_AGEMA_signal_26309 ;
    wire new_AGEMA_signal_26310 ;
    wire new_AGEMA_signal_26311 ;
    wire new_AGEMA_signal_26312 ;
    wire new_AGEMA_signal_26313 ;
    wire new_AGEMA_signal_26314 ;
    wire new_AGEMA_signal_26315 ;
    wire new_AGEMA_signal_26316 ;
    wire new_AGEMA_signal_26317 ;
    wire new_AGEMA_signal_26318 ;
    wire new_AGEMA_signal_26319 ;
    wire new_AGEMA_signal_26320 ;
    wire new_AGEMA_signal_26321 ;
    wire new_AGEMA_signal_26322 ;
    wire new_AGEMA_signal_26323 ;
    wire new_AGEMA_signal_26324 ;
    wire new_AGEMA_signal_26325 ;
    wire new_AGEMA_signal_26326 ;
    wire new_AGEMA_signal_26327 ;
    wire new_AGEMA_signal_26328 ;
    wire new_AGEMA_signal_26329 ;
    wire new_AGEMA_signal_26330 ;
    wire new_AGEMA_signal_26331 ;
    wire new_AGEMA_signal_26332 ;
    wire new_AGEMA_signal_26333 ;
    wire new_AGEMA_signal_26334 ;
    wire new_AGEMA_signal_26335 ;
    wire new_AGEMA_signal_26336 ;
    wire new_AGEMA_signal_26337 ;
    wire new_AGEMA_signal_26338 ;
    wire new_AGEMA_signal_26339 ;
    wire new_AGEMA_signal_26340 ;
    wire new_AGEMA_signal_26341 ;
    wire new_AGEMA_signal_26342 ;
    wire new_AGEMA_signal_26343 ;
    wire new_AGEMA_signal_26344 ;
    wire new_AGEMA_signal_26345 ;
    wire new_AGEMA_signal_26346 ;
    wire new_AGEMA_signal_26347 ;
    wire new_AGEMA_signal_26348 ;
    wire new_AGEMA_signal_26349 ;
    wire new_AGEMA_signal_26350 ;
    wire new_AGEMA_signal_26351 ;
    wire new_AGEMA_signal_26352 ;
    wire new_AGEMA_signal_26353 ;
    wire new_AGEMA_signal_26354 ;
    wire new_AGEMA_signal_26355 ;
    wire new_AGEMA_signal_26356 ;
    wire new_AGEMA_signal_26357 ;
    wire new_AGEMA_signal_26358 ;
    wire new_AGEMA_signal_26359 ;
    wire new_AGEMA_signal_26360 ;
    wire new_AGEMA_signal_26361 ;
    wire new_AGEMA_signal_26362 ;
    wire new_AGEMA_signal_26363 ;
    wire new_AGEMA_signal_26364 ;
    wire new_AGEMA_signal_26365 ;
    wire new_AGEMA_signal_26366 ;
    wire new_AGEMA_signal_26367 ;
    wire new_AGEMA_signal_26368 ;
    wire new_AGEMA_signal_26369 ;
    wire new_AGEMA_signal_26370 ;
    wire new_AGEMA_signal_26371 ;
    wire new_AGEMA_signal_26372 ;
    wire new_AGEMA_signal_26373 ;
    wire new_AGEMA_signal_26374 ;
    wire new_AGEMA_signal_26375 ;
    wire new_AGEMA_signal_26376 ;
    wire new_AGEMA_signal_26377 ;
    wire new_AGEMA_signal_26378 ;
    wire new_AGEMA_signal_26379 ;
    wire new_AGEMA_signal_26380 ;
    wire new_AGEMA_signal_26381 ;
    wire new_AGEMA_signal_26382 ;
    wire new_AGEMA_signal_26383 ;
    wire new_AGEMA_signal_26384 ;
    wire new_AGEMA_signal_26385 ;
    wire new_AGEMA_signal_26386 ;
    wire new_AGEMA_signal_26387 ;
    wire new_AGEMA_signal_26388 ;
    wire new_AGEMA_signal_26389 ;
    wire new_AGEMA_signal_26390 ;
    wire new_AGEMA_signal_26391 ;
    wire new_AGEMA_signal_26392 ;
    wire new_AGEMA_signal_26393 ;
    wire new_AGEMA_signal_26394 ;
    wire new_AGEMA_signal_26395 ;
    wire new_AGEMA_signal_26396 ;
    wire new_AGEMA_signal_26397 ;
    wire new_AGEMA_signal_26398 ;
    wire new_AGEMA_signal_26399 ;
    wire new_AGEMA_signal_26400 ;
    wire new_AGEMA_signal_26401 ;
    wire new_AGEMA_signal_26402 ;
    wire new_AGEMA_signal_26403 ;
    wire new_AGEMA_signal_26404 ;
    wire new_AGEMA_signal_26405 ;
    wire new_AGEMA_signal_26406 ;
    wire new_AGEMA_signal_26407 ;
    wire new_AGEMA_signal_26408 ;
    wire new_AGEMA_signal_26409 ;
    wire new_AGEMA_signal_26410 ;
    wire new_AGEMA_signal_26411 ;
    wire new_AGEMA_signal_26412 ;
    wire new_AGEMA_signal_26413 ;
    wire new_AGEMA_signal_26414 ;
    wire new_AGEMA_signal_26415 ;
    wire new_AGEMA_signal_26416 ;
    wire new_AGEMA_signal_26417 ;
    wire new_AGEMA_signal_26418 ;
    wire new_AGEMA_signal_26419 ;
    wire new_AGEMA_signal_26420 ;
    wire new_AGEMA_signal_26421 ;
    wire new_AGEMA_signal_26422 ;
    wire new_AGEMA_signal_26423 ;
    wire new_AGEMA_signal_26424 ;
    wire new_AGEMA_signal_26425 ;
    wire new_AGEMA_signal_26426 ;
    wire new_AGEMA_signal_26427 ;
    wire new_AGEMA_signal_26428 ;
    wire new_AGEMA_signal_26429 ;
    wire new_AGEMA_signal_26430 ;
    wire new_AGEMA_signal_26431 ;
    wire new_AGEMA_signal_26432 ;
    wire new_AGEMA_signal_26433 ;
    wire new_AGEMA_signal_26434 ;
    wire new_AGEMA_signal_26435 ;
    wire new_AGEMA_signal_26436 ;
    wire new_AGEMA_signal_26437 ;
    wire new_AGEMA_signal_26438 ;
    wire new_AGEMA_signal_26439 ;
    wire new_AGEMA_signal_26440 ;
    wire new_AGEMA_signal_26441 ;
    wire new_AGEMA_signal_26442 ;
    wire new_AGEMA_signal_26443 ;
    wire new_AGEMA_signal_26444 ;
    wire new_AGEMA_signal_26445 ;
    wire new_AGEMA_signal_26446 ;
    wire new_AGEMA_signal_26447 ;
    wire new_AGEMA_signal_26448 ;
    wire new_AGEMA_signal_26449 ;
    wire new_AGEMA_signal_26450 ;
    wire new_AGEMA_signal_26451 ;
    wire new_AGEMA_signal_26452 ;
    wire new_AGEMA_signal_26453 ;
    wire new_AGEMA_signal_26454 ;
    wire new_AGEMA_signal_26455 ;
    wire new_AGEMA_signal_26456 ;
    wire new_AGEMA_signal_26457 ;
    wire new_AGEMA_signal_26458 ;
    wire new_AGEMA_signal_26459 ;
    wire new_AGEMA_signal_26460 ;
    wire new_AGEMA_signal_26461 ;
    wire new_AGEMA_signal_26462 ;
    wire new_AGEMA_signal_26463 ;
    wire new_AGEMA_signal_26464 ;
    wire new_AGEMA_signal_26465 ;
    wire new_AGEMA_signal_26466 ;
    wire new_AGEMA_signal_26467 ;
    wire new_AGEMA_signal_26468 ;
    wire new_AGEMA_signal_26469 ;
    wire new_AGEMA_signal_26470 ;
    wire new_AGEMA_signal_26471 ;
    wire new_AGEMA_signal_26472 ;
    wire new_AGEMA_signal_26473 ;
    wire new_AGEMA_signal_26474 ;
    wire new_AGEMA_signal_26475 ;
    wire new_AGEMA_signal_26476 ;
    wire new_AGEMA_signal_26477 ;
    wire new_AGEMA_signal_26478 ;
    wire new_AGEMA_signal_26479 ;
    wire new_AGEMA_signal_26480 ;
    wire new_AGEMA_signal_26481 ;
    wire new_AGEMA_signal_26482 ;
    wire new_AGEMA_signal_26483 ;
    wire new_AGEMA_signal_26484 ;
    wire new_AGEMA_signal_26485 ;
    wire new_AGEMA_signal_26486 ;
    wire new_AGEMA_signal_26487 ;
    wire new_AGEMA_signal_26488 ;
    wire new_AGEMA_signal_26489 ;
    wire new_AGEMA_signal_26490 ;
    wire new_AGEMA_signal_26491 ;
    wire new_AGEMA_signal_26492 ;
    wire new_AGEMA_signal_26493 ;
    wire new_AGEMA_signal_26494 ;
    wire new_AGEMA_signal_26495 ;
    wire new_AGEMA_signal_26496 ;
    wire new_AGEMA_signal_26497 ;
    wire new_AGEMA_signal_26498 ;
    wire new_AGEMA_signal_26499 ;
    wire new_AGEMA_signal_26500 ;
    wire new_AGEMA_signal_26501 ;
    wire new_AGEMA_signal_26502 ;
    wire new_AGEMA_signal_26503 ;
    wire new_AGEMA_signal_26504 ;
    wire new_AGEMA_signal_26505 ;
    wire new_AGEMA_signal_26506 ;
    wire new_AGEMA_signal_26507 ;
    wire new_AGEMA_signal_26508 ;
    wire new_AGEMA_signal_26509 ;
    wire new_AGEMA_signal_26510 ;
    wire new_AGEMA_signal_26511 ;
    wire new_AGEMA_signal_26512 ;
    wire new_AGEMA_signal_26513 ;
    wire new_AGEMA_signal_26514 ;
    wire new_AGEMA_signal_26515 ;
    wire new_AGEMA_signal_26516 ;
    wire new_AGEMA_signal_26517 ;
    wire new_AGEMA_signal_26518 ;
    wire new_AGEMA_signal_26519 ;
    wire new_AGEMA_signal_26520 ;
    wire new_AGEMA_signal_26521 ;
    wire new_AGEMA_signal_26522 ;
    wire new_AGEMA_signal_26523 ;
    wire new_AGEMA_signal_26524 ;
    wire new_AGEMA_signal_26525 ;
    wire new_AGEMA_signal_26526 ;
    wire new_AGEMA_signal_26527 ;
    wire new_AGEMA_signal_26528 ;
    wire new_AGEMA_signal_26529 ;
    wire new_AGEMA_signal_26530 ;
    wire new_AGEMA_signal_26531 ;
    wire new_AGEMA_signal_26532 ;
    wire new_AGEMA_signal_26533 ;
    wire new_AGEMA_signal_26534 ;
    wire new_AGEMA_signal_26535 ;
    wire new_AGEMA_signal_26536 ;
    wire new_AGEMA_signal_26537 ;
    wire new_AGEMA_signal_26538 ;
    wire new_AGEMA_signal_26539 ;
    wire new_AGEMA_signal_26540 ;
    wire new_AGEMA_signal_26541 ;
    wire new_AGEMA_signal_26542 ;
    wire new_AGEMA_signal_26543 ;
    wire new_AGEMA_signal_26544 ;
    wire new_AGEMA_signal_26545 ;
    wire new_AGEMA_signal_26546 ;
    wire new_AGEMA_signal_26547 ;
    wire new_AGEMA_signal_26548 ;
    wire new_AGEMA_signal_26549 ;
    wire new_AGEMA_signal_26550 ;
    wire new_AGEMA_signal_26551 ;
    wire new_AGEMA_signal_26552 ;
    wire new_AGEMA_signal_26553 ;
    wire new_AGEMA_signal_26554 ;
    wire new_AGEMA_signal_26555 ;
    wire new_AGEMA_signal_26556 ;
    wire new_AGEMA_signal_26557 ;
    wire new_AGEMA_signal_26558 ;
    wire new_AGEMA_signal_26559 ;
    wire new_AGEMA_signal_26560 ;
    wire new_AGEMA_signal_26561 ;
    wire new_AGEMA_signal_26562 ;
    wire new_AGEMA_signal_26563 ;
    wire new_AGEMA_signal_26564 ;
    wire new_AGEMA_signal_26565 ;
    wire new_AGEMA_signal_26566 ;
    wire new_AGEMA_signal_26567 ;
    wire new_AGEMA_signal_26568 ;
    wire new_AGEMA_signal_26569 ;
    wire new_AGEMA_signal_26570 ;
    wire new_AGEMA_signal_26571 ;
    wire new_AGEMA_signal_26572 ;
    wire new_AGEMA_signal_26573 ;
    wire new_AGEMA_signal_26574 ;
    wire new_AGEMA_signal_26575 ;
    wire new_AGEMA_signal_26576 ;
    wire new_AGEMA_signal_26577 ;
    wire new_AGEMA_signal_26578 ;
    wire new_AGEMA_signal_26579 ;
    wire new_AGEMA_signal_26580 ;
    wire new_AGEMA_signal_26581 ;
    wire new_AGEMA_signal_26582 ;
    wire new_AGEMA_signal_26583 ;
    wire new_AGEMA_signal_26584 ;
    wire new_AGEMA_signal_26585 ;
    wire new_AGEMA_signal_26586 ;
    wire new_AGEMA_signal_26587 ;
    wire new_AGEMA_signal_26588 ;
    wire new_AGEMA_signal_26589 ;
    wire new_AGEMA_signal_26590 ;
    wire new_AGEMA_signal_26591 ;
    wire new_AGEMA_signal_26592 ;
    wire new_AGEMA_signal_26593 ;
    wire new_AGEMA_signal_26594 ;
    wire new_AGEMA_signal_26595 ;
    wire new_AGEMA_signal_26596 ;
    wire new_AGEMA_signal_26597 ;
    wire new_AGEMA_signal_26598 ;
    wire new_AGEMA_signal_26599 ;
    wire new_AGEMA_signal_26600 ;
    wire new_AGEMA_signal_26601 ;
    wire new_AGEMA_signal_26602 ;
    wire new_AGEMA_signal_26603 ;
    wire new_AGEMA_signal_26604 ;
    wire new_AGEMA_signal_26605 ;
    wire new_AGEMA_signal_26606 ;
    wire new_AGEMA_signal_26607 ;
    wire new_AGEMA_signal_26608 ;
    wire new_AGEMA_signal_26609 ;
    wire new_AGEMA_signal_26610 ;
    wire new_AGEMA_signal_26611 ;
    wire new_AGEMA_signal_26612 ;
    wire new_AGEMA_signal_26613 ;
    wire new_AGEMA_signal_26614 ;
    wire new_AGEMA_signal_26615 ;
    wire new_AGEMA_signal_26616 ;
    wire new_AGEMA_signal_26617 ;
    wire new_AGEMA_signal_26618 ;
    wire new_AGEMA_signal_26619 ;
    wire new_AGEMA_signal_26620 ;
    wire new_AGEMA_signal_26621 ;
    wire new_AGEMA_signal_26622 ;
    wire new_AGEMA_signal_26623 ;
    wire new_AGEMA_signal_26624 ;
    wire new_AGEMA_signal_26625 ;
    wire new_AGEMA_signal_26626 ;
    wire new_AGEMA_signal_26627 ;
    wire new_AGEMA_signal_26628 ;
    wire new_AGEMA_signal_26629 ;
    wire new_AGEMA_signal_26630 ;
    wire new_AGEMA_signal_26631 ;
    wire new_AGEMA_signal_26632 ;
    wire new_AGEMA_signal_26633 ;
    wire new_AGEMA_signal_26634 ;
    wire new_AGEMA_signal_26635 ;
    wire new_AGEMA_signal_26636 ;
    wire new_AGEMA_signal_26637 ;
    wire new_AGEMA_signal_26638 ;
    wire new_AGEMA_signal_26639 ;
    wire new_AGEMA_signal_26640 ;
    wire new_AGEMA_signal_26641 ;
    wire new_AGEMA_signal_26642 ;
    wire new_AGEMA_signal_26643 ;
    wire new_AGEMA_signal_26644 ;
    wire new_AGEMA_signal_26645 ;
    wire new_AGEMA_signal_26646 ;
    wire new_AGEMA_signal_26647 ;
    wire new_AGEMA_signal_26648 ;
    wire new_AGEMA_signal_26649 ;
    wire new_AGEMA_signal_26650 ;
    wire new_AGEMA_signal_26651 ;
    wire new_AGEMA_signal_26652 ;
    wire new_AGEMA_signal_26653 ;
    wire new_AGEMA_signal_26654 ;
    wire new_AGEMA_signal_26655 ;
    wire new_AGEMA_signal_26656 ;
    wire new_AGEMA_signal_26657 ;
    wire new_AGEMA_signal_26658 ;
    wire new_AGEMA_signal_26659 ;
    wire new_AGEMA_signal_26660 ;
    wire new_AGEMA_signal_26661 ;
    wire new_AGEMA_signal_26662 ;
    wire new_AGEMA_signal_26663 ;
    wire new_AGEMA_signal_26664 ;
    wire new_AGEMA_signal_26665 ;
    wire new_AGEMA_signal_26666 ;
    wire new_AGEMA_signal_26667 ;
    wire new_AGEMA_signal_26668 ;
    wire new_AGEMA_signal_26669 ;
    wire new_AGEMA_signal_26670 ;
    wire new_AGEMA_signal_26671 ;
    wire new_AGEMA_signal_26672 ;
    wire new_AGEMA_signal_26673 ;
    wire new_AGEMA_signal_26674 ;
    wire new_AGEMA_signal_26675 ;
    wire new_AGEMA_signal_26676 ;
    wire new_AGEMA_signal_26677 ;
    wire new_AGEMA_signal_26678 ;
    wire new_AGEMA_signal_26679 ;
    wire new_AGEMA_signal_26680 ;
    wire new_AGEMA_signal_26681 ;
    wire new_AGEMA_signal_26682 ;
    wire new_AGEMA_signal_26683 ;
    wire new_AGEMA_signal_26684 ;
    wire new_AGEMA_signal_26685 ;
    wire new_AGEMA_signal_26686 ;
    wire new_AGEMA_signal_26687 ;
    wire new_AGEMA_signal_26688 ;
    wire new_AGEMA_signal_26689 ;
    wire new_AGEMA_signal_26690 ;
    wire new_AGEMA_signal_26691 ;
    wire new_AGEMA_signal_26692 ;
    wire new_AGEMA_signal_26693 ;
    wire new_AGEMA_signal_26694 ;
    wire new_AGEMA_signal_26695 ;
    wire new_AGEMA_signal_26696 ;
    wire new_AGEMA_signal_26697 ;
    wire new_AGEMA_signal_26698 ;
    wire new_AGEMA_signal_26699 ;
    wire new_AGEMA_signal_26700 ;
    wire new_AGEMA_signal_26701 ;
    wire new_AGEMA_signal_26702 ;
    wire new_AGEMA_signal_26703 ;
    wire new_AGEMA_signal_26704 ;
    wire new_AGEMA_signal_26705 ;
    wire new_AGEMA_signal_26706 ;
    wire new_AGEMA_signal_26707 ;
    wire new_AGEMA_signal_26708 ;
    wire new_AGEMA_signal_26709 ;
    wire new_AGEMA_signal_26710 ;
    wire new_AGEMA_signal_26711 ;
    wire new_AGEMA_signal_26712 ;
    wire new_AGEMA_signal_26713 ;
    wire new_AGEMA_signal_26714 ;
    wire new_AGEMA_signal_26715 ;
    wire new_AGEMA_signal_26716 ;
    wire new_AGEMA_signal_26717 ;
    wire new_AGEMA_signal_26718 ;
    wire new_AGEMA_signal_26719 ;
    wire new_AGEMA_signal_26720 ;
    wire new_AGEMA_signal_26721 ;
    wire new_AGEMA_signal_26722 ;
    wire new_AGEMA_signal_26723 ;
    wire new_AGEMA_signal_26724 ;
    wire new_AGEMA_signal_26725 ;
    wire new_AGEMA_signal_26726 ;
    wire new_AGEMA_signal_26727 ;
    wire new_AGEMA_signal_26728 ;
    wire new_AGEMA_signal_26729 ;
    wire new_AGEMA_signal_26730 ;
    wire new_AGEMA_signal_26731 ;
    wire new_AGEMA_signal_26732 ;
    wire new_AGEMA_signal_26733 ;
    wire new_AGEMA_signal_26734 ;
    wire new_AGEMA_signal_26735 ;
    wire new_AGEMA_signal_26736 ;
    wire new_AGEMA_signal_26737 ;
    wire new_AGEMA_signal_26738 ;
    wire new_AGEMA_signal_26739 ;
    wire new_AGEMA_signal_26740 ;
    wire new_AGEMA_signal_26741 ;
    wire new_AGEMA_signal_26742 ;
    wire new_AGEMA_signal_26743 ;
    wire new_AGEMA_signal_26744 ;
    wire new_AGEMA_signal_26745 ;
    wire new_AGEMA_signal_26746 ;
    wire new_AGEMA_signal_26747 ;
    wire new_AGEMA_signal_26748 ;
    wire new_AGEMA_signal_26749 ;
    wire new_AGEMA_signal_26750 ;
    wire new_AGEMA_signal_26751 ;
    wire new_AGEMA_signal_26752 ;
    wire new_AGEMA_signal_26753 ;
    wire new_AGEMA_signal_26754 ;
    wire new_AGEMA_signal_26755 ;
    wire new_AGEMA_signal_26756 ;
    wire new_AGEMA_signal_26757 ;
    wire new_AGEMA_signal_26758 ;
    wire new_AGEMA_signal_26759 ;
    wire new_AGEMA_signal_26760 ;
    wire new_AGEMA_signal_26761 ;
    wire new_AGEMA_signal_26762 ;
    wire new_AGEMA_signal_26763 ;
    wire new_AGEMA_signal_26764 ;
    wire new_AGEMA_signal_26765 ;
    wire new_AGEMA_signal_26766 ;
    wire new_AGEMA_signal_26767 ;
    wire new_AGEMA_signal_26768 ;
    wire new_AGEMA_signal_26769 ;
    wire new_AGEMA_signal_26770 ;
    wire new_AGEMA_signal_26771 ;
    wire new_AGEMA_signal_26772 ;
    wire new_AGEMA_signal_26773 ;
    wire new_AGEMA_signal_26774 ;
    wire new_AGEMA_signal_26775 ;
    wire new_AGEMA_signal_26776 ;
    wire new_AGEMA_signal_26777 ;
    wire new_AGEMA_signal_26778 ;
    wire new_AGEMA_signal_26779 ;
    wire new_AGEMA_signal_26780 ;
    wire new_AGEMA_signal_26781 ;
    wire new_AGEMA_signal_26782 ;
    wire new_AGEMA_signal_26783 ;
    wire new_AGEMA_signal_26784 ;
    wire new_AGEMA_signal_26785 ;
    wire new_AGEMA_signal_26786 ;
    wire new_AGEMA_signal_26787 ;
    wire new_AGEMA_signal_26788 ;
    wire new_AGEMA_signal_26789 ;
    wire new_AGEMA_signal_26790 ;
    wire new_AGEMA_signal_26791 ;
    wire new_AGEMA_signal_26792 ;
    wire new_AGEMA_signal_26793 ;
    wire new_AGEMA_signal_26794 ;
    wire new_AGEMA_signal_26795 ;
    wire new_AGEMA_signal_26796 ;
    wire new_AGEMA_signal_26797 ;
    wire new_AGEMA_signal_26798 ;
    wire new_AGEMA_signal_26799 ;
    wire new_AGEMA_signal_26800 ;
    wire new_AGEMA_signal_26801 ;
    wire new_AGEMA_signal_26802 ;
    wire new_AGEMA_signal_26803 ;
    wire new_AGEMA_signal_26804 ;
    wire new_AGEMA_signal_26805 ;
    wire new_AGEMA_signal_26806 ;
    wire new_AGEMA_signal_26807 ;
    wire new_AGEMA_signal_26808 ;
    wire new_AGEMA_signal_26809 ;
    wire new_AGEMA_signal_26810 ;
    wire new_AGEMA_signal_26811 ;
    wire new_AGEMA_signal_26812 ;
    wire new_AGEMA_signal_26813 ;
    wire new_AGEMA_signal_26814 ;
    wire new_AGEMA_signal_26815 ;
    wire new_AGEMA_signal_26816 ;
    wire new_AGEMA_signal_26817 ;
    wire new_AGEMA_signal_26818 ;
    wire new_AGEMA_signal_26819 ;
    wire new_AGEMA_signal_26820 ;
    wire new_AGEMA_signal_26821 ;
    wire new_AGEMA_signal_26822 ;
    wire new_AGEMA_signal_26823 ;
    wire new_AGEMA_signal_26824 ;
    wire new_AGEMA_signal_26825 ;
    wire new_AGEMA_signal_26826 ;
    wire new_AGEMA_signal_26827 ;
    wire new_AGEMA_signal_26828 ;
    wire new_AGEMA_signal_26829 ;
    wire new_AGEMA_signal_26830 ;
    wire new_AGEMA_signal_26831 ;
    wire new_AGEMA_signal_26832 ;
    wire new_AGEMA_signal_26833 ;
    wire new_AGEMA_signal_26834 ;
    wire new_AGEMA_signal_26835 ;
    wire new_AGEMA_signal_26836 ;
    wire new_AGEMA_signal_26837 ;
    wire new_AGEMA_signal_26838 ;
    wire new_AGEMA_signal_26839 ;
    wire new_AGEMA_signal_26840 ;
    wire new_AGEMA_signal_26841 ;
    wire new_AGEMA_signal_26842 ;
    wire new_AGEMA_signal_26843 ;
    wire new_AGEMA_signal_26844 ;
    wire new_AGEMA_signal_26845 ;
    wire new_AGEMA_signal_26846 ;
    wire new_AGEMA_signal_26847 ;
    wire new_AGEMA_signal_26848 ;
    wire new_AGEMA_signal_26849 ;
    wire new_AGEMA_signal_26850 ;
    wire new_AGEMA_signal_26851 ;
    wire new_AGEMA_signal_26852 ;
    wire new_AGEMA_signal_26853 ;
    wire new_AGEMA_signal_26854 ;
    wire new_AGEMA_signal_26855 ;
    wire new_AGEMA_signal_26856 ;
    wire new_AGEMA_signal_26857 ;
    wire new_AGEMA_signal_26858 ;
    wire new_AGEMA_signal_26859 ;
    wire new_AGEMA_signal_26860 ;
    wire new_AGEMA_signal_26861 ;
    wire new_AGEMA_signal_26862 ;
    wire new_AGEMA_signal_26863 ;
    wire new_AGEMA_signal_26864 ;
    wire new_AGEMA_signal_26865 ;
    wire new_AGEMA_signal_26866 ;
    wire new_AGEMA_signal_26867 ;
    wire new_AGEMA_signal_26868 ;
    wire new_AGEMA_signal_26869 ;
    wire new_AGEMA_signal_26870 ;
    wire new_AGEMA_signal_26871 ;
    wire new_AGEMA_signal_26872 ;
    wire new_AGEMA_signal_26873 ;
    wire new_AGEMA_signal_26874 ;
    wire new_AGEMA_signal_26875 ;
    wire new_AGEMA_signal_26876 ;
    wire new_AGEMA_signal_26877 ;
    wire new_AGEMA_signal_26878 ;
    wire new_AGEMA_signal_26879 ;
    wire new_AGEMA_signal_26880 ;
    wire new_AGEMA_signal_26881 ;
    wire new_AGEMA_signal_26882 ;
    wire new_AGEMA_signal_26883 ;
    wire new_AGEMA_signal_26884 ;
    wire new_AGEMA_signal_26885 ;
    wire new_AGEMA_signal_26886 ;
    wire new_AGEMA_signal_26887 ;
    wire new_AGEMA_signal_26888 ;
    wire new_AGEMA_signal_26889 ;
    wire new_AGEMA_signal_26890 ;
    wire new_AGEMA_signal_26891 ;
    wire new_AGEMA_signal_26892 ;
    wire new_AGEMA_signal_26893 ;
    wire new_AGEMA_signal_26894 ;
    wire new_AGEMA_signal_26895 ;
    wire new_AGEMA_signal_26896 ;
    wire new_AGEMA_signal_26897 ;
    wire new_AGEMA_signal_26898 ;
    wire new_AGEMA_signal_26899 ;
    wire new_AGEMA_signal_26900 ;
    wire new_AGEMA_signal_26901 ;
    wire new_AGEMA_signal_26902 ;
    wire new_AGEMA_signal_26903 ;
    wire new_AGEMA_signal_26904 ;
    wire new_AGEMA_signal_26905 ;
    wire new_AGEMA_signal_26906 ;
    wire new_AGEMA_signal_26907 ;
    wire new_AGEMA_signal_26908 ;
    wire new_AGEMA_signal_26909 ;
    wire new_AGEMA_signal_26910 ;
    wire new_AGEMA_signal_26911 ;
    wire new_AGEMA_signal_26912 ;
    wire new_AGEMA_signal_26913 ;
    wire new_AGEMA_signal_26914 ;
    wire new_AGEMA_signal_26915 ;
    wire new_AGEMA_signal_26916 ;
    wire new_AGEMA_signal_26917 ;
    wire new_AGEMA_signal_26918 ;
    wire new_AGEMA_signal_26919 ;
    wire new_AGEMA_signal_26920 ;
    wire new_AGEMA_signal_26921 ;
    wire new_AGEMA_signal_26922 ;
    wire new_AGEMA_signal_26923 ;
    wire new_AGEMA_signal_26924 ;
    wire new_AGEMA_signal_26925 ;
    wire new_AGEMA_signal_26926 ;
    wire new_AGEMA_signal_26927 ;
    wire new_AGEMA_signal_26928 ;
    wire new_AGEMA_signal_26929 ;
    wire new_AGEMA_signal_26930 ;
    wire new_AGEMA_signal_26931 ;
    wire new_AGEMA_signal_26932 ;
    wire new_AGEMA_signal_26933 ;
    wire new_AGEMA_signal_26934 ;
    wire new_AGEMA_signal_26935 ;
    wire new_AGEMA_signal_26936 ;
    wire new_AGEMA_signal_26937 ;
    wire new_AGEMA_signal_26938 ;
    wire new_AGEMA_signal_26939 ;
    wire new_AGEMA_signal_26940 ;
    wire new_AGEMA_signal_26941 ;
    wire new_AGEMA_signal_26942 ;
    wire new_AGEMA_signal_26943 ;
    wire new_AGEMA_signal_26944 ;
    wire new_AGEMA_signal_26945 ;
    wire new_AGEMA_signal_26946 ;
    wire new_AGEMA_signal_26947 ;
    wire new_AGEMA_signal_26948 ;
    wire new_AGEMA_signal_26949 ;
    wire new_AGEMA_signal_26950 ;
    wire new_AGEMA_signal_26951 ;
    wire new_AGEMA_signal_26952 ;
    wire new_AGEMA_signal_26953 ;
    wire new_AGEMA_signal_26954 ;
    wire new_AGEMA_signal_26955 ;
    wire new_AGEMA_signal_26956 ;
    wire new_AGEMA_signal_26957 ;
    wire new_AGEMA_signal_26958 ;
    wire new_AGEMA_signal_26959 ;
    wire new_AGEMA_signal_26960 ;
    wire new_AGEMA_signal_26961 ;
    wire new_AGEMA_signal_26962 ;
    wire new_AGEMA_signal_26963 ;
    wire new_AGEMA_signal_26964 ;
    wire new_AGEMA_signal_26965 ;
    wire new_AGEMA_signal_26966 ;
    wire new_AGEMA_signal_26967 ;
    wire new_AGEMA_signal_26968 ;
    wire new_AGEMA_signal_26969 ;
    wire new_AGEMA_signal_26970 ;
    wire new_AGEMA_signal_26971 ;
    wire new_AGEMA_signal_26972 ;
    wire new_AGEMA_signal_26973 ;
    wire new_AGEMA_signal_26974 ;
    wire new_AGEMA_signal_26975 ;
    wire new_AGEMA_signal_26976 ;
    wire new_AGEMA_signal_26977 ;
    wire new_AGEMA_signal_26978 ;
    wire new_AGEMA_signal_26979 ;
    wire new_AGEMA_signal_26980 ;
    wire new_AGEMA_signal_26981 ;
    wire new_AGEMA_signal_26982 ;
    wire new_AGEMA_signal_26983 ;
    wire new_AGEMA_signal_26984 ;
    wire new_AGEMA_signal_26985 ;
    wire new_AGEMA_signal_26986 ;
    wire new_AGEMA_signal_26987 ;
    wire new_AGEMA_signal_26988 ;
    wire new_AGEMA_signal_26989 ;
    wire new_AGEMA_signal_26990 ;
    wire new_AGEMA_signal_26991 ;
    wire new_AGEMA_signal_26992 ;
    wire new_AGEMA_signal_26993 ;
    wire new_AGEMA_signal_26994 ;
    wire new_AGEMA_signal_26995 ;
    wire new_AGEMA_signal_26996 ;
    wire new_AGEMA_signal_26997 ;
    wire new_AGEMA_signal_26998 ;
    wire new_AGEMA_signal_26999 ;
    wire new_AGEMA_signal_27000 ;
    wire new_AGEMA_signal_27001 ;
    wire new_AGEMA_signal_27002 ;
    wire new_AGEMA_signal_27003 ;
    wire new_AGEMA_signal_27004 ;
    wire new_AGEMA_signal_27005 ;
    wire new_AGEMA_signal_27006 ;
    wire new_AGEMA_signal_27007 ;
    wire new_AGEMA_signal_27008 ;
    wire new_AGEMA_signal_27009 ;
    wire new_AGEMA_signal_27010 ;
    wire new_AGEMA_signal_27011 ;
    wire new_AGEMA_signal_27012 ;
    wire new_AGEMA_signal_27013 ;
    wire new_AGEMA_signal_27014 ;
    wire new_AGEMA_signal_27015 ;
    wire new_AGEMA_signal_27016 ;
    wire new_AGEMA_signal_27017 ;
    wire new_AGEMA_signal_27018 ;
    wire new_AGEMA_signal_27019 ;
    wire new_AGEMA_signal_27020 ;
    wire new_AGEMA_signal_27021 ;
    wire new_AGEMA_signal_27022 ;
    wire new_AGEMA_signal_27023 ;
    wire new_AGEMA_signal_27024 ;
    wire new_AGEMA_signal_27025 ;
    wire new_AGEMA_signal_27026 ;
    wire new_AGEMA_signal_27027 ;
    wire new_AGEMA_signal_27028 ;
    wire new_AGEMA_signal_27029 ;
    wire new_AGEMA_signal_27030 ;
    wire new_AGEMA_signal_27031 ;
    wire new_AGEMA_signal_27032 ;
    wire new_AGEMA_signal_27033 ;
    wire new_AGEMA_signal_27034 ;
    wire new_AGEMA_signal_27035 ;
    wire new_AGEMA_signal_27036 ;
    wire new_AGEMA_signal_27037 ;
    wire new_AGEMA_signal_27038 ;
    wire new_AGEMA_signal_27039 ;
    wire new_AGEMA_signal_27040 ;
    wire new_AGEMA_signal_27041 ;
    wire new_AGEMA_signal_27042 ;
    wire new_AGEMA_signal_27043 ;
    wire new_AGEMA_signal_27044 ;
    wire new_AGEMA_signal_27045 ;
    wire new_AGEMA_signal_27046 ;
    wire new_AGEMA_signal_27047 ;
    wire new_AGEMA_signal_27048 ;
    wire new_AGEMA_signal_27049 ;
    wire new_AGEMA_signal_27050 ;
    wire new_AGEMA_signal_27051 ;
    wire new_AGEMA_signal_27052 ;
    wire new_AGEMA_signal_27053 ;
    wire new_AGEMA_signal_27054 ;
    wire new_AGEMA_signal_27055 ;
    wire new_AGEMA_signal_27056 ;
    wire new_AGEMA_signal_27057 ;
    wire new_AGEMA_signal_27058 ;
    wire new_AGEMA_signal_27059 ;
    wire new_AGEMA_signal_27060 ;
    wire new_AGEMA_signal_27061 ;
    wire new_AGEMA_signal_27062 ;
    wire new_AGEMA_signal_27063 ;
    wire new_AGEMA_signal_27064 ;
    wire new_AGEMA_signal_27065 ;
    wire new_AGEMA_signal_27066 ;
    wire new_AGEMA_signal_27067 ;
    wire new_AGEMA_signal_27068 ;
    wire new_AGEMA_signal_27069 ;
    wire new_AGEMA_signal_27070 ;
    wire new_AGEMA_signal_27071 ;
    wire new_AGEMA_signal_27072 ;
    wire new_AGEMA_signal_27073 ;
    wire new_AGEMA_signal_27074 ;
    wire new_AGEMA_signal_27075 ;
    wire new_AGEMA_signal_27076 ;
    wire new_AGEMA_signal_27077 ;
    wire new_AGEMA_signal_27078 ;
    wire new_AGEMA_signal_27079 ;
    wire new_AGEMA_signal_27080 ;
    wire new_AGEMA_signal_27081 ;
    wire new_AGEMA_signal_27082 ;
    wire new_AGEMA_signal_27083 ;
    wire new_AGEMA_signal_27084 ;
    wire new_AGEMA_signal_27085 ;
    wire new_AGEMA_signal_27086 ;
    wire new_AGEMA_signal_27087 ;
    wire new_AGEMA_signal_27088 ;
    wire new_AGEMA_signal_27089 ;
    wire new_AGEMA_signal_27090 ;
    wire new_AGEMA_signal_27091 ;
    wire new_AGEMA_signal_27092 ;
    wire new_AGEMA_signal_27093 ;
    wire new_AGEMA_signal_27094 ;
    wire new_AGEMA_signal_27095 ;
    wire new_AGEMA_signal_27096 ;
    wire new_AGEMA_signal_27097 ;
    wire new_AGEMA_signal_27098 ;
    wire new_AGEMA_signal_27099 ;
    wire new_AGEMA_signal_27100 ;
    wire new_AGEMA_signal_27101 ;
    wire new_AGEMA_signal_27102 ;
    wire new_AGEMA_signal_27103 ;
    wire new_AGEMA_signal_27104 ;
    wire new_AGEMA_signal_27105 ;
    wire new_AGEMA_signal_27106 ;
    wire new_AGEMA_signal_27107 ;
    wire new_AGEMA_signal_27108 ;
    wire new_AGEMA_signal_27109 ;
    wire new_AGEMA_signal_27110 ;
    wire new_AGEMA_signal_27111 ;
    wire new_AGEMA_signal_27112 ;
    wire new_AGEMA_signal_27113 ;
    wire new_AGEMA_signal_27114 ;
    wire new_AGEMA_signal_27115 ;
    wire new_AGEMA_signal_27116 ;
    wire new_AGEMA_signal_27117 ;
    wire new_AGEMA_signal_27118 ;
    wire new_AGEMA_signal_27119 ;
    wire new_AGEMA_signal_27120 ;
    wire new_AGEMA_signal_27121 ;
    wire new_AGEMA_signal_27122 ;
    wire new_AGEMA_signal_27123 ;
    wire new_AGEMA_signal_27124 ;
    wire new_AGEMA_signal_27125 ;
    wire new_AGEMA_signal_27126 ;
    wire new_AGEMA_signal_27127 ;
    wire new_AGEMA_signal_27128 ;
    wire new_AGEMA_signal_27129 ;
    wire new_AGEMA_signal_27130 ;
    wire new_AGEMA_signal_27131 ;
    wire new_AGEMA_signal_27132 ;
    wire new_AGEMA_signal_27133 ;
    wire new_AGEMA_signal_27134 ;
    wire new_AGEMA_signal_27135 ;
    wire new_AGEMA_signal_27136 ;
    wire new_AGEMA_signal_27137 ;
    wire new_AGEMA_signal_27138 ;
    wire new_AGEMA_signal_27139 ;
    wire new_AGEMA_signal_27140 ;
    wire new_AGEMA_signal_27141 ;
    wire new_AGEMA_signal_27142 ;
    wire new_AGEMA_signal_27143 ;
    wire new_AGEMA_signal_27144 ;
    wire new_AGEMA_signal_27145 ;
    wire new_AGEMA_signal_27146 ;
    wire new_AGEMA_signal_27147 ;
    wire new_AGEMA_signal_27148 ;
    wire new_AGEMA_signal_27149 ;
    wire new_AGEMA_signal_27150 ;
    wire new_AGEMA_signal_27151 ;
    wire new_AGEMA_signal_27152 ;
    wire new_AGEMA_signal_27153 ;
    wire new_AGEMA_signal_27154 ;
    wire new_AGEMA_signal_27155 ;
    wire new_AGEMA_signal_27156 ;
    wire new_AGEMA_signal_27157 ;
    wire new_AGEMA_signal_27158 ;
    wire new_AGEMA_signal_27159 ;
    wire new_AGEMA_signal_27160 ;
    wire new_AGEMA_signal_27161 ;
    wire new_AGEMA_signal_27162 ;
    wire new_AGEMA_signal_27163 ;
    wire new_AGEMA_signal_27164 ;
    wire new_AGEMA_signal_27165 ;
    wire new_AGEMA_signal_27166 ;
    wire new_AGEMA_signal_27167 ;
    wire new_AGEMA_signal_27168 ;
    wire new_AGEMA_signal_27169 ;
    wire new_AGEMA_signal_27170 ;
    wire new_AGEMA_signal_27171 ;
    wire new_AGEMA_signal_27172 ;
    wire new_AGEMA_signal_27173 ;
    wire new_AGEMA_signal_27174 ;
    wire new_AGEMA_signal_27175 ;
    wire new_AGEMA_signal_27176 ;
    wire new_AGEMA_signal_27177 ;
    wire new_AGEMA_signal_27178 ;
    wire new_AGEMA_signal_27179 ;
    wire new_AGEMA_signal_27180 ;
    wire new_AGEMA_signal_27181 ;
    wire new_AGEMA_signal_27182 ;
    wire new_AGEMA_signal_27183 ;
    wire new_AGEMA_signal_27184 ;
    wire new_AGEMA_signal_27185 ;
    wire new_AGEMA_signal_27186 ;
    wire new_AGEMA_signal_27187 ;
    wire new_AGEMA_signal_27188 ;
    wire new_AGEMA_signal_27189 ;
    wire new_AGEMA_signal_27190 ;
    wire new_AGEMA_signal_27191 ;
    wire new_AGEMA_signal_27192 ;
    wire new_AGEMA_signal_27193 ;
    wire new_AGEMA_signal_27194 ;
    wire new_AGEMA_signal_27195 ;
    wire new_AGEMA_signal_27196 ;
    wire new_AGEMA_signal_27197 ;
    wire new_AGEMA_signal_27198 ;
    wire new_AGEMA_signal_27199 ;
    wire new_AGEMA_signal_27200 ;
    wire new_AGEMA_signal_27201 ;
    wire new_AGEMA_signal_27202 ;
    wire new_AGEMA_signal_27203 ;
    wire new_AGEMA_signal_27204 ;
    wire new_AGEMA_signal_27205 ;
    wire new_AGEMA_signal_27206 ;
    wire new_AGEMA_signal_27207 ;
    wire new_AGEMA_signal_27208 ;
    wire new_AGEMA_signal_27209 ;
    wire new_AGEMA_signal_27210 ;
    wire new_AGEMA_signal_27211 ;
    wire new_AGEMA_signal_27212 ;
    wire new_AGEMA_signal_27213 ;
    wire new_AGEMA_signal_27214 ;
    wire new_AGEMA_signal_27215 ;
    wire new_AGEMA_signal_27216 ;
    wire new_AGEMA_signal_27217 ;
    wire new_AGEMA_signal_27218 ;
    wire new_AGEMA_signal_27219 ;
    wire new_AGEMA_signal_27220 ;
    wire new_AGEMA_signal_27221 ;
    wire new_AGEMA_signal_27222 ;
    wire new_AGEMA_signal_27223 ;
    wire new_AGEMA_signal_27224 ;
    wire new_AGEMA_signal_27225 ;
    wire new_AGEMA_signal_27226 ;
    wire new_AGEMA_signal_27227 ;
    wire new_AGEMA_signal_27228 ;
    wire new_AGEMA_signal_27229 ;
    wire new_AGEMA_signal_27230 ;
    wire new_AGEMA_signal_27231 ;
    wire new_AGEMA_signal_27232 ;
    wire new_AGEMA_signal_27233 ;
    wire new_AGEMA_signal_27234 ;
    wire new_AGEMA_signal_27235 ;
    wire new_AGEMA_signal_27236 ;
    wire new_AGEMA_signal_27237 ;
    wire new_AGEMA_signal_27238 ;
    wire new_AGEMA_signal_27239 ;
    wire new_AGEMA_signal_27240 ;
    wire new_AGEMA_signal_27241 ;
    wire new_AGEMA_signal_27242 ;
    wire new_AGEMA_signal_27243 ;
    wire new_AGEMA_signal_27244 ;
    wire new_AGEMA_signal_27245 ;
    wire new_AGEMA_signal_27246 ;
    wire new_AGEMA_signal_27247 ;
    wire new_AGEMA_signal_27248 ;
    wire new_AGEMA_signal_27249 ;
    wire new_AGEMA_signal_27250 ;
    wire new_AGEMA_signal_27251 ;
    wire new_AGEMA_signal_27252 ;
    wire new_AGEMA_signal_27253 ;
    wire new_AGEMA_signal_27254 ;
    wire new_AGEMA_signal_27255 ;
    wire new_AGEMA_signal_27256 ;
    wire new_AGEMA_signal_27257 ;
    wire new_AGEMA_signal_27258 ;
    wire new_AGEMA_signal_27259 ;
    wire new_AGEMA_signal_27260 ;
    wire new_AGEMA_signal_27261 ;
    wire new_AGEMA_signal_27262 ;
    wire new_AGEMA_signal_27263 ;
    wire new_AGEMA_signal_27264 ;
    wire new_AGEMA_signal_27265 ;
    wire new_AGEMA_signal_27266 ;
    wire new_AGEMA_signal_27267 ;
    wire new_AGEMA_signal_27268 ;
    wire new_AGEMA_signal_27269 ;
    wire new_AGEMA_signal_27270 ;
    wire new_AGEMA_signal_27271 ;
    wire new_AGEMA_signal_27272 ;
    wire new_AGEMA_signal_27273 ;
    wire new_AGEMA_signal_27274 ;
    wire new_AGEMA_signal_27275 ;
    wire new_AGEMA_signal_27276 ;
    wire new_AGEMA_signal_27277 ;
    wire new_AGEMA_signal_27278 ;
    wire new_AGEMA_signal_27279 ;
    wire new_AGEMA_signal_27280 ;
    wire new_AGEMA_signal_27281 ;
    wire new_AGEMA_signal_27282 ;
    wire new_AGEMA_signal_27283 ;
    wire new_AGEMA_signal_27284 ;
    wire new_AGEMA_signal_27285 ;
    wire new_AGEMA_signal_27286 ;
    wire new_AGEMA_signal_27287 ;
    wire new_AGEMA_signal_27288 ;
    wire new_AGEMA_signal_27289 ;
    wire new_AGEMA_signal_27290 ;
    wire new_AGEMA_signal_27291 ;
    wire new_AGEMA_signal_27292 ;
    wire new_AGEMA_signal_27293 ;
    wire new_AGEMA_signal_27294 ;
    wire new_AGEMA_signal_27295 ;
    wire new_AGEMA_signal_27296 ;
    wire new_AGEMA_signal_27297 ;
    wire new_AGEMA_signal_27298 ;
    wire new_AGEMA_signal_27299 ;
    wire new_AGEMA_signal_27300 ;
    wire new_AGEMA_signal_27301 ;
    wire new_AGEMA_signal_27302 ;
    wire new_AGEMA_signal_27303 ;
    wire new_AGEMA_signal_27304 ;
    wire new_AGEMA_signal_27305 ;
    wire new_AGEMA_signal_27306 ;
    wire new_AGEMA_signal_27307 ;
    wire new_AGEMA_signal_27308 ;
    wire new_AGEMA_signal_27309 ;
    wire new_AGEMA_signal_27310 ;
    wire new_AGEMA_signal_27311 ;
    wire new_AGEMA_signal_27312 ;
    wire new_AGEMA_signal_27313 ;
    wire new_AGEMA_signal_27314 ;
    wire new_AGEMA_signal_27315 ;
    wire new_AGEMA_signal_27316 ;
    wire new_AGEMA_signal_27317 ;
    wire new_AGEMA_signal_27318 ;
    wire new_AGEMA_signal_27319 ;
    wire new_AGEMA_signal_27320 ;
    wire new_AGEMA_signal_27321 ;
    wire new_AGEMA_signal_27322 ;
    wire new_AGEMA_signal_27323 ;
    wire new_AGEMA_signal_27324 ;
    wire new_AGEMA_signal_27325 ;
    wire new_AGEMA_signal_27326 ;
    wire new_AGEMA_signal_27327 ;
    wire new_AGEMA_signal_27328 ;
    wire new_AGEMA_signal_27329 ;
    wire new_AGEMA_signal_27330 ;
    wire new_AGEMA_signal_27331 ;
    wire new_AGEMA_signal_27332 ;
    wire new_AGEMA_signal_27333 ;
    wire new_AGEMA_signal_27334 ;
    wire new_AGEMA_signal_27335 ;
    wire new_AGEMA_signal_27336 ;
    wire new_AGEMA_signal_27337 ;
    wire new_AGEMA_signal_27338 ;
    wire new_AGEMA_signal_27339 ;
    wire new_AGEMA_signal_27340 ;
    wire new_AGEMA_signal_27341 ;
    wire new_AGEMA_signal_27342 ;
    wire new_AGEMA_signal_27343 ;
    wire new_AGEMA_signal_27344 ;
    wire new_AGEMA_signal_27345 ;
    wire new_AGEMA_signal_27346 ;
    wire new_AGEMA_signal_27347 ;
    wire new_AGEMA_signal_27348 ;
    wire new_AGEMA_signal_27349 ;
    wire new_AGEMA_signal_27350 ;
    wire new_AGEMA_signal_27351 ;
    wire new_AGEMA_signal_27352 ;
    wire new_AGEMA_signal_27353 ;
    wire new_AGEMA_signal_27354 ;
    wire new_AGEMA_signal_27355 ;
    wire new_AGEMA_signal_27356 ;
    wire new_AGEMA_signal_27357 ;
    wire new_AGEMA_signal_27358 ;
    wire new_AGEMA_signal_27359 ;
    wire new_AGEMA_signal_27360 ;
    wire new_AGEMA_signal_27361 ;
    wire new_AGEMA_signal_27362 ;
    wire new_AGEMA_signal_27363 ;
    wire new_AGEMA_signal_27364 ;
    wire new_AGEMA_signal_27365 ;
    wire new_AGEMA_signal_27366 ;
    wire new_AGEMA_signal_27367 ;
    wire new_AGEMA_signal_27368 ;
    wire new_AGEMA_signal_27369 ;
    wire new_AGEMA_signal_27370 ;
    wire new_AGEMA_signal_27371 ;
    wire new_AGEMA_signal_27372 ;
    wire new_AGEMA_signal_27373 ;
    wire new_AGEMA_signal_27374 ;
    wire new_AGEMA_signal_27375 ;
    wire new_AGEMA_signal_27376 ;
    wire new_AGEMA_signal_27377 ;
    wire new_AGEMA_signal_27378 ;
    wire new_AGEMA_signal_27379 ;
    wire new_AGEMA_signal_27380 ;
    wire new_AGEMA_signal_27381 ;
    wire new_AGEMA_signal_27382 ;
    wire new_AGEMA_signal_27383 ;
    wire new_AGEMA_signal_27384 ;
    wire new_AGEMA_signal_27385 ;
    wire new_AGEMA_signal_27386 ;
    wire new_AGEMA_signal_27387 ;
    wire new_AGEMA_signal_27388 ;
    wire new_AGEMA_signal_27389 ;
    wire new_AGEMA_signal_27390 ;
    wire new_AGEMA_signal_27391 ;
    wire new_AGEMA_signal_27392 ;
    wire new_AGEMA_signal_27393 ;
    wire new_AGEMA_signal_27394 ;
    wire new_AGEMA_signal_27395 ;
    wire new_AGEMA_signal_27396 ;
    wire new_AGEMA_signal_27397 ;
    wire new_AGEMA_signal_27398 ;
    wire new_AGEMA_signal_27399 ;
    wire new_AGEMA_signal_27400 ;
    wire new_AGEMA_signal_27401 ;
    wire new_AGEMA_signal_27402 ;
    wire new_AGEMA_signal_27403 ;
    wire new_AGEMA_signal_27404 ;
    wire new_AGEMA_signal_27405 ;
    wire new_AGEMA_signal_27406 ;
    wire new_AGEMA_signal_27407 ;
    wire new_AGEMA_signal_27408 ;
    wire new_AGEMA_signal_27409 ;
    wire new_AGEMA_signal_27410 ;
    wire new_AGEMA_signal_27411 ;
    wire new_AGEMA_signal_27412 ;
    wire new_AGEMA_signal_27413 ;
    wire new_AGEMA_signal_27414 ;
    wire new_AGEMA_signal_27415 ;
    wire new_AGEMA_signal_27416 ;
    wire new_AGEMA_signal_27417 ;
    wire new_AGEMA_signal_27418 ;
    wire new_AGEMA_signal_27419 ;
    wire new_AGEMA_signal_27420 ;
    wire new_AGEMA_signal_27421 ;
    wire new_AGEMA_signal_27422 ;
    wire new_AGEMA_signal_27423 ;
    wire new_AGEMA_signal_27424 ;
    wire new_AGEMA_signal_27425 ;
    wire new_AGEMA_signal_27426 ;
    wire new_AGEMA_signal_27427 ;
    wire new_AGEMA_signal_27428 ;
    wire new_AGEMA_signal_27429 ;
    wire new_AGEMA_signal_27430 ;
    wire new_AGEMA_signal_27431 ;
    wire new_AGEMA_signal_27432 ;
    wire new_AGEMA_signal_27433 ;
    wire new_AGEMA_signal_27434 ;
    wire new_AGEMA_signal_27435 ;
    wire new_AGEMA_signal_27436 ;
    wire new_AGEMA_signal_27437 ;
    wire new_AGEMA_signal_27438 ;
    wire new_AGEMA_signal_27439 ;
    wire new_AGEMA_signal_27440 ;
    wire new_AGEMA_signal_27441 ;
    wire new_AGEMA_signal_27442 ;
    wire new_AGEMA_signal_27443 ;
    wire new_AGEMA_signal_27444 ;
    wire new_AGEMA_signal_27445 ;
    wire new_AGEMA_signal_27446 ;
    wire new_AGEMA_signal_27447 ;
    wire new_AGEMA_signal_27448 ;
    wire new_AGEMA_signal_27449 ;
    wire new_AGEMA_signal_27450 ;
    wire new_AGEMA_signal_27451 ;
    wire new_AGEMA_signal_27452 ;
    wire new_AGEMA_signal_27453 ;
    wire new_AGEMA_signal_27454 ;
    wire new_AGEMA_signal_27455 ;
    wire new_AGEMA_signal_27456 ;
    wire new_AGEMA_signal_27457 ;
    wire new_AGEMA_signal_27458 ;
    wire new_AGEMA_signal_27459 ;
    wire new_AGEMA_signal_27460 ;
    wire new_AGEMA_signal_27461 ;
    wire new_AGEMA_signal_27462 ;
    wire new_AGEMA_signal_27463 ;
    wire new_AGEMA_signal_27464 ;
    wire new_AGEMA_signal_27465 ;
    wire new_AGEMA_signal_27466 ;
    wire new_AGEMA_signal_27467 ;
    wire new_AGEMA_signal_27468 ;
    wire new_AGEMA_signal_27469 ;
    wire new_AGEMA_signal_27470 ;
    wire new_AGEMA_signal_27471 ;
    wire new_AGEMA_signal_27472 ;
    wire new_AGEMA_signal_27473 ;
    wire new_AGEMA_signal_27474 ;
    wire new_AGEMA_signal_27475 ;
    wire new_AGEMA_signal_27476 ;
    wire new_AGEMA_signal_27477 ;
    wire new_AGEMA_signal_27478 ;
    wire new_AGEMA_signal_27479 ;
    wire new_AGEMA_signal_27480 ;
    wire new_AGEMA_signal_27481 ;
    wire new_AGEMA_signal_27482 ;
    wire new_AGEMA_signal_27483 ;
    wire new_AGEMA_signal_27484 ;
    wire new_AGEMA_signal_27485 ;
    wire new_AGEMA_signal_27486 ;
    wire new_AGEMA_signal_27487 ;
    wire new_AGEMA_signal_27488 ;
    wire new_AGEMA_signal_27489 ;
    wire new_AGEMA_signal_27490 ;
    wire new_AGEMA_signal_27491 ;
    wire new_AGEMA_signal_27492 ;
    wire new_AGEMA_signal_27493 ;
    wire new_AGEMA_signal_27494 ;
    wire new_AGEMA_signal_27495 ;
    wire new_AGEMA_signal_27496 ;
    wire new_AGEMA_signal_27497 ;
    wire new_AGEMA_signal_27498 ;
    wire new_AGEMA_signal_27499 ;
    wire new_AGEMA_signal_27500 ;
    wire new_AGEMA_signal_27501 ;
    wire new_AGEMA_signal_27502 ;
    wire new_AGEMA_signal_27503 ;
    wire new_AGEMA_signal_27504 ;
    wire new_AGEMA_signal_27505 ;
    wire new_AGEMA_signal_27506 ;
    wire new_AGEMA_signal_27507 ;
    wire new_AGEMA_signal_27508 ;
    wire new_AGEMA_signal_27509 ;
    wire new_AGEMA_signal_27510 ;
    wire new_AGEMA_signal_27511 ;
    wire new_AGEMA_signal_27512 ;
    wire new_AGEMA_signal_27513 ;
    wire new_AGEMA_signal_27514 ;
    wire new_AGEMA_signal_27515 ;
    wire new_AGEMA_signal_27516 ;
    wire new_AGEMA_signal_27517 ;
    wire new_AGEMA_signal_27518 ;
    wire new_AGEMA_signal_27519 ;
    wire new_AGEMA_signal_27520 ;
    wire new_AGEMA_signal_27521 ;
    wire new_AGEMA_signal_27522 ;
    wire new_AGEMA_signal_27523 ;
    wire new_AGEMA_signal_27524 ;
    wire new_AGEMA_signal_27525 ;
    wire new_AGEMA_signal_27526 ;
    wire new_AGEMA_signal_27527 ;
    wire new_AGEMA_signal_27528 ;
    wire new_AGEMA_signal_27529 ;
    wire new_AGEMA_signal_27530 ;
    wire new_AGEMA_signal_27531 ;
    wire new_AGEMA_signal_27532 ;
    wire new_AGEMA_signal_27533 ;
    wire new_AGEMA_signal_27534 ;
    wire new_AGEMA_signal_27535 ;
    wire new_AGEMA_signal_27536 ;
    wire new_AGEMA_signal_27537 ;
    wire new_AGEMA_signal_27538 ;
    wire new_AGEMA_signal_27539 ;
    wire new_AGEMA_signal_27540 ;
    wire new_AGEMA_signal_27541 ;
    wire new_AGEMA_signal_27542 ;
    wire new_AGEMA_signal_27543 ;
    wire new_AGEMA_signal_27544 ;
    wire new_AGEMA_signal_27545 ;
    wire new_AGEMA_signal_27546 ;
    wire new_AGEMA_signal_27547 ;
    wire new_AGEMA_signal_27548 ;
    wire new_AGEMA_signal_27549 ;
    wire new_AGEMA_signal_27550 ;
    wire new_AGEMA_signal_27551 ;
    wire new_AGEMA_signal_27552 ;
    wire new_AGEMA_signal_27553 ;
    wire new_AGEMA_signal_27554 ;
    wire new_AGEMA_signal_27555 ;
    wire new_AGEMA_signal_27556 ;
    wire new_AGEMA_signal_27557 ;
    wire new_AGEMA_signal_27558 ;
    wire new_AGEMA_signal_27559 ;
    wire new_AGEMA_signal_27560 ;
    wire new_AGEMA_signal_27561 ;
    wire new_AGEMA_signal_27562 ;
    wire new_AGEMA_signal_27563 ;
    wire new_AGEMA_signal_27564 ;
    wire new_AGEMA_signal_27565 ;
    wire new_AGEMA_signal_27566 ;
    wire new_AGEMA_signal_27567 ;
    wire new_AGEMA_signal_27568 ;
    wire new_AGEMA_signal_27569 ;
    wire new_AGEMA_signal_27570 ;
    wire new_AGEMA_signal_27571 ;
    wire new_AGEMA_signal_27572 ;
    wire new_AGEMA_signal_27573 ;
    wire new_AGEMA_signal_27574 ;
    wire new_AGEMA_signal_27575 ;
    wire new_AGEMA_signal_27576 ;
    wire new_AGEMA_signal_27577 ;
    wire new_AGEMA_signal_27578 ;
    wire new_AGEMA_signal_27579 ;
    wire new_AGEMA_signal_27580 ;
    wire new_AGEMA_signal_27581 ;
    wire new_AGEMA_signal_27582 ;
    wire new_AGEMA_signal_27583 ;
    wire new_AGEMA_signal_27584 ;
    wire new_AGEMA_signal_27585 ;
    wire new_AGEMA_signal_27586 ;
    wire new_AGEMA_signal_27587 ;
    wire new_AGEMA_signal_27588 ;
    wire new_AGEMA_signal_27589 ;
    wire new_AGEMA_signal_27590 ;
    wire new_AGEMA_signal_27591 ;
    wire new_AGEMA_signal_27592 ;
    wire new_AGEMA_signal_27593 ;
    wire new_AGEMA_signal_27594 ;
    wire new_AGEMA_signal_27595 ;
    wire new_AGEMA_signal_27596 ;
    wire new_AGEMA_signal_27597 ;
    wire new_AGEMA_signal_27598 ;
    wire new_AGEMA_signal_27599 ;
    wire new_AGEMA_signal_27600 ;
    wire new_AGEMA_signal_27601 ;
    wire new_AGEMA_signal_27602 ;
    wire new_AGEMA_signal_27603 ;
    wire new_AGEMA_signal_27604 ;
    wire new_AGEMA_signal_27605 ;
    wire new_AGEMA_signal_27606 ;
    wire new_AGEMA_signal_27607 ;
    wire new_AGEMA_signal_27608 ;
    wire new_AGEMA_signal_27609 ;
    wire new_AGEMA_signal_27610 ;
    wire new_AGEMA_signal_27611 ;
    wire new_AGEMA_signal_27612 ;
    wire new_AGEMA_signal_27613 ;
    wire new_AGEMA_signal_27614 ;
    wire new_AGEMA_signal_27615 ;
    wire new_AGEMA_signal_27616 ;
    wire new_AGEMA_signal_27617 ;
    wire new_AGEMA_signal_27618 ;
    wire new_AGEMA_signal_27619 ;
    wire new_AGEMA_signal_27620 ;
    wire new_AGEMA_signal_27621 ;
    wire new_AGEMA_signal_27622 ;
    wire new_AGEMA_signal_27623 ;
    wire new_AGEMA_signal_27624 ;
    wire new_AGEMA_signal_27625 ;
    wire new_AGEMA_signal_27626 ;
    wire new_AGEMA_signal_27627 ;
    wire new_AGEMA_signal_27628 ;
    wire new_AGEMA_signal_27629 ;
    wire new_AGEMA_signal_27630 ;
    wire new_AGEMA_signal_27631 ;
    wire new_AGEMA_signal_27632 ;
    wire new_AGEMA_signal_27633 ;
    wire new_AGEMA_signal_27634 ;
    wire new_AGEMA_signal_27635 ;
    wire new_AGEMA_signal_27636 ;
    wire new_AGEMA_signal_27637 ;
    wire new_AGEMA_signal_27638 ;
    wire new_AGEMA_signal_27639 ;
    wire new_AGEMA_signal_27640 ;
    wire new_AGEMA_signal_27641 ;
    wire new_AGEMA_signal_27642 ;
    wire new_AGEMA_signal_27643 ;
    wire new_AGEMA_signal_27644 ;
    wire new_AGEMA_signal_27645 ;
    wire new_AGEMA_signal_27646 ;
    wire new_AGEMA_signal_27647 ;
    wire new_AGEMA_signal_27648 ;
    wire new_AGEMA_signal_27649 ;
    wire new_AGEMA_signal_27650 ;
    wire new_AGEMA_signal_27651 ;
    wire new_AGEMA_signal_27652 ;
    wire new_AGEMA_signal_27653 ;
    wire new_AGEMA_signal_27654 ;
    wire new_AGEMA_signal_27655 ;
    wire new_AGEMA_signal_27656 ;
    wire new_AGEMA_signal_27657 ;
    wire new_AGEMA_signal_27658 ;
    wire new_AGEMA_signal_27659 ;
    wire new_AGEMA_signal_27660 ;
    wire new_AGEMA_signal_27661 ;
    wire new_AGEMA_signal_27662 ;
    wire new_AGEMA_signal_27663 ;
    wire new_AGEMA_signal_27664 ;
    wire new_AGEMA_signal_27665 ;
    wire new_AGEMA_signal_27666 ;
    wire new_AGEMA_signal_27667 ;
    wire new_AGEMA_signal_27668 ;
    wire new_AGEMA_signal_27669 ;
    wire new_AGEMA_signal_27670 ;
    wire new_AGEMA_signal_27671 ;
    wire new_AGEMA_signal_27672 ;
    wire new_AGEMA_signal_27673 ;
    wire new_AGEMA_signal_27674 ;
    wire new_AGEMA_signal_27675 ;
    wire new_AGEMA_signal_27676 ;
    wire new_AGEMA_signal_27677 ;
    wire new_AGEMA_signal_27678 ;
    wire new_AGEMA_signal_27679 ;
    wire new_AGEMA_signal_27680 ;
    wire new_AGEMA_signal_27681 ;
    wire new_AGEMA_signal_27682 ;
    wire new_AGEMA_signal_27683 ;
    wire new_AGEMA_signal_27684 ;
    wire new_AGEMA_signal_27685 ;
    wire new_AGEMA_signal_27686 ;
    wire new_AGEMA_signal_27687 ;
    wire new_AGEMA_signal_27688 ;
    wire new_AGEMA_signal_27689 ;
    wire new_AGEMA_signal_27690 ;
    wire new_AGEMA_signal_27691 ;
    wire new_AGEMA_signal_27692 ;
    wire new_AGEMA_signal_27693 ;
    wire new_AGEMA_signal_27694 ;
    wire new_AGEMA_signal_27695 ;
    wire new_AGEMA_signal_27696 ;
    wire new_AGEMA_signal_27697 ;
    wire new_AGEMA_signal_27698 ;
    wire new_AGEMA_signal_27699 ;
    wire new_AGEMA_signal_27700 ;
    wire new_AGEMA_signal_27701 ;
    wire new_AGEMA_signal_27702 ;
    wire new_AGEMA_signal_27703 ;
    wire new_AGEMA_signal_27704 ;
    wire new_AGEMA_signal_27705 ;
    wire new_AGEMA_signal_27706 ;
    wire new_AGEMA_signal_27707 ;
    wire new_AGEMA_signal_27708 ;
    wire new_AGEMA_signal_27709 ;
    wire new_AGEMA_signal_27710 ;
    wire new_AGEMA_signal_27711 ;
    wire new_AGEMA_signal_27712 ;
    wire new_AGEMA_signal_27713 ;
    wire new_AGEMA_signal_27714 ;
    wire new_AGEMA_signal_27715 ;
    wire new_AGEMA_signal_27716 ;
    wire new_AGEMA_signal_27717 ;
    wire new_AGEMA_signal_27718 ;
    wire new_AGEMA_signal_27719 ;
    wire new_AGEMA_signal_27720 ;
    wire new_AGEMA_signal_27721 ;
    wire new_AGEMA_signal_27722 ;
    wire new_AGEMA_signal_27723 ;
    wire new_AGEMA_signal_27724 ;
    wire new_AGEMA_signal_27725 ;
    wire new_AGEMA_signal_27726 ;
    wire new_AGEMA_signal_27727 ;
    wire new_AGEMA_signal_27728 ;
    wire new_AGEMA_signal_27729 ;
    wire new_AGEMA_signal_27730 ;
    wire new_AGEMA_signal_27731 ;
    wire new_AGEMA_signal_27732 ;
    wire new_AGEMA_signal_27733 ;
    wire new_AGEMA_signal_27734 ;
    wire new_AGEMA_signal_27735 ;
    wire new_AGEMA_signal_27736 ;
    wire new_AGEMA_signal_27737 ;
    wire new_AGEMA_signal_27738 ;
    wire new_AGEMA_signal_27739 ;
    wire new_AGEMA_signal_27740 ;
    wire new_AGEMA_signal_27741 ;
    wire new_AGEMA_signal_27742 ;
    wire new_AGEMA_signal_27743 ;
    wire new_AGEMA_signal_27744 ;
    wire new_AGEMA_signal_27745 ;
    wire new_AGEMA_signal_27746 ;
    wire new_AGEMA_signal_27747 ;
    wire new_AGEMA_signal_27748 ;
    wire new_AGEMA_signal_27749 ;
    wire new_AGEMA_signal_27750 ;
    wire new_AGEMA_signal_27751 ;
    wire new_AGEMA_signal_27752 ;
    wire new_AGEMA_signal_27753 ;
    wire new_AGEMA_signal_27754 ;
    wire new_AGEMA_signal_27755 ;
    wire new_AGEMA_signal_27756 ;
    wire new_AGEMA_signal_27757 ;
    wire new_AGEMA_signal_27758 ;
    wire new_AGEMA_signal_27759 ;
    wire new_AGEMA_signal_27760 ;
    wire new_AGEMA_signal_27761 ;
    wire new_AGEMA_signal_27762 ;
    wire new_AGEMA_signal_27763 ;
    wire new_AGEMA_signal_27764 ;
    wire new_AGEMA_signal_27765 ;
    wire new_AGEMA_signal_27766 ;
    wire new_AGEMA_signal_27767 ;
    wire new_AGEMA_signal_27768 ;
    wire new_AGEMA_signal_27769 ;
    wire new_AGEMA_signal_27770 ;
    wire new_AGEMA_signal_27771 ;
    wire new_AGEMA_signal_27772 ;
    wire new_AGEMA_signal_27773 ;
    wire new_AGEMA_signal_27774 ;
    wire new_AGEMA_signal_27775 ;
    wire new_AGEMA_signal_27776 ;
    wire new_AGEMA_signal_27777 ;
    wire new_AGEMA_signal_27778 ;
    wire new_AGEMA_signal_27779 ;
    wire new_AGEMA_signal_27780 ;
    wire new_AGEMA_signal_27781 ;
    wire new_AGEMA_signal_27782 ;
    wire new_AGEMA_signal_27783 ;
    wire new_AGEMA_signal_27784 ;
    wire new_AGEMA_signal_27785 ;
    wire new_AGEMA_signal_27786 ;
    wire new_AGEMA_signal_27787 ;
    wire new_AGEMA_signal_27788 ;
    wire new_AGEMA_signal_27789 ;
    wire new_AGEMA_signal_27790 ;
    wire new_AGEMA_signal_27791 ;
    wire new_AGEMA_signal_27792 ;
    wire new_AGEMA_signal_27793 ;
    wire new_AGEMA_signal_27794 ;
    wire new_AGEMA_signal_27795 ;
    wire new_AGEMA_signal_27796 ;
    wire new_AGEMA_signal_27797 ;
    wire new_AGEMA_signal_27798 ;
    wire new_AGEMA_signal_27799 ;
    wire new_AGEMA_signal_27800 ;
    wire new_AGEMA_signal_27801 ;
    wire new_AGEMA_signal_27802 ;
    wire new_AGEMA_signal_27803 ;
    wire new_AGEMA_signal_27804 ;
    wire new_AGEMA_signal_27805 ;
    wire new_AGEMA_signal_27806 ;
    wire new_AGEMA_signal_27807 ;
    wire new_AGEMA_signal_27808 ;
    wire new_AGEMA_signal_27809 ;
    wire new_AGEMA_signal_27810 ;
    wire new_AGEMA_signal_27811 ;
    wire new_AGEMA_signal_27812 ;
    wire new_AGEMA_signal_27813 ;
    wire new_AGEMA_signal_27814 ;
    wire new_AGEMA_signal_27815 ;
    wire new_AGEMA_signal_27816 ;
    wire new_AGEMA_signal_27817 ;
    wire new_AGEMA_signal_27818 ;
    wire new_AGEMA_signal_27819 ;
    wire new_AGEMA_signal_27820 ;
    wire new_AGEMA_signal_27821 ;
    wire new_AGEMA_signal_27822 ;
    wire new_AGEMA_signal_27823 ;
    wire new_AGEMA_signal_27824 ;
    wire new_AGEMA_signal_27825 ;
    wire new_AGEMA_signal_27826 ;
    wire new_AGEMA_signal_27827 ;
    wire new_AGEMA_signal_27828 ;
    wire new_AGEMA_signal_27829 ;
    wire new_AGEMA_signal_27830 ;
    wire new_AGEMA_signal_27831 ;
    wire new_AGEMA_signal_27832 ;
    wire new_AGEMA_signal_27833 ;
    wire new_AGEMA_signal_27834 ;
    wire new_AGEMA_signal_27835 ;
    wire new_AGEMA_signal_27836 ;
    wire new_AGEMA_signal_27837 ;
    wire new_AGEMA_signal_27838 ;
    wire new_AGEMA_signal_27839 ;
    wire new_AGEMA_signal_27840 ;
    wire new_AGEMA_signal_27841 ;
    wire new_AGEMA_signal_27842 ;
    wire new_AGEMA_signal_27843 ;
    wire new_AGEMA_signal_27844 ;
    wire new_AGEMA_signal_27845 ;
    wire new_AGEMA_signal_27846 ;
    wire new_AGEMA_signal_27847 ;
    wire new_AGEMA_signal_27848 ;
    wire new_AGEMA_signal_27849 ;
    wire new_AGEMA_signal_27850 ;
    wire new_AGEMA_signal_27851 ;
    wire new_AGEMA_signal_27852 ;
    wire new_AGEMA_signal_27853 ;
    wire new_AGEMA_signal_27854 ;
    wire new_AGEMA_signal_27855 ;
    wire new_AGEMA_signal_27856 ;
    wire new_AGEMA_signal_27857 ;
    wire new_AGEMA_signal_27858 ;
    wire new_AGEMA_signal_27859 ;
    wire new_AGEMA_signal_27860 ;
    wire new_AGEMA_signal_27861 ;
    wire new_AGEMA_signal_27862 ;
    wire new_AGEMA_signal_27863 ;
    wire new_AGEMA_signal_27864 ;
    wire new_AGEMA_signal_27865 ;
    wire new_AGEMA_signal_27866 ;
    wire new_AGEMA_signal_27867 ;
    wire new_AGEMA_signal_27868 ;
    wire new_AGEMA_signal_27869 ;
    wire new_AGEMA_signal_27870 ;
    wire new_AGEMA_signal_27871 ;
    wire new_AGEMA_signal_27872 ;
    wire new_AGEMA_signal_27873 ;
    wire new_AGEMA_signal_27874 ;
    wire new_AGEMA_signal_27875 ;
    wire new_AGEMA_signal_27876 ;
    wire new_AGEMA_signal_27877 ;
    wire new_AGEMA_signal_27878 ;
    wire new_AGEMA_signal_27879 ;
    wire new_AGEMA_signal_27880 ;
    wire new_AGEMA_signal_27881 ;
    wire new_AGEMA_signal_27882 ;
    wire new_AGEMA_signal_27883 ;
    wire new_AGEMA_signal_27884 ;
    wire new_AGEMA_signal_27885 ;
    wire new_AGEMA_signal_27886 ;
    wire new_AGEMA_signal_27887 ;
    wire new_AGEMA_signal_27888 ;
    wire new_AGEMA_signal_27889 ;
    wire new_AGEMA_signal_27890 ;
    wire new_AGEMA_signal_27891 ;
    wire new_AGEMA_signal_27892 ;
    wire new_AGEMA_signal_27893 ;
    wire new_AGEMA_signal_27894 ;
    wire new_AGEMA_signal_27895 ;
    wire new_AGEMA_signal_27896 ;
    wire new_AGEMA_signal_27897 ;
    wire new_AGEMA_signal_27898 ;
    wire new_AGEMA_signal_27899 ;
    wire new_AGEMA_signal_27900 ;
    wire new_AGEMA_signal_27901 ;
    wire new_AGEMA_signal_27902 ;
    wire new_AGEMA_signal_27903 ;
    wire new_AGEMA_signal_27904 ;
    wire new_AGEMA_signal_27905 ;
    wire new_AGEMA_signal_27906 ;
    wire new_AGEMA_signal_27907 ;
    wire new_AGEMA_signal_27908 ;
    wire new_AGEMA_signal_27909 ;
    wire new_AGEMA_signal_27910 ;
    wire new_AGEMA_signal_27911 ;
    wire new_AGEMA_signal_27912 ;
    wire new_AGEMA_signal_27913 ;
    wire new_AGEMA_signal_27914 ;
    wire new_AGEMA_signal_27915 ;
    wire new_AGEMA_signal_27916 ;
    wire new_AGEMA_signal_27917 ;
    wire new_AGEMA_signal_27918 ;
    wire new_AGEMA_signal_27919 ;
    wire new_AGEMA_signal_27920 ;
    wire new_AGEMA_signal_27921 ;
    wire new_AGEMA_signal_27922 ;
    wire new_AGEMA_signal_27923 ;
    wire new_AGEMA_signal_27924 ;
    wire new_AGEMA_signal_27925 ;
    wire new_AGEMA_signal_27926 ;
    wire new_AGEMA_signal_27927 ;
    wire new_AGEMA_signal_27928 ;
    wire new_AGEMA_signal_27929 ;
    wire new_AGEMA_signal_27930 ;
    wire new_AGEMA_signal_27931 ;
    wire new_AGEMA_signal_27932 ;
    wire new_AGEMA_signal_27933 ;
    wire new_AGEMA_signal_27934 ;
    wire new_AGEMA_signal_27935 ;
    wire new_AGEMA_signal_27936 ;
    wire new_AGEMA_signal_27937 ;
    wire new_AGEMA_signal_27938 ;
    wire new_AGEMA_signal_27939 ;
    wire new_AGEMA_signal_27940 ;
    wire new_AGEMA_signal_27941 ;
    wire new_AGEMA_signal_27942 ;
    wire new_AGEMA_signal_27943 ;
    wire new_AGEMA_signal_27944 ;
    wire new_AGEMA_signal_27945 ;
    wire new_AGEMA_signal_27946 ;
    wire new_AGEMA_signal_27947 ;
    wire new_AGEMA_signal_27948 ;
    wire new_AGEMA_signal_27949 ;
    wire new_AGEMA_signal_27950 ;
    wire new_AGEMA_signal_27951 ;
    wire new_AGEMA_signal_27952 ;
    wire new_AGEMA_signal_27953 ;
    wire new_AGEMA_signal_27954 ;
    wire new_AGEMA_signal_27955 ;
    wire new_AGEMA_signal_27956 ;
    wire new_AGEMA_signal_27957 ;
    wire new_AGEMA_signal_27958 ;
    wire new_AGEMA_signal_27959 ;
    wire new_AGEMA_signal_27960 ;
    wire new_AGEMA_signal_27961 ;
    wire new_AGEMA_signal_27962 ;
    wire new_AGEMA_signal_27963 ;
    wire new_AGEMA_signal_27964 ;
    wire new_AGEMA_signal_27965 ;
    wire new_AGEMA_signal_27966 ;
    wire new_AGEMA_signal_27967 ;
    wire new_AGEMA_signal_27968 ;
    wire new_AGEMA_signal_27969 ;
    wire new_AGEMA_signal_27970 ;
    wire new_AGEMA_signal_27971 ;
    wire new_AGEMA_signal_27972 ;
    wire new_AGEMA_signal_27973 ;
    wire new_AGEMA_signal_27974 ;
    wire new_AGEMA_signal_27975 ;
    wire new_AGEMA_signal_27976 ;
    wire new_AGEMA_signal_27977 ;
    wire new_AGEMA_signal_27978 ;
    wire new_AGEMA_signal_27979 ;
    wire new_AGEMA_signal_27980 ;
    wire new_AGEMA_signal_27981 ;
    wire new_AGEMA_signal_27982 ;
    wire new_AGEMA_signal_27983 ;
    wire new_AGEMA_signal_27984 ;
    wire new_AGEMA_signal_27985 ;
    wire new_AGEMA_signal_27986 ;
    wire new_AGEMA_signal_27987 ;
    wire new_AGEMA_signal_27988 ;
    wire new_AGEMA_signal_27989 ;
    wire new_AGEMA_signal_27990 ;
    wire new_AGEMA_signal_27991 ;
    wire new_AGEMA_signal_27992 ;
    wire new_AGEMA_signal_27993 ;
    wire new_AGEMA_signal_27994 ;
    wire new_AGEMA_signal_27995 ;
    wire new_AGEMA_signal_27996 ;
    wire new_AGEMA_signal_27997 ;
    wire new_AGEMA_signal_27998 ;
    wire new_AGEMA_signal_27999 ;
    wire new_AGEMA_signal_28000 ;
    wire new_AGEMA_signal_28001 ;
    wire new_AGEMA_signal_28002 ;
    wire new_AGEMA_signal_28003 ;
    wire new_AGEMA_signal_28004 ;
    wire new_AGEMA_signal_28005 ;
    wire new_AGEMA_signal_28006 ;
    wire new_AGEMA_signal_28007 ;
    wire new_AGEMA_signal_28008 ;
    wire new_AGEMA_signal_28009 ;
    wire new_AGEMA_signal_28010 ;
    wire new_AGEMA_signal_28011 ;
    wire new_AGEMA_signal_28012 ;
    wire new_AGEMA_signal_28013 ;
    wire new_AGEMA_signal_28014 ;
    wire new_AGEMA_signal_28015 ;
    wire new_AGEMA_signal_28016 ;
    wire new_AGEMA_signal_28017 ;
    wire new_AGEMA_signal_28018 ;
    wire new_AGEMA_signal_28019 ;
    wire new_AGEMA_signal_28020 ;
    wire new_AGEMA_signal_28021 ;
    wire new_AGEMA_signal_28022 ;
    wire new_AGEMA_signal_28023 ;
    wire new_AGEMA_signal_28024 ;
    wire new_AGEMA_signal_28025 ;
    wire new_AGEMA_signal_28026 ;
    wire new_AGEMA_signal_28027 ;
    wire new_AGEMA_signal_28028 ;
    wire new_AGEMA_signal_28029 ;
    wire new_AGEMA_signal_28030 ;
    wire new_AGEMA_signal_28031 ;
    wire new_AGEMA_signal_28032 ;
    wire new_AGEMA_signal_28033 ;
    wire new_AGEMA_signal_28034 ;
    wire new_AGEMA_signal_28035 ;
    wire new_AGEMA_signal_28036 ;
    wire new_AGEMA_signal_28037 ;
    wire new_AGEMA_signal_28038 ;
    wire new_AGEMA_signal_28039 ;
    wire new_AGEMA_signal_28040 ;
    wire new_AGEMA_signal_28041 ;
    wire new_AGEMA_signal_28042 ;
    wire new_AGEMA_signal_28043 ;
    wire new_AGEMA_signal_28044 ;
    wire new_AGEMA_signal_28045 ;
    wire new_AGEMA_signal_28046 ;
    wire new_AGEMA_signal_28047 ;
    wire new_AGEMA_signal_28048 ;
    wire new_AGEMA_signal_28049 ;
    wire new_AGEMA_signal_28050 ;
    wire new_AGEMA_signal_28051 ;
    wire new_AGEMA_signal_28052 ;
    wire new_AGEMA_signal_28053 ;
    wire new_AGEMA_signal_28054 ;
    wire new_AGEMA_signal_28055 ;
    wire new_AGEMA_signal_28056 ;
    wire new_AGEMA_signal_28057 ;
    wire new_AGEMA_signal_28058 ;
    wire new_AGEMA_signal_28059 ;
    wire new_AGEMA_signal_28060 ;
    wire new_AGEMA_signal_28061 ;
    wire new_AGEMA_signal_28062 ;
    wire new_AGEMA_signal_28063 ;
    wire new_AGEMA_signal_28064 ;
    wire new_AGEMA_signal_28065 ;
    wire new_AGEMA_signal_28066 ;
    wire new_AGEMA_signal_28067 ;
    wire new_AGEMA_signal_28068 ;
    wire new_AGEMA_signal_28069 ;
    wire new_AGEMA_signal_28070 ;
    wire new_AGEMA_signal_28071 ;
    wire new_AGEMA_signal_28072 ;
    wire new_AGEMA_signal_28073 ;
    wire new_AGEMA_signal_28074 ;
    wire new_AGEMA_signal_28075 ;
    wire new_AGEMA_signal_28076 ;
    wire new_AGEMA_signal_28077 ;
    wire new_AGEMA_signal_28078 ;
    wire new_AGEMA_signal_28079 ;
    wire new_AGEMA_signal_28080 ;
    wire new_AGEMA_signal_28081 ;
    wire new_AGEMA_signal_28082 ;
    wire new_AGEMA_signal_28083 ;
    wire new_AGEMA_signal_28084 ;
    wire new_AGEMA_signal_28085 ;
    wire new_AGEMA_signal_28086 ;
    wire new_AGEMA_signal_28087 ;
    wire new_AGEMA_signal_28088 ;
    wire new_AGEMA_signal_28089 ;
    wire new_AGEMA_signal_28090 ;
    wire new_AGEMA_signal_28091 ;
    wire new_AGEMA_signal_28092 ;
    wire new_AGEMA_signal_28093 ;
    wire new_AGEMA_signal_28094 ;
    wire new_AGEMA_signal_28095 ;
    wire new_AGEMA_signal_28096 ;
    wire new_AGEMA_signal_28097 ;
    wire new_AGEMA_signal_28098 ;
    wire new_AGEMA_signal_28099 ;
    wire new_AGEMA_signal_28100 ;
    wire new_AGEMA_signal_28101 ;
    wire new_AGEMA_signal_28102 ;
    wire new_AGEMA_signal_28103 ;
    wire new_AGEMA_signal_28104 ;
    wire new_AGEMA_signal_28105 ;
    wire new_AGEMA_signal_28106 ;
    wire new_AGEMA_signal_28107 ;
    wire new_AGEMA_signal_28108 ;
    wire new_AGEMA_signal_28109 ;
    wire new_AGEMA_signal_28110 ;
    wire new_AGEMA_signal_28111 ;
    wire new_AGEMA_signal_28112 ;
    wire new_AGEMA_signal_28113 ;
    wire new_AGEMA_signal_28114 ;
    wire new_AGEMA_signal_28115 ;
    wire new_AGEMA_signal_28116 ;
    wire new_AGEMA_signal_28117 ;
    wire new_AGEMA_signal_28118 ;
    wire new_AGEMA_signal_28119 ;
    wire new_AGEMA_signal_28120 ;
    wire new_AGEMA_signal_28121 ;
    wire new_AGEMA_signal_28122 ;
    wire new_AGEMA_signal_28123 ;
    wire new_AGEMA_signal_28124 ;
    wire new_AGEMA_signal_28125 ;
    wire new_AGEMA_signal_28126 ;
    wire new_AGEMA_signal_28127 ;
    wire new_AGEMA_signal_28128 ;
    wire new_AGEMA_signal_28129 ;
    wire new_AGEMA_signal_28130 ;
    wire new_AGEMA_signal_28131 ;
    wire new_AGEMA_signal_28132 ;
    wire new_AGEMA_signal_28133 ;
    wire new_AGEMA_signal_28134 ;
    wire new_AGEMA_signal_28135 ;
    wire new_AGEMA_signal_28136 ;
    wire new_AGEMA_signal_28137 ;
    wire new_AGEMA_signal_28138 ;
    wire new_AGEMA_signal_28139 ;
    wire new_AGEMA_signal_28140 ;
    wire new_AGEMA_signal_28141 ;
    wire new_AGEMA_signal_28142 ;
    wire new_AGEMA_signal_28143 ;
    wire new_AGEMA_signal_28144 ;
    wire new_AGEMA_signal_28145 ;
    wire new_AGEMA_signal_28146 ;
    wire new_AGEMA_signal_28147 ;
    wire new_AGEMA_signal_28148 ;
    wire new_AGEMA_signal_28149 ;
    wire new_AGEMA_signal_28150 ;
    wire new_AGEMA_signal_28151 ;
    wire new_AGEMA_signal_28152 ;
    wire new_AGEMA_signal_28153 ;
    wire new_AGEMA_signal_28154 ;
    wire new_AGEMA_signal_28155 ;
    wire new_AGEMA_signal_28156 ;
    wire new_AGEMA_signal_28157 ;
    wire new_AGEMA_signal_28158 ;
    wire new_AGEMA_signal_28159 ;
    wire new_AGEMA_signal_28160 ;
    wire new_AGEMA_signal_28161 ;
    wire new_AGEMA_signal_28162 ;
    wire new_AGEMA_signal_28163 ;
    wire new_AGEMA_signal_28164 ;
    wire new_AGEMA_signal_28165 ;
    wire new_AGEMA_signal_28166 ;
    wire new_AGEMA_signal_28167 ;
    wire new_AGEMA_signal_28168 ;
    wire new_AGEMA_signal_28169 ;
    wire new_AGEMA_signal_28170 ;
    wire new_AGEMA_signal_28171 ;
    wire new_AGEMA_signal_28172 ;
    wire new_AGEMA_signal_28173 ;
    wire new_AGEMA_signal_28174 ;
    wire new_AGEMA_signal_28175 ;
    wire new_AGEMA_signal_28176 ;
    wire new_AGEMA_signal_28177 ;
    wire new_AGEMA_signal_28178 ;
    wire new_AGEMA_signal_28179 ;
    wire new_AGEMA_signal_28180 ;
    wire new_AGEMA_signal_28181 ;
    wire new_AGEMA_signal_28182 ;
    wire new_AGEMA_signal_28183 ;
    wire new_AGEMA_signal_28184 ;
    wire new_AGEMA_signal_28185 ;
    wire new_AGEMA_signal_28186 ;
    wire new_AGEMA_signal_28187 ;
    wire new_AGEMA_signal_28188 ;
    wire new_AGEMA_signal_28189 ;
    wire new_AGEMA_signal_28190 ;
    wire new_AGEMA_signal_28191 ;
    wire new_AGEMA_signal_28192 ;
    wire new_AGEMA_signal_28193 ;
    wire new_AGEMA_signal_28194 ;
    wire new_AGEMA_signal_28195 ;
    wire new_AGEMA_signal_28196 ;
    wire new_AGEMA_signal_28197 ;
    wire new_AGEMA_signal_28198 ;
    wire new_AGEMA_signal_28199 ;
    wire new_AGEMA_signal_28200 ;
    wire new_AGEMA_signal_28201 ;
    wire new_AGEMA_signal_28202 ;
    wire new_AGEMA_signal_28203 ;
    wire new_AGEMA_signal_28204 ;
    wire new_AGEMA_signal_28205 ;
    wire new_AGEMA_signal_28206 ;
    wire new_AGEMA_signal_28207 ;
    wire new_AGEMA_signal_28208 ;
    wire new_AGEMA_signal_28209 ;
    wire new_AGEMA_signal_28210 ;
    wire new_AGEMA_signal_28211 ;
    wire new_AGEMA_signal_28212 ;
    wire new_AGEMA_signal_28213 ;
    wire new_AGEMA_signal_28214 ;
    wire new_AGEMA_signal_28215 ;
    wire new_AGEMA_signal_28216 ;
    wire new_AGEMA_signal_28217 ;
    wire new_AGEMA_signal_28218 ;
    wire new_AGEMA_signal_28219 ;
    wire new_AGEMA_signal_28220 ;
    wire new_AGEMA_signal_28221 ;
    wire new_AGEMA_signal_28222 ;
    wire new_AGEMA_signal_28223 ;
    wire new_AGEMA_signal_28224 ;
    wire new_AGEMA_signal_28225 ;
    wire new_AGEMA_signal_28226 ;
    wire new_AGEMA_signal_28227 ;
    wire new_AGEMA_signal_28228 ;
    wire new_AGEMA_signal_28229 ;
    wire new_AGEMA_signal_28230 ;
    wire new_AGEMA_signal_28231 ;
    wire new_AGEMA_signal_28232 ;
    wire new_AGEMA_signal_28233 ;
    wire new_AGEMA_signal_28234 ;
    wire new_AGEMA_signal_28235 ;
    wire new_AGEMA_signal_28236 ;
    wire new_AGEMA_signal_28237 ;
    wire new_AGEMA_signal_28238 ;
    wire new_AGEMA_signal_28239 ;
    wire new_AGEMA_signal_28240 ;
    wire new_AGEMA_signal_28241 ;
    wire new_AGEMA_signal_28242 ;
    wire new_AGEMA_signal_28243 ;
    wire new_AGEMA_signal_28244 ;
    wire new_AGEMA_signal_28245 ;
    wire new_AGEMA_signal_28246 ;
    wire new_AGEMA_signal_28247 ;
    wire new_AGEMA_signal_28248 ;
    wire new_AGEMA_signal_28249 ;
    wire new_AGEMA_signal_28250 ;
    wire new_AGEMA_signal_28251 ;
    wire new_AGEMA_signal_28252 ;
    wire new_AGEMA_signal_28253 ;
    wire new_AGEMA_signal_28254 ;
    wire new_AGEMA_signal_28255 ;
    wire new_AGEMA_signal_28256 ;
    wire new_AGEMA_signal_28257 ;
    wire new_AGEMA_signal_28258 ;
    wire new_AGEMA_signal_28259 ;
    wire new_AGEMA_signal_28260 ;
    wire new_AGEMA_signal_28261 ;
    wire new_AGEMA_signal_28262 ;
    wire new_AGEMA_signal_28263 ;
    wire new_AGEMA_signal_28264 ;
    wire new_AGEMA_signal_28265 ;
    wire new_AGEMA_signal_28266 ;
    wire new_AGEMA_signal_28267 ;
    wire new_AGEMA_signal_28268 ;
    wire new_AGEMA_signal_28269 ;
    wire new_AGEMA_signal_28270 ;
    wire new_AGEMA_signal_28271 ;
    wire new_AGEMA_signal_28272 ;
    wire new_AGEMA_signal_28273 ;
    wire new_AGEMA_signal_28274 ;
    wire new_AGEMA_signal_28275 ;
    wire new_AGEMA_signal_28276 ;
    wire new_AGEMA_signal_28277 ;
    wire new_AGEMA_signal_28278 ;
    wire new_AGEMA_signal_28279 ;
    wire new_AGEMA_signal_28280 ;
    wire new_AGEMA_signal_28281 ;
    wire new_AGEMA_signal_28282 ;
    wire new_AGEMA_signal_28283 ;
    wire new_AGEMA_signal_28284 ;
    wire new_AGEMA_signal_28285 ;
    wire new_AGEMA_signal_28286 ;
    wire new_AGEMA_signal_28287 ;
    wire new_AGEMA_signal_28288 ;
    wire new_AGEMA_signal_28289 ;
    wire new_AGEMA_signal_28290 ;
    wire new_AGEMA_signal_28291 ;
    wire new_AGEMA_signal_28292 ;
    wire new_AGEMA_signal_28293 ;
    wire new_AGEMA_signal_28294 ;
    wire new_AGEMA_signal_28295 ;
    wire new_AGEMA_signal_28296 ;
    wire new_AGEMA_signal_28297 ;
    wire new_AGEMA_signal_28298 ;
    wire new_AGEMA_signal_28299 ;
    wire new_AGEMA_signal_28300 ;
    wire new_AGEMA_signal_28301 ;
    wire new_AGEMA_signal_28302 ;
    wire new_AGEMA_signal_28303 ;
    wire new_AGEMA_signal_28304 ;
    wire new_AGEMA_signal_28305 ;
    wire new_AGEMA_signal_28306 ;
    wire new_AGEMA_signal_28307 ;
    wire new_AGEMA_signal_28308 ;
    wire new_AGEMA_signal_28309 ;
    wire new_AGEMA_signal_28310 ;
    wire new_AGEMA_signal_28311 ;
    wire new_AGEMA_signal_28312 ;
    wire new_AGEMA_signal_28313 ;
    wire new_AGEMA_signal_28314 ;
    wire new_AGEMA_signal_28315 ;
    wire new_AGEMA_signal_28316 ;
    wire new_AGEMA_signal_28317 ;
    wire new_AGEMA_signal_28318 ;
    wire new_AGEMA_signal_28319 ;
    wire new_AGEMA_signal_28320 ;
    wire new_AGEMA_signal_28321 ;
    wire new_AGEMA_signal_28322 ;
    wire new_AGEMA_signal_28323 ;
    wire new_AGEMA_signal_28324 ;
    wire new_AGEMA_signal_28325 ;
    wire new_AGEMA_signal_28326 ;
    wire new_AGEMA_signal_28327 ;
    wire new_AGEMA_signal_28328 ;
    wire new_AGEMA_signal_28329 ;
    wire new_AGEMA_signal_28330 ;
    wire new_AGEMA_signal_28331 ;
    wire new_AGEMA_signal_28332 ;
    wire new_AGEMA_signal_28333 ;
    wire new_AGEMA_signal_28334 ;
    wire new_AGEMA_signal_28335 ;
    wire new_AGEMA_signal_28336 ;
    wire new_AGEMA_signal_28337 ;
    wire new_AGEMA_signal_28338 ;
    wire new_AGEMA_signal_28339 ;
    wire new_AGEMA_signal_28340 ;
    wire new_AGEMA_signal_28341 ;
    wire new_AGEMA_signal_28342 ;
    wire new_AGEMA_signal_28343 ;
    wire new_AGEMA_signal_28344 ;
    wire new_AGEMA_signal_28345 ;
    wire new_AGEMA_signal_28346 ;
    wire new_AGEMA_signal_28347 ;
    wire new_AGEMA_signal_28348 ;
    wire new_AGEMA_signal_28349 ;
    wire new_AGEMA_signal_28350 ;
    wire new_AGEMA_signal_28351 ;
    wire new_AGEMA_signal_28352 ;
    wire new_AGEMA_signal_28353 ;
    wire new_AGEMA_signal_28354 ;
    wire new_AGEMA_signal_28355 ;
    wire new_AGEMA_signal_28356 ;
    wire new_AGEMA_signal_28357 ;
    wire new_AGEMA_signal_28358 ;
    wire new_AGEMA_signal_28359 ;
    wire new_AGEMA_signal_28360 ;
    wire new_AGEMA_signal_28361 ;
    wire new_AGEMA_signal_28362 ;
    wire new_AGEMA_signal_28363 ;
    wire new_AGEMA_signal_28364 ;
    wire new_AGEMA_signal_28365 ;
    wire new_AGEMA_signal_28366 ;
    wire new_AGEMA_signal_28367 ;
    wire new_AGEMA_signal_28368 ;
    wire new_AGEMA_signal_28369 ;
    wire new_AGEMA_signal_28370 ;
    wire new_AGEMA_signal_28371 ;
    wire new_AGEMA_signal_28372 ;
    wire new_AGEMA_signal_28373 ;
    wire new_AGEMA_signal_28374 ;
    wire new_AGEMA_signal_28375 ;
    wire new_AGEMA_signal_28376 ;
    wire new_AGEMA_signal_28377 ;
    wire new_AGEMA_signal_28378 ;
    wire new_AGEMA_signal_28379 ;
    wire new_AGEMA_signal_28380 ;
    wire new_AGEMA_signal_28381 ;
    wire new_AGEMA_signal_28382 ;
    wire new_AGEMA_signal_28383 ;
    wire new_AGEMA_signal_28384 ;
    wire new_AGEMA_signal_28385 ;
    wire new_AGEMA_signal_28386 ;
    wire new_AGEMA_signal_28387 ;
    wire new_AGEMA_signal_28388 ;
    wire new_AGEMA_signal_28389 ;
    wire new_AGEMA_signal_28390 ;
    wire new_AGEMA_signal_28391 ;
    wire new_AGEMA_signal_28392 ;
    wire new_AGEMA_signal_28393 ;
    wire new_AGEMA_signal_28394 ;
    wire new_AGEMA_signal_28395 ;
    wire new_AGEMA_signal_28396 ;
    wire new_AGEMA_signal_28397 ;
    wire new_AGEMA_signal_28398 ;
    wire new_AGEMA_signal_28399 ;
    wire new_AGEMA_signal_28400 ;
    wire new_AGEMA_signal_28401 ;
    wire new_AGEMA_signal_28402 ;
    wire new_AGEMA_signal_28403 ;
    wire new_AGEMA_signal_28404 ;
    wire new_AGEMA_signal_28405 ;
    wire new_AGEMA_signal_28406 ;
    wire new_AGEMA_signal_28407 ;
    wire new_AGEMA_signal_28408 ;
    wire new_AGEMA_signal_28409 ;
    wire new_AGEMA_signal_28410 ;
    wire new_AGEMA_signal_28411 ;
    wire new_AGEMA_signal_28412 ;
    wire new_AGEMA_signal_28413 ;
    wire new_AGEMA_signal_28414 ;
    wire new_AGEMA_signal_28415 ;
    wire new_AGEMA_signal_28416 ;
    wire new_AGEMA_signal_28417 ;
    wire new_AGEMA_signal_28418 ;
    wire new_AGEMA_signal_28419 ;
    wire new_AGEMA_signal_28420 ;
    wire new_AGEMA_signal_28421 ;
    wire new_AGEMA_signal_28422 ;
    wire new_AGEMA_signal_28423 ;
    wire new_AGEMA_signal_28424 ;
    wire new_AGEMA_signal_28425 ;
    wire new_AGEMA_signal_28426 ;
    wire new_AGEMA_signal_28427 ;
    wire new_AGEMA_signal_28428 ;
    wire new_AGEMA_signal_28429 ;
    wire new_AGEMA_signal_28430 ;
    wire new_AGEMA_signal_28431 ;
    wire new_AGEMA_signal_28432 ;
    wire new_AGEMA_signal_28433 ;
    wire new_AGEMA_signal_28434 ;
    wire new_AGEMA_signal_28435 ;
    wire new_AGEMA_signal_28436 ;
    wire new_AGEMA_signal_28437 ;
    wire new_AGEMA_signal_28438 ;
    wire new_AGEMA_signal_28439 ;
    wire new_AGEMA_signal_28440 ;
    wire new_AGEMA_signal_28441 ;
    wire new_AGEMA_signal_28442 ;
    wire new_AGEMA_signal_28443 ;
    wire new_AGEMA_signal_28444 ;
    wire new_AGEMA_signal_28445 ;
    wire new_AGEMA_signal_28446 ;
    wire new_AGEMA_signal_28447 ;
    wire new_AGEMA_signal_28448 ;
    wire new_AGEMA_signal_28449 ;
    wire new_AGEMA_signal_28450 ;
    wire new_AGEMA_signal_28451 ;
    wire new_AGEMA_signal_28452 ;
    wire new_AGEMA_signal_28453 ;
    wire new_AGEMA_signal_28454 ;
    wire new_AGEMA_signal_28455 ;
    wire new_AGEMA_signal_28456 ;
    wire new_AGEMA_signal_28457 ;
    wire new_AGEMA_signal_28458 ;
    wire new_AGEMA_signal_28459 ;
    wire new_AGEMA_signal_28460 ;
    wire new_AGEMA_signal_28461 ;
    wire new_AGEMA_signal_28462 ;
    wire new_AGEMA_signal_28463 ;
    wire new_AGEMA_signal_28464 ;
    wire new_AGEMA_signal_28465 ;
    wire new_AGEMA_signal_28466 ;
    wire new_AGEMA_signal_28467 ;
    wire new_AGEMA_signal_28468 ;
    wire new_AGEMA_signal_28469 ;
    wire new_AGEMA_signal_28470 ;
    wire new_AGEMA_signal_28471 ;
    wire new_AGEMA_signal_28472 ;
    wire new_AGEMA_signal_28473 ;
    wire new_AGEMA_signal_28474 ;
    wire new_AGEMA_signal_28475 ;
    wire new_AGEMA_signal_28476 ;
    wire new_AGEMA_signal_28477 ;
    wire new_AGEMA_signal_28478 ;
    wire new_AGEMA_signal_28479 ;
    wire new_AGEMA_signal_28480 ;
    wire new_AGEMA_signal_28481 ;
    wire new_AGEMA_signal_28482 ;
    wire new_AGEMA_signal_28483 ;
    wire new_AGEMA_signal_28484 ;
    wire new_AGEMA_signal_28485 ;
    wire new_AGEMA_signal_28486 ;
    wire new_AGEMA_signal_28487 ;
    wire new_AGEMA_signal_28488 ;
    wire new_AGEMA_signal_28489 ;
    wire new_AGEMA_signal_28490 ;
    wire new_AGEMA_signal_28491 ;
    wire new_AGEMA_signal_28492 ;
    wire new_AGEMA_signal_28493 ;
    wire new_AGEMA_signal_28494 ;
    wire new_AGEMA_signal_28495 ;
    wire new_AGEMA_signal_28496 ;
    wire new_AGEMA_signal_28497 ;
    wire new_AGEMA_signal_28498 ;
    wire new_AGEMA_signal_28499 ;
    wire new_AGEMA_signal_28500 ;
    wire new_AGEMA_signal_28501 ;
    wire new_AGEMA_signal_28502 ;
    wire new_AGEMA_signal_28503 ;
    wire new_AGEMA_signal_28504 ;
    wire new_AGEMA_signal_28505 ;
    wire new_AGEMA_signal_28506 ;
    wire new_AGEMA_signal_28507 ;
    wire new_AGEMA_signal_28508 ;
    wire new_AGEMA_signal_28509 ;
    wire new_AGEMA_signal_28510 ;
    wire new_AGEMA_signal_28511 ;
    wire new_AGEMA_signal_28512 ;
    wire new_AGEMA_signal_28513 ;
    wire new_AGEMA_signal_28514 ;
    wire new_AGEMA_signal_28515 ;
    wire new_AGEMA_signal_28516 ;
    wire new_AGEMA_signal_28517 ;
    wire new_AGEMA_signal_28518 ;
    wire new_AGEMA_signal_28519 ;
    wire new_AGEMA_signal_28520 ;
    wire new_AGEMA_signal_28521 ;
    wire new_AGEMA_signal_28522 ;
    wire new_AGEMA_signal_28523 ;
    wire new_AGEMA_signal_28524 ;
    wire new_AGEMA_signal_28525 ;
    wire new_AGEMA_signal_28526 ;
    wire new_AGEMA_signal_28527 ;
    wire new_AGEMA_signal_28528 ;
    wire new_AGEMA_signal_28529 ;
    wire new_AGEMA_signal_28530 ;
    wire new_AGEMA_signal_28531 ;
    wire new_AGEMA_signal_28532 ;
    wire new_AGEMA_signal_28533 ;
    wire new_AGEMA_signal_28534 ;
    wire new_AGEMA_signal_28535 ;
    wire new_AGEMA_signal_28536 ;
    wire new_AGEMA_signal_28537 ;
    wire new_AGEMA_signal_28538 ;
    wire new_AGEMA_signal_28539 ;
    wire new_AGEMA_signal_28540 ;
    wire new_AGEMA_signal_28541 ;
    wire new_AGEMA_signal_28542 ;
    wire new_AGEMA_signal_28543 ;
    wire new_AGEMA_signal_28544 ;
    wire new_AGEMA_signal_28545 ;
    wire new_AGEMA_signal_28546 ;
    wire new_AGEMA_signal_28547 ;
    wire new_AGEMA_signal_28548 ;
    wire new_AGEMA_signal_28549 ;
    wire new_AGEMA_signal_28550 ;
    wire new_AGEMA_signal_28551 ;
    wire new_AGEMA_signal_28552 ;
    wire new_AGEMA_signal_28553 ;
    wire new_AGEMA_signal_28554 ;
    wire new_AGEMA_signal_28555 ;
    wire new_AGEMA_signal_28556 ;
    wire new_AGEMA_signal_28557 ;
    wire new_AGEMA_signal_28558 ;
    wire new_AGEMA_signal_28559 ;
    wire new_AGEMA_signal_28560 ;
    wire new_AGEMA_signal_28561 ;
    wire new_AGEMA_signal_28562 ;
    wire new_AGEMA_signal_28563 ;
    wire new_AGEMA_signal_28564 ;
    wire new_AGEMA_signal_28565 ;
    wire new_AGEMA_signal_28566 ;
    wire new_AGEMA_signal_28567 ;
    wire new_AGEMA_signal_28568 ;
    wire new_AGEMA_signal_28569 ;
    wire new_AGEMA_signal_28570 ;
    wire new_AGEMA_signal_28571 ;
    wire new_AGEMA_signal_28572 ;
    wire new_AGEMA_signal_28573 ;
    wire new_AGEMA_signal_28574 ;
    wire new_AGEMA_signal_28575 ;
    wire new_AGEMA_signal_28576 ;
    wire new_AGEMA_signal_28577 ;
    wire new_AGEMA_signal_28578 ;
    wire new_AGEMA_signal_28579 ;
    wire new_AGEMA_signal_28580 ;
    wire new_AGEMA_signal_28581 ;
    wire new_AGEMA_signal_28582 ;
    wire new_AGEMA_signal_28583 ;
    wire new_AGEMA_signal_28584 ;
    wire new_AGEMA_signal_28585 ;
    wire new_AGEMA_signal_28586 ;
    wire new_AGEMA_signal_28587 ;
    wire new_AGEMA_signal_28588 ;
    wire new_AGEMA_signal_28589 ;
    wire new_AGEMA_signal_28590 ;
    wire new_AGEMA_signal_28591 ;
    wire new_AGEMA_signal_28592 ;
    wire new_AGEMA_signal_28593 ;
    wire new_AGEMA_signal_28594 ;
    wire new_AGEMA_signal_28595 ;
    wire new_AGEMA_signal_28596 ;
    wire new_AGEMA_signal_28597 ;
    wire new_AGEMA_signal_28598 ;
    wire new_AGEMA_signal_28599 ;
    wire new_AGEMA_signal_28600 ;
    wire new_AGEMA_signal_28601 ;
    wire new_AGEMA_signal_28602 ;
    wire new_AGEMA_signal_28603 ;
    wire new_AGEMA_signal_28604 ;
    wire new_AGEMA_signal_28605 ;
    wire new_AGEMA_signal_28606 ;
    wire new_AGEMA_signal_28607 ;
    wire new_AGEMA_signal_28608 ;
    wire new_AGEMA_signal_28609 ;
    wire new_AGEMA_signal_28610 ;
    wire new_AGEMA_signal_28611 ;
    wire new_AGEMA_signal_28612 ;
    wire new_AGEMA_signal_28613 ;
    wire new_AGEMA_signal_28614 ;
    wire new_AGEMA_signal_28615 ;
    wire new_AGEMA_signal_28616 ;
    wire new_AGEMA_signal_28617 ;
    wire new_AGEMA_signal_28618 ;
    wire new_AGEMA_signal_28619 ;
    wire new_AGEMA_signal_28620 ;
    wire new_AGEMA_signal_28621 ;
    wire new_AGEMA_signal_28622 ;
    wire new_AGEMA_signal_28623 ;
    wire new_AGEMA_signal_28624 ;
    wire new_AGEMA_signal_28625 ;
    wire new_AGEMA_signal_28626 ;
    wire new_AGEMA_signal_28627 ;
    wire new_AGEMA_signal_28628 ;
    wire new_AGEMA_signal_28629 ;
    wire new_AGEMA_signal_28630 ;
    wire new_AGEMA_signal_28631 ;
    wire new_AGEMA_signal_28632 ;
    wire new_AGEMA_signal_28633 ;
    wire new_AGEMA_signal_28634 ;
    wire new_AGEMA_signal_28635 ;
    wire new_AGEMA_signal_28636 ;
    wire new_AGEMA_signal_28637 ;
    wire new_AGEMA_signal_28638 ;
    wire new_AGEMA_signal_28639 ;
    wire new_AGEMA_signal_28640 ;
    wire new_AGEMA_signal_28641 ;
    wire new_AGEMA_signal_28642 ;
    wire new_AGEMA_signal_28643 ;
    wire new_AGEMA_signal_28644 ;
    wire new_AGEMA_signal_28645 ;
    wire new_AGEMA_signal_28646 ;
    wire new_AGEMA_signal_28647 ;
    wire new_AGEMA_signal_28648 ;
    wire new_AGEMA_signal_28649 ;
    wire new_AGEMA_signal_28650 ;
    wire new_AGEMA_signal_28651 ;
    wire new_AGEMA_signal_28652 ;
    wire new_AGEMA_signal_28653 ;
    wire new_AGEMA_signal_28654 ;
    wire new_AGEMA_signal_28655 ;
    wire new_AGEMA_signal_28656 ;
    wire new_AGEMA_signal_28657 ;
    wire new_AGEMA_signal_28658 ;
    wire new_AGEMA_signal_28659 ;
    wire new_AGEMA_signal_28660 ;
    wire new_AGEMA_signal_28661 ;
    wire new_AGEMA_signal_28662 ;
    wire new_AGEMA_signal_28663 ;
    wire new_AGEMA_signal_28664 ;
    wire new_AGEMA_signal_28665 ;
    wire new_AGEMA_signal_28666 ;
    wire new_AGEMA_signal_28667 ;
    wire new_AGEMA_signal_28668 ;
    wire new_AGEMA_signal_28669 ;
    wire new_AGEMA_signal_28670 ;
    wire new_AGEMA_signal_28671 ;
    wire new_AGEMA_signal_28672 ;
    wire new_AGEMA_signal_28673 ;
    wire new_AGEMA_signal_28674 ;
    wire new_AGEMA_signal_28675 ;
    wire new_AGEMA_signal_28676 ;
    wire new_AGEMA_signal_28677 ;
    wire new_AGEMA_signal_28678 ;
    wire new_AGEMA_signal_28679 ;
    wire new_AGEMA_signal_28680 ;
    wire new_AGEMA_signal_28681 ;
    wire new_AGEMA_signal_28682 ;
    wire new_AGEMA_signal_28683 ;
    wire new_AGEMA_signal_28684 ;
    wire new_AGEMA_signal_28685 ;
    wire new_AGEMA_signal_28686 ;
    wire new_AGEMA_signal_28687 ;
    wire new_AGEMA_signal_28688 ;
    wire new_AGEMA_signal_28689 ;
    wire new_AGEMA_signal_28690 ;
    wire new_AGEMA_signal_28691 ;
    wire new_AGEMA_signal_28692 ;
    wire new_AGEMA_signal_28693 ;
    wire new_AGEMA_signal_28694 ;
    wire new_AGEMA_signal_28695 ;
    wire new_AGEMA_signal_28696 ;
    wire new_AGEMA_signal_28697 ;
    wire new_AGEMA_signal_28698 ;
    wire new_AGEMA_signal_28699 ;
    wire new_AGEMA_signal_28700 ;
    wire new_AGEMA_signal_28701 ;
    wire new_AGEMA_signal_28702 ;
    wire new_AGEMA_signal_28703 ;
    wire new_AGEMA_signal_28704 ;
    wire new_AGEMA_signal_28705 ;
    wire new_AGEMA_signal_28706 ;
    wire new_AGEMA_signal_28707 ;
    wire new_AGEMA_signal_28708 ;
    wire new_AGEMA_signal_28709 ;
    wire new_AGEMA_signal_28710 ;
    wire new_AGEMA_signal_28711 ;
    wire new_AGEMA_signal_28712 ;
    wire new_AGEMA_signal_28713 ;
    wire new_AGEMA_signal_28714 ;
    wire new_AGEMA_signal_28715 ;
    wire new_AGEMA_signal_28716 ;
    wire new_AGEMA_signal_28717 ;
    wire new_AGEMA_signal_28718 ;
    wire new_AGEMA_signal_28719 ;
    wire new_AGEMA_signal_28720 ;
    wire new_AGEMA_signal_28721 ;
    wire new_AGEMA_signal_28722 ;
    wire new_AGEMA_signal_28723 ;
    wire new_AGEMA_signal_28724 ;
    wire new_AGEMA_signal_28725 ;
    wire new_AGEMA_signal_28726 ;
    wire new_AGEMA_signal_28727 ;
    wire new_AGEMA_signal_28728 ;
    wire new_AGEMA_signal_28729 ;
    wire new_AGEMA_signal_28730 ;
    wire new_AGEMA_signal_28731 ;
    wire new_AGEMA_signal_28732 ;
    wire new_AGEMA_signal_28733 ;
    wire new_AGEMA_signal_28734 ;
    wire new_AGEMA_signal_28735 ;
    wire new_AGEMA_signal_28736 ;
    wire new_AGEMA_signal_28737 ;
    wire new_AGEMA_signal_28738 ;
    wire new_AGEMA_signal_28739 ;
    wire new_AGEMA_signal_28740 ;
    wire new_AGEMA_signal_28741 ;
    wire new_AGEMA_signal_28742 ;
    wire new_AGEMA_signal_28743 ;
    wire new_AGEMA_signal_28744 ;
    wire new_AGEMA_signal_28745 ;
    wire new_AGEMA_signal_28746 ;
    wire new_AGEMA_signal_28747 ;
    wire new_AGEMA_signal_28748 ;
    wire new_AGEMA_signal_28749 ;
    wire new_AGEMA_signal_28750 ;
    wire new_AGEMA_signal_28751 ;
    wire new_AGEMA_signal_28752 ;
    wire new_AGEMA_signal_28753 ;
    wire new_AGEMA_signal_28754 ;
    wire new_AGEMA_signal_28755 ;
    wire new_AGEMA_signal_28756 ;
    wire new_AGEMA_signal_28757 ;
    wire new_AGEMA_signal_28758 ;
    wire new_AGEMA_signal_28759 ;
    wire new_AGEMA_signal_28760 ;
    wire new_AGEMA_signal_28761 ;
    wire new_AGEMA_signal_28762 ;
    wire new_AGEMA_signal_28763 ;
    wire new_AGEMA_signal_28764 ;
    wire new_AGEMA_signal_28765 ;
    wire new_AGEMA_signal_28766 ;
    wire new_AGEMA_signal_28767 ;
    wire new_AGEMA_signal_28768 ;
    wire new_AGEMA_signal_28769 ;
    wire new_AGEMA_signal_28770 ;
    wire new_AGEMA_signal_28771 ;
    wire new_AGEMA_signal_28772 ;
    wire new_AGEMA_signal_28773 ;
    wire new_AGEMA_signal_28774 ;
    wire new_AGEMA_signal_28775 ;
    wire new_AGEMA_signal_28776 ;
    wire new_AGEMA_signal_28777 ;
    wire new_AGEMA_signal_28778 ;
    wire new_AGEMA_signal_28779 ;
    wire new_AGEMA_signal_28780 ;
    wire new_AGEMA_signal_28781 ;
    wire new_AGEMA_signal_28782 ;
    wire new_AGEMA_signal_28783 ;
    wire new_AGEMA_signal_28784 ;
    wire new_AGEMA_signal_28785 ;
    wire new_AGEMA_signal_28786 ;
    wire new_AGEMA_signal_28787 ;
    wire new_AGEMA_signal_28788 ;
    wire new_AGEMA_signal_28789 ;
    wire new_AGEMA_signal_28790 ;
    wire new_AGEMA_signal_28791 ;
    wire new_AGEMA_signal_28792 ;
    wire new_AGEMA_signal_28793 ;
    wire new_AGEMA_signal_28794 ;
    wire new_AGEMA_signal_28795 ;
    wire new_AGEMA_signal_28796 ;
    wire new_AGEMA_signal_28797 ;
    wire new_AGEMA_signal_28798 ;
    wire new_AGEMA_signal_28799 ;
    wire new_AGEMA_signal_28800 ;
    wire new_AGEMA_signal_28801 ;
    wire new_AGEMA_signal_28802 ;
    wire new_AGEMA_signal_28803 ;
    wire new_AGEMA_signal_28804 ;
    wire new_AGEMA_signal_28805 ;
    wire new_AGEMA_signal_28806 ;
    wire new_AGEMA_signal_28807 ;
    wire new_AGEMA_signal_28808 ;
    wire new_AGEMA_signal_28809 ;
    wire new_AGEMA_signal_28810 ;
    wire new_AGEMA_signal_28811 ;
    wire new_AGEMA_signal_28812 ;
    wire new_AGEMA_signal_28813 ;
    wire new_AGEMA_signal_28814 ;
    wire new_AGEMA_signal_28815 ;
    wire new_AGEMA_signal_28816 ;
    wire new_AGEMA_signal_28817 ;
    wire new_AGEMA_signal_28818 ;
    wire new_AGEMA_signal_28819 ;
    wire new_AGEMA_signal_28820 ;
    wire new_AGEMA_signal_28821 ;
    wire new_AGEMA_signal_28822 ;
    wire new_AGEMA_signal_28823 ;
    wire new_AGEMA_signal_28824 ;
    wire new_AGEMA_signal_28825 ;
    wire new_AGEMA_signal_28826 ;
    wire new_AGEMA_signal_28827 ;
    wire new_AGEMA_signal_28828 ;
    wire new_AGEMA_signal_28829 ;
    wire new_AGEMA_signal_28830 ;
    wire new_AGEMA_signal_28831 ;
    wire new_AGEMA_signal_28832 ;
    wire new_AGEMA_signal_28833 ;
    wire new_AGEMA_signal_28834 ;
    wire new_AGEMA_signal_28835 ;
    wire new_AGEMA_signal_28836 ;
    wire new_AGEMA_signal_28837 ;
    wire new_AGEMA_signal_28838 ;
    wire new_AGEMA_signal_28839 ;
    wire new_AGEMA_signal_28840 ;
    wire new_AGEMA_signal_28841 ;
    wire new_AGEMA_signal_28842 ;
    wire new_AGEMA_signal_28843 ;
    wire new_AGEMA_signal_28844 ;
    wire new_AGEMA_signal_28845 ;
    wire new_AGEMA_signal_28846 ;
    wire new_AGEMA_signal_28847 ;
    wire new_AGEMA_signal_28848 ;
    wire new_AGEMA_signal_28849 ;
    wire new_AGEMA_signal_28850 ;
    wire new_AGEMA_signal_28851 ;
    wire new_AGEMA_signal_28852 ;
    wire new_AGEMA_signal_28853 ;
    wire new_AGEMA_signal_28854 ;
    wire new_AGEMA_signal_28855 ;
    wire new_AGEMA_signal_28856 ;
    wire new_AGEMA_signal_28857 ;
    wire new_AGEMA_signal_28858 ;
    wire new_AGEMA_signal_28859 ;
    wire new_AGEMA_signal_28860 ;
    wire new_AGEMA_signal_28861 ;
    wire new_AGEMA_signal_28862 ;
    wire new_AGEMA_signal_28863 ;
    wire new_AGEMA_signal_28864 ;
    wire new_AGEMA_signal_28865 ;
    wire new_AGEMA_signal_28866 ;
    wire new_AGEMA_signal_28867 ;
    wire new_AGEMA_signal_28868 ;
    wire new_AGEMA_signal_28869 ;
    wire new_AGEMA_signal_28870 ;
    wire new_AGEMA_signal_28871 ;
    wire new_AGEMA_signal_28872 ;
    wire new_AGEMA_signal_28873 ;
    wire new_AGEMA_signal_28874 ;
    wire new_AGEMA_signal_28875 ;
    wire new_AGEMA_signal_28876 ;
    wire new_AGEMA_signal_28877 ;
    wire new_AGEMA_signal_28878 ;
    wire new_AGEMA_signal_28879 ;
    wire new_AGEMA_signal_28880 ;
    wire new_AGEMA_signal_28881 ;
    wire new_AGEMA_signal_28882 ;
    wire new_AGEMA_signal_28883 ;
    wire new_AGEMA_signal_28884 ;
    wire new_AGEMA_signal_28885 ;
    wire new_AGEMA_signal_28886 ;
    wire new_AGEMA_signal_28887 ;
    wire new_AGEMA_signal_28888 ;
    wire new_AGEMA_signal_28889 ;
    wire new_AGEMA_signal_28890 ;
    wire new_AGEMA_signal_28891 ;
    wire new_AGEMA_signal_28892 ;
    wire new_AGEMA_signal_28893 ;
    wire new_AGEMA_signal_28894 ;
    wire new_AGEMA_signal_28895 ;
    wire new_AGEMA_signal_28896 ;
    wire new_AGEMA_signal_28897 ;
    wire new_AGEMA_signal_28898 ;
    wire new_AGEMA_signal_28899 ;
    wire new_AGEMA_signal_28900 ;
    wire new_AGEMA_signal_28901 ;
    wire new_AGEMA_signal_28902 ;
    wire new_AGEMA_signal_28903 ;
    wire new_AGEMA_signal_28904 ;
    wire new_AGEMA_signal_28905 ;
    wire new_AGEMA_signal_28906 ;
    wire new_AGEMA_signal_28907 ;
    wire new_AGEMA_signal_28908 ;
    wire new_AGEMA_signal_28909 ;
    wire new_AGEMA_signal_28910 ;
    wire new_AGEMA_signal_28911 ;
    wire new_AGEMA_signal_28912 ;
    wire new_AGEMA_signal_28913 ;
    wire new_AGEMA_signal_28914 ;
    wire new_AGEMA_signal_28915 ;
    wire new_AGEMA_signal_28916 ;
    wire new_AGEMA_signal_28917 ;
    wire new_AGEMA_signal_28918 ;
    wire new_AGEMA_signal_28919 ;
    wire new_AGEMA_signal_28920 ;
    wire new_AGEMA_signal_28921 ;
    wire new_AGEMA_signal_28922 ;
    wire new_AGEMA_signal_28923 ;
    wire new_AGEMA_signal_28924 ;
    wire new_AGEMA_signal_28925 ;
    wire new_AGEMA_signal_28926 ;
    wire new_AGEMA_signal_28927 ;
    wire new_AGEMA_signal_28928 ;
    wire new_AGEMA_signal_28929 ;
    wire new_AGEMA_signal_28930 ;
    wire new_AGEMA_signal_28931 ;
    wire new_AGEMA_signal_28932 ;
    wire new_AGEMA_signal_28933 ;
    wire new_AGEMA_signal_28934 ;
    wire new_AGEMA_signal_28935 ;
    wire new_AGEMA_signal_28936 ;
    wire new_AGEMA_signal_28937 ;
    wire new_AGEMA_signal_28938 ;
    wire new_AGEMA_signal_28939 ;
    wire new_AGEMA_signal_28940 ;
    wire new_AGEMA_signal_28941 ;
    wire new_AGEMA_signal_28942 ;
    wire new_AGEMA_signal_28943 ;
    wire new_AGEMA_signal_28944 ;
    wire new_AGEMA_signal_28945 ;
    wire new_AGEMA_signal_28946 ;
    wire new_AGEMA_signal_28947 ;
    wire new_AGEMA_signal_28948 ;
    wire new_AGEMA_signal_28949 ;
    wire new_AGEMA_signal_28950 ;
    wire new_AGEMA_signal_28951 ;
    wire new_AGEMA_signal_28952 ;
    wire new_AGEMA_signal_28953 ;
    wire new_AGEMA_signal_28954 ;
    wire new_AGEMA_signal_28955 ;
    wire new_AGEMA_signal_28956 ;
    wire new_AGEMA_signal_28957 ;
    wire new_AGEMA_signal_28958 ;
    wire new_AGEMA_signal_28959 ;
    wire new_AGEMA_signal_28960 ;
    wire new_AGEMA_signal_28961 ;
    wire new_AGEMA_signal_28962 ;
    wire new_AGEMA_signal_28963 ;
    wire new_AGEMA_signal_28964 ;
    wire new_AGEMA_signal_28965 ;
    wire new_AGEMA_signal_28966 ;
    wire new_AGEMA_signal_28967 ;
    wire new_AGEMA_signal_28968 ;
    wire new_AGEMA_signal_28969 ;
    wire new_AGEMA_signal_28970 ;
    wire new_AGEMA_signal_28971 ;
    wire new_AGEMA_signal_28972 ;
    wire new_AGEMA_signal_28973 ;
    wire new_AGEMA_signal_28974 ;
    wire new_AGEMA_signal_28975 ;
    wire new_AGEMA_signal_28976 ;
    wire new_AGEMA_signal_28977 ;
    wire new_AGEMA_signal_28978 ;
    wire new_AGEMA_signal_28979 ;
    wire new_AGEMA_signal_28980 ;
    wire new_AGEMA_signal_28981 ;
    wire new_AGEMA_signal_28982 ;
    wire new_AGEMA_signal_28983 ;
    wire new_AGEMA_signal_28984 ;
    wire new_AGEMA_signal_28985 ;
    wire new_AGEMA_signal_28986 ;
    wire new_AGEMA_signal_28987 ;
    wire new_AGEMA_signal_28988 ;
    wire new_AGEMA_signal_28989 ;
    wire new_AGEMA_signal_28990 ;
    wire new_AGEMA_signal_28991 ;
    wire new_AGEMA_signal_28992 ;
    wire new_AGEMA_signal_28993 ;
    wire new_AGEMA_signal_28994 ;
    wire new_AGEMA_signal_28995 ;
    wire new_AGEMA_signal_28996 ;
    wire new_AGEMA_signal_28997 ;
    wire new_AGEMA_signal_28998 ;
    wire new_AGEMA_signal_28999 ;
    wire new_AGEMA_signal_29000 ;
    wire new_AGEMA_signal_29001 ;
    wire new_AGEMA_signal_29002 ;
    wire new_AGEMA_signal_29003 ;
    wire new_AGEMA_signal_29004 ;
    wire new_AGEMA_signal_29005 ;
    wire new_AGEMA_signal_29006 ;
    wire new_AGEMA_signal_29007 ;
    wire new_AGEMA_signal_29008 ;
    wire new_AGEMA_signal_29009 ;
    wire new_AGEMA_signal_29010 ;
    wire new_AGEMA_signal_29011 ;
    wire new_AGEMA_signal_29012 ;
    wire new_AGEMA_signal_29013 ;
    wire new_AGEMA_signal_29014 ;
    wire new_AGEMA_signal_29015 ;
    wire new_AGEMA_signal_29016 ;
    wire new_AGEMA_signal_29017 ;
    wire new_AGEMA_signal_29018 ;
    wire new_AGEMA_signal_29019 ;
    wire new_AGEMA_signal_29020 ;
    wire new_AGEMA_signal_29021 ;
    wire new_AGEMA_signal_29022 ;
    wire new_AGEMA_signal_29023 ;
    wire new_AGEMA_signal_29024 ;
    wire new_AGEMA_signal_29025 ;
    wire new_AGEMA_signal_29026 ;
    wire new_AGEMA_signal_29027 ;
    wire new_AGEMA_signal_29028 ;
    wire new_AGEMA_signal_29029 ;
    wire new_AGEMA_signal_29030 ;
    wire new_AGEMA_signal_29031 ;
    wire new_AGEMA_signal_29032 ;
    wire new_AGEMA_signal_29033 ;
    wire new_AGEMA_signal_29034 ;
    wire new_AGEMA_signal_29035 ;
    wire new_AGEMA_signal_29036 ;
    wire new_AGEMA_signal_29037 ;
    wire new_AGEMA_signal_29038 ;
    wire new_AGEMA_signal_29039 ;
    wire new_AGEMA_signal_29040 ;
    wire new_AGEMA_signal_29041 ;
    wire new_AGEMA_signal_29042 ;
    wire new_AGEMA_signal_29043 ;
    wire new_AGEMA_signal_29044 ;
    wire new_AGEMA_signal_29045 ;
    wire new_AGEMA_signal_29046 ;
    wire new_AGEMA_signal_29047 ;
    wire new_AGEMA_signal_29048 ;
    wire new_AGEMA_signal_29049 ;
    wire new_AGEMA_signal_29050 ;
    wire new_AGEMA_signal_29051 ;
    wire new_AGEMA_signal_29052 ;
    wire new_AGEMA_signal_29053 ;
    wire new_AGEMA_signal_29054 ;
    wire new_AGEMA_signal_29055 ;
    wire new_AGEMA_signal_29056 ;
    wire new_AGEMA_signal_29057 ;
    wire new_AGEMA_signal_29058 ;
    wire new_AGEMA_signal_29059 ;
    wire new_AGEMA_signal_29060 ;
    wire new_AGEMA_signal_29061 ;
    wire new_AGEMA_signal_29062 ;
    wire new_AGEMA_signal_29063 ;
    wire new_AGEMA_signal_29064 ;
    wire new_AGEMA_signal_29065 ;
    wire new_AGEMA_signal_29066 ;
    wire new_AGEMA_signal_29067 ;
    wire new_AGEMA_signal_29068 ;
    wire new_AGEMA_signal_29069 ;
    wire new_AGEMA_signal_29070 ;
    wire new_AGEMA_signal_29071 ;
    wire new_AGEMA_signal_29072 ;
    wire new_AGEMA_signal_29073 ;
    wire new_AGEMA_signal_29074 ;
    wire new_AGEMA_signal_29075 ;
    wire new_AGEMA_signal_29076 ;
    wire new_AGEMA_signal_29077 ;
    wire new_AGEMA_signal_29078 ;
    wire new_AGEMA_signal_29079 ;
    wire new_AGEMA_signal_29080 ;
    wire new_AGEMA_signal_29081 ;
    wire new_AGEMA_signal_29082 ;
    wire new_AGEMA_signal_29083 ;
    wire new_AGEMA_signal_29084 ;
    wire new_AGEMA_signal_29085 ;
    wire new_AGEMA_signal_29086 ;
    wire new_AGEMA_signal_29087 ;
    wire new_AGEMA_signal_29088 ;
    wire new_AGEMA_signal_29089 ;
    wire new_AGEMA_signal_29090 ;
    wire new_AGEMA_signal_29091 ;
    wire new_AGEMA_signal_29092 ;
    wire new_AGEMA_signal_29093 ;
    wire new_AGEMA_signal_29094 ;
    wire new_AGEMA_signal_29095 ;
    wire new_AGEMA_signal_29096 ;
    wire new_AGEMA_signal_29097 ;
    wire new_AGEMA_signal_29098 ;
    wire new_AGEMA_signal_29099 ;
    wire new_AGEMA_signal_29100 ;
    wire new_AGEMA_signal_29101 ;
    wire new_AGEMA_signal_29102 ;
    wire new_AGEMA_signal_29103 ;
    wire new_AGEMA_signal_29104 ;
    wire new_AGEMA_signal_29105 ;
    wire new_AGEMA_signal_29106 ;
    wire new_AGEMA_signal_29107 ;
    wire new_AGEMA_signal_29108 ;
    wire new_AGEMA_signal_29109 ;
    wire new_AGEMA_signal_29110 ;
    wire new_AGEMA_signal_29111 ;
    wire new_AGEMA_signal_29112 ;
    wire new_AGEMA_signal_29113 ;
    wire new_AGEMA_signal_29114 ;
    wire new_AGEMA_signal_29115 ;
    wire new_AGEMA_signal_29116 ;
    wire new_AGEMA_signal_29117 ;
    wire new_AGEMA_signal_29118 ;
    wire new_AGEMA_signal_29119 ;
    wire new_AGEMA_signal_29120 ;
    wire new_AGEMA_signal_29121 ;
    wire new_AGEMA_signal_29122 ;
    wire new_AGEMA_signal_29123 ;
    wire new_AGEMA_signal_29124 ;
    wire new_AGEMA_signal_29125 ;
    wire new_AGEMA_signal_29126 ;
    wire new_AGEMA_signal_29127 ;
    wire new_AGEMA_signal_29128 ;
    wire new_AGEMA_signal_29129 ;
    wire new_AGEMA_signal_29130 ;
    wire new_AGEMA_signal_29131 ;
    wire new_AGEMA_signal_29132 ;
    wire new_AGEMA_signal_29133 ;
    wire new_AGEMA_signal_29134 ;
    wire new_AGEMA_signal_29135 ;
    wire new_AGEMA_signal_29136 ;
    wire new_AGEMA_signal_29137 ;
    wire new_AGEMA_signal_29138 ;
    wire new_AGEMA_signal_29139 ;
    wire new_AGEMA_signal_29140 ;
    wire new_AGEMA_signal_29141 ;
    wire new_AGEMA_signal_29142 ;
    wire new_AGEMA_signal_29143 ;
    wire new_AGEMA_signal_29144 ;
    wire new_AGEMA_signal_29145 ;
    wire new_AGEMA_signal_29146 ;
    wire new_AGEMA_signal_29147 ;
    wire new_AGEMA_signal_29148 ;
    wire new_AGEMA_signal_29149 ;
    wire new_AGEMA_signal_29150 ;
    wire new_AGEMA_signal_29151 ;
    wire new_AGEMA_signal_29152 ;
    wire new_AGEMA_signal_29153 ;
    wire new_AGEMA_signal_29154 ;
    wire new_AGEMA_signal_29155 ;
    wire new_AGEMA_signal_29156 ;
    wire new_AGEMA_signal_29157 ;
    wire new_AGEMA_signal_29158 ;
    wire new_AGEMA_signal_29159 ;
    wire new_AGEMA_signal_29160 ;
    wire new_AGEMA_signal_29161 ;
    wire new_AGEMA_signal_29162 ;
    wire new_AGEMA_signal_29163 ;
    wire new_AGEMA_signal_29164 ;
    wire new_AGEMA_signal_29165 ;
    wire new_AGEMA_signal_29166 ;
    wire new_AGEMA_signal_29167 ;
    wire new_AGEMA_signal_29168 ;
    wire new_AGEMA_signal_29169 ;
    wire new_AGEMA_signal_29170 ;
    wire new_AGEMA_signal_29171 ;
    wire new_AGEMA_signal_29172 ;
    wire new_AGEMA_signal_29173 ;
    wire new_AGEMA_signal_29174 ;
    wire new_AGEMA_signal_29175 ;
    wire new_AGEMA_signal_29176 ;
    wire new_AGEMA_signal_29177 ;
    wire new_AGEMA_signal_29178 ;
    wire new_AGEMA_signal_29179 ;
    wire new_AGEMA_signal_29180 ;
    wire new_AGEMA_signal_29181 ;
    wire new_AGEMA_signal_29182 ;
    wire new_AGEMA_signal_29183 ;
    wire new_AGEMA_signal_29184 ;
    wire new_AGEMA_signal_29185 ;
    wire new_AGEMA_signal_29186 ;
    wire new_AGEMA_signal_29187 ;
    wire new_AGEMA_signal_29188 ;
    wire new_AGEMA_signal_29189 ;
    wire new_AGEMA_signal_29190 ;
    wire new_AGEMA_signal_29191 ;
    wire new_AGEMA_signal_29192 ;
    wire new_AGEMA_signal_29193 ;
    wire new_AGEMA_signal_29194 ;
    wire new_AGEMA_signal_29195 ;
    wire new_AGEMA_signal_29196 ;
    wire new_AGEMA_signal_29197 ;
    wire new_AGEMA_signal_29198 ;
    wire new_AGEMA_signal_29199 ;
    wire new_AGEMA_signal_29200 ;
    wire new_AGEMA_signal_29201 ;
    wire new_AGEMA_signal_29202 ;
    wire new_AGEMA_signal_29203 ;
    wire new_AGEMA_signal_29204 ;
    wire new_AGEMA_signal_29205 ;
    wire new_AGEMA_signal_29206 ;
    wire new_AGEMA_signal_29207 ;
    wire new_AGEMA_signal_29208 ;
    wire new_AGEMA_signal_29209 ;
    wire new_AGEMA_signal_29210 ;
    wire new_AGEMA_signal_29211 ;
    wire new_AGEMA_signal_29212 ;
    wire new_AGEMA_signal_29213 ;
    wire new_AGEMA_signal_29214 ;
    wire new_AGEMA_signal_29215 ;
    wire new_AGEMA_signal_29216 ;
    wire new_AGEMA_signal_29217 ;
    wire new_AGEMA_signal_29218 ;
    wire new_AGEMA_signal_29219 ;
    wire new_AGEMA_signal_29220 ;
    wire new_AGEMA_signal_29221 ;
    wire new_AGEMA_signal_29222 ;
    wire new_AGEMA_signal_29223 ;
    wire new_AGEMA_signal_29224 ;
    wire new_AGEMA_signal_29225 ;
    wire new_AGEMA_signal_29226 ;
    wire new_AGEMA_signal_29227 ;
    wire new_AGEMA_signal_29228 ;
    wire new_AGEMA_signal_29229 ;
    wire new_AGEMA_signal_29230 ;
    wire new_AGEMA_signal_29231 ;
    wire new_AGEMA_signal_29232 ;
    wire new_AGEMA_signal_29233 ;
    wire new_AGEMA_signal_29234 ;
    wire new_AGEMA_signal_29235 ;
    wire new_AGEMA_signal_29236 ;
    wire new_AGEMA_signal_29237 ;
    wire new_AGEMA_signal_29238 ;
    wire new_AGEMA_signal_29239 ;
    wire new_AGEMA_signal_29240 ;
    wire new_AGEMA_signal_29241 ;
    wire new_AGEMA_signal_29242 ;
    wire new_AGEMA_signal_29243 ;
    wire new_AGEMA_signal_29244 ;
    wire new_AGEMA_signal_29245 ;
    wire new_AGEMA_signal_29246 ;
    wire new_AGEMA_signal_29247 ;
    wire new_AGEMA_signal_29248 ;
    wire new_AGEMA_signal_29249 ;
    wire new_AGEMA_signal_29250 ;
    wire new_AGEMA_signal_29251 ;
    wire new_AGEMA_signal_29252 ;
    wire new_AGEMA_signal_29253 ;
    wire new_AGEMA_signal_29254 ;
    wire new_AGEMA_signal_29255 ;
    wire new_AGEMA_signal_29256 ;
    wire new_AGEMA_signal_29257 ;
    wire new_AGEMA_signal_29258 ;
    wire new_AGEMA_signal_29259 ;
    wire new_AGEMA_signal_29260 ;
    wire new_AGEMA_signal_29261 ;
    wire new_AGEMA_signal_29262 ;
    wire new_AGEMA_signal_29263 ;
    wire new_AGEMA_signal_29264 ;
    wire new_AGEMA_signal_29265 ;
    wire new_AGEMA_signal_29266 ;
    wire new_AGEMA_signal_29267 ;
    wire new_AGEMA_signal_29268 ;
    wire new_AGEMA_signal_29269 ;
    wire new_AGEMA_signal_29270 ;
    wire new_AGEMA_signal_29271 ;
    wire new_AGEMA_signal_29272 ;
    wire new_AGEMA_signal_29273 ;
    wire new_AGEMA_signal_29274 ;
    wire new_AGEMA_signal_29275 ;
    wire new_AGEMA_signal_29276 ;
    wire new_AGEMA_signal_29277 ;
    wire new_AGEMA_signal_29278 ;
    wire new_AGEMA_signal_29279 ;
    wire new_AGEMA_signal_29280 ;
    wire new_AGEMA_signal_29281 ;
    wire new_AGEMA_signal_29282 ;
    wire new_AGEMA_signal_29283 ;
    wire new_AGEMA_signal_29284 ;
    wire new_AGEMA_signal_29285 ;
    wire new_AGEMA_signal_29286 ;
    wire new_AGEMA_signal_29287 ;
    wire new_AGEMA_signal_29288 ;
    wire new_AGEMA_signal_29289 ;
    wire new_AGEMA_signal_29290 ;
    wire new_AGEMA_signal_29291 ;
    wire new_AGEMA_signal_29292 ;
    wire new_AGEMA_signal_29293 ;
    wire new_AGEMA_signal_29294 ;
    wire new_AGEMA_signal_29295 ;
    wire new_AGEMA_signal_29296 ;
    wire new_AGEMA_signal_29297 ;
    wire new_AGEMA_signal_29298 ;
    wire new_AGEMA_signal_29299 ;
    wire new_AGEMA_signal_29300 ;
    wire new_AGEMA_signal_29301 ;
    wire new_AGEMA_signal_29302 ;
    wire new_AGEMA_signal_29303 ;
    wire new_AGEMA_signal_29304 ;
    wire new_AGEMA_signal_29305 ;
    wire new_AGEMA_signal_29306 ;
    wire new_AGEMA_signal_29307 ;
    wire new_AGEMA_signal_29308 ;
    wire new_AGEMA_signal_29309 ;
    wire new_AGEMA_signal_29310 ;
    wire new_AGEMA_signal_29311 ;
    wire new_AGEMA_signal_29312 ;
    wire new_AGEMA_signal_29313 ;
    wire new_AGEMA_signal_29314 ;
    wire new_AGEMA_signal_29315 ;
    wire new_AGEMA_signal_29316 ;
    wire new_AGEMA_signal_29317 ;
    wire new_AGEMA_signal_29318 ;
    wire new_AGEMA_signal_29319 ;
    wire new_AGEMA_signal_29320 ;
    wire new_AGEMA_signal_29321 ;
    wire new_AGEMA_signal_29322 ;
    wire new_AGEMA_signal_29323 ;
    wire new_AGEMA_signal_29324 ;
    wire new_AGEMA_signal_29325 ;
    wire new_AGEMA_signal_29326 ;
    wire new_AGEMA_signal_29327 ;
    wire new_AGEMA_signal_29328 ;
    wire new_AGEMA_signal_29329 ;
    wire new_AGEMA_signal_29330 ;
    wire new_AGEMA_signal_29331 ;
    wire new_AGEMA_signal_29332 ;
    wire new_AGEMA_signal_29333 ;
    wire new_AGEMA_signal_29334 ;
    wire new_AGEMA_signal_29335 ;
    wire new_AGEMA_signal_29336 ;
    wire new_AGEMA_signal_29337 ;
    wire new_AGEMA_signal_29338 ;
    wire new_AGEMA_signal_29339 ;
    wire new_AGEMA_signal_29340 ;
    wire new_AGEMA_signal_29341 ;
    wire new_AGEMA_signal_29342 ;
    wire new_AGEMA_signal_29343 ;
    wire new_AGEMA_signal_29344 ;
    wire new_AGEMA_signal_29345 ;
    wire new_AGEMA_signal_29346 ;
    wire new_AGEMA_signal_29347 ;
    wire new_AGEMA_signal_29348 ;
    wire new_AGEMA_signal_29349 ;
    wire new_AGEMA_signal_29350 ;
    wire new_AGEMA_signal_29351 ;
    wire new_AGEMA_signal_29352 ;
    wire new_AGEMA_signal_29353 ;
    wire new_AGEMA_signal_29354 ;
    wire new_AGEMA_signal_29355 ;
    wire new_AGEMA_signal_29356 ;
    wire new_AGEMA_signal_29357 ;
    wire new_AGEMA_signal_29358 ;
    wire new_AGEMA_signal_29359 ;
    wire new_AGEMA_signal_29360 ;
    wire new_AGEMA_signal_29361 ;
    wire new_AGEMA_signal_29362 ;
    wire new_AGEMA_signal_29363 ;
    wire new_AGEMA_signal_29364 ;
    wire new_AGEMA_signal_29365 ;
    wire new_AGEMA_signal_29366 ;
    wire new_AGEMA_signal_29367 ;
    wire new_AGEMA_signal_29368 ;
    wire new_AGEMA_signal_29369 ;
    wire new_AGEMA_signal_29370 ;
    wire new_AGEMA_signal_29371 ;
    wire new_AGEMA_signal_29372 ;
    wire new_AGEMA_signal_29373 ;
    wire new_AGEMA_signal_29374 ;
    wire new_AGEMA_signal_29375 ;
    wire new_AGEMA_signal_29376 ;
    wire new_AGEMA_signal_29377 ;
    wire new_AGEMA_signal_29378 ;
    wire new_AGEMA_signal_29379 ;
    wire new_AGEMA_signal_29380 ;
    wire new_AGEMA_signal_29381 ;
    wire new_AGEMA_signal_29382 ;
    wire new_AGEMA_signal_29383 ;
    wire new_AGEMA_signal_29384 ;
    wire new_AGEMA_signal_29385 ;
    wire new_AGEMA_signal_29386 ;
    wire new_AGEMA_signal_29387 ;
    wire new_AGEMA_signal_29388 ;
    wire new_AGEMA_signal_29389 ;
    wire new_AGEMA_signal_29390 ;
    wire new_AGEMA_signal_29391 ;
    wire new_AGEMA_signal_29392 ;
    wire new_AGEMA_signal_29393 ;
    wire new_AGEMA_signal_29394 ;
    wire new_AGEMA_signal_29395 ;
    wire new_AGEMA_signal_29396 ;
    wire new_AGEMA_signal_29397 ;
    wire new_AGEMA_signal_29398 ;
    wire new_AGEMA_signal_29399 ;
    wire new_AGEMA_signal_29400 ;
    wire new_AGEMA_signal_29401 ;
    wire new_AGEMA_signal_29402 ;
    wire new_AGEMA_signal_29403 ;
    wire new_AGEMA_signal_29404 ;
    wire new_AGEMA_signal_29405 ;
    wire new_AGEMA_signal_29406 ;
    wire new_AGEMA_signal_29407 ;
    wire new_AGEMA_signal_29408 ;
    wire new_AGEMA_signal_29409 ;
    wire new_AGEMA_signal_29410 ;
    wire new_AGEMA_signal_29411 ;
    wire new_AGEMA_signal_29412 ;
    wire new_AGEMA_signal_29413 ;
    wire new_AGEMA_signal_29414 ;
    wire new_AGEMA_signal_29415 ;
    wire new_AGEMA_signal_29416 ;
    wire new_AGEMA_signal_29417 ;
    wire new_AGEMA_signal_29418 ;
    wire new_AGEMA_signal_29419 ;
    wire new_AGEMA_signal_29420 ;
    wire new_AGEMA_signal_29421 ;
    wire new_AGEMA_signal_29422 ;
    wire new_AGEMA_signal_29423 ;
    wire new_AGEMA_signal_29424 ;
    wire new_AGEMA_signal_29425 ;
    wire new_AGEMA_signal_29426 ;
    wire new_AGEMA_signal_29427 ;
    wire new_AGEMA_signal_29428 ;
    wire new_AGEMA_signal_29429 ;
    wire new_AGEMA_signal_29430 ;
    wire new_AGEMA_signal_29431 ;
    wire new_AGEMA_signal_29432 ;
    wire new_AGEMA_signal_29433 ;
    wire new_AGEMA_signal_29434 ;
    wire new_AGEMA_signal_29435 ;
    wire new_AGEMA_signal_29436 ;
    wire new_AGEMA_signal_29437 ;
    wire new_AGEMA_signal_29438 ;
    wire new_AGEMA_signal_29439 ;
    wire new_AGEMA_signal_29440 ;
    wire new_AGEMA_signal_29441 ;
    wire new_AGEMA_signal_29442 ;
    wire new_AGEMA_signal_29443 ;
    wire new_AGEMA_signal_29444 ;
    wire new_AGEMA_signal_29445 ;
    wire new_AGEMA_signal_29446 ;
    wire new_AGEMA_signal_29447 ;
    wire new_AGEMA_signal_29448 ;
    wire new_AGEMA_signal_29449 ;
    wire new_AGEMA_signal_29450 ;
    wire new_AGEMA_signal_29451 ;
    wire new_AGEMA_signal_29452 ;
    wire new_AGEMA_signal_29453 ;
    wire new_AGEMA_signal_29454 ;
    wire new_AGEMA_signal_29455 ;
    wire new_AGEMA_signal_29456 ;
    wire new_AGEMA_signal_29457 ;
    wire new_AGEMA_signal_29458 ;
    wire new_AGEMA_signal_29459 ;
    wire new_AGEMA_signal_29460 ;
    wire new_AGEMA_signal_29461 ;
    wire new_AGEMA_signal_29462 ;
    wire new_AGEMA_signal_29463 ;
    wire new_AGEMA_signal_29464 ;
    wire new_AGEMA_signal_29465 ;
    wire new_AGEMA_signal_29466 ;
    wire new_AGEMA_signal_29467 ;
    wire new_AGEMA_signal_29468 ;
    wire new_AGEMA_signal_29469 ;
    wire new_AGEMA_signal_29470 ;
    wire new_AGEMA_signal_29471 ;
    wire new_AGEMA_signal_29472 ;
    wire new_AGEMA_signal_29473 ;
    wire new_AGEMA_signal_29474 ;
    wire new_AGEMA_signal_29475 ;
    wire new_AGEMA_signal_29476 ;
    wire new_AGEMA_signal_29477 ;
    wire new_AGEMA_signal_29478 ;
    wire new_AGEMA_signal_29479 ;
    wire new_AGEMA_signal_29480 ;
    wire new_AGEMA_signal_29481 ;
    wire new_AGEMA_signal_29482 ;
    wire new_AGEMA_signal_29483 ;
    wire new_AGEMA_signal_29484 ;
    wire new_AGEMA_signal_29485 ;
    wire new_AGEMA_signal_29486 ;
    wire new_AGEMA_signal_29487 ;
    wire new_AGEMA_signal_29488 ;
    wire new_AGEMA_signal_29489 ;
    wire new_AGEMA_signal_29490 ;
    wire new_AGEMA_signal_29491 ;
    wire new_AGEMA_signal_29492 ;
    wire new_AGEMA_signal_29493 ;
    wire new_AGEMA_signal_29494 ;
    wire new_AGEMA_signal_29495 ;
    wire new_AGEMA_signal_29496 ;
    wire new_AGEMA_signal_29497 ;
    wire new_AGEMA_signal_29498 ;
    wire new_AGEMA_signal_29499 ;
    wire new_AGEMA_signal_29500 ;
    wire new_AGEMA_signal_29501 ;
    wire new_AGEMA_signal_29502 ;
    wire new_AGEMA_signal_29503 ;
    wire new_AGEMA_signal_29504 ;
    wire new_AGEMA_signal_29505 ;
    wire new_AGEMA_signal_29506 ;
    wire new_AGEMA_signal_29507 ;
    wire new_AGEMA_signal_29508 ;
    wire new_AGEMA_signal_29509 ;
    wire new_AGEMA_signal_29510 ;
    wire new_AGEMA_signal_29511 ;
    wire new_AGEMA_signal_29512 ;
    wire new_AGEMA_signal_29513 ;
    wire new_AGEMA_signal_29514 ;
    wire new_AGEMA_signal_29515 ;
    wire new_AGEMA_signal_29516 ;
    wire new_AGEMA_signal_29517 ;
    wire new_AGEMA_signal_29518 ;
    wire new_AGEMA_signal_29519 ;
    wire new_AGEMA_signal_29520 ;
    wire new_AGEMA_signal_29521 ;
    wire new_AGEMA_signal_29522 ;
    wire new_AGEMA_signal_29523 ;
    wire new_AGEMA_signal_29524 ;
    wire new_AGEMA_signal_29525 ;
    wire new_AGEMA_signal_29526 ;
    wire new_AGEMA_signal_29527 ;
    wire new_AGEMA_signal_29528 ;
    wire new_AGEMA_signal_29529 ;
    wire new_AGEMA_signal_29530 ;
    wire new_AGEMA_signal_29531 ;
    wire new_AGEMA_signal_29532 ;
    wire new_AGEMA_signal_29533 ;
    wire new_AGEMA_signal_29534 ;
    wire new_AGEMA_signal_29535 ;
    wire new_AGEMA_signal_29536 ;
    wire new_AGEMA_signal_29537 ;
    wire new_AGEMA_signal_29538 ;
    wire new_AGEMA_signal_29539 ;
    wire new_AGEMA_signal_29540 ;
    wire new_AGEMA_signal_29541 ;
    wire new_AGEMA_signal_29542 ;
    wire new_AGEMA_signal_29543 ;
    wire new_AGEMA_signal_29544 ;
    wire new_AGEMA_signal_29545 ;
    wire new_AGEMA_signal_29546 ;
    wire new_AGEMA_signal_29547 ;
    wire new_AGEMA_signal_29548 ;
    wire new_AGEMA_signal_29549 ;
    wire new_AGEMA_signal_29550 ;
    wire new_AGEMA_signal_29551 ;
    wire new_AGEMA_signal_29552 ;
    wire new_AGEMA_signal_29553 ;
    wire new_AGEMA_signal_29554 ;
    wire new_AGEMA_signal_29555 ;
    wire new_AGEMA_signal_29556 ;
    wire new_AGEMA_signal_29557 ;
    wire new_AGEMA_signal_29558 ;
    wire new_AGEMA_signal_29559 ;
    wire new_AGEMA_signal_29560 ;
    wire new_AGEMA_signal_29561 ;
    wire new_AGEMA_signal_29562 ;
    wire new_AGEMA_signal_29563 ;
    wire new_AGEMA_signal_29564 ;
    wire new_AGEMA_signal_29565 ;
    wire new_AGEMA_signal_29566 ;
    wire new_AGEMA_signal_29567 ;
    wire new_AGEMA_signal_29568 ;
    wire new_AGEMA_signal_29569 ;
    wire new_AGEMA_signal_29570 ;
    wire new_AGEMA_signal_29571 ;
    wire new_AGEMA_signal_29572 ;
    wire new_AGEMA_signal_29573 ;
    wire new_AGEMA_signal_29574 ;
    wire new_AGEMA_signal_29575 ;
    wire new_AGEMA_signal_29576 ;
    wire new_AGEMA_signal_29577 ;
    wire new_AGEMA_signal_29578 ;
    wire new_AGEMA_signal_29579 ;
    wire new_AGEMA_signal_29580 ;
    wire new_AGEMA_signal_29581 ;
    wire new_AGEMA_signal_29582 ;
    wire new_AGEMA_signal_29583 ;
    wire new_AGEMA_signal_29584 ;
    wire new_AGEMA_signal_29585 ;
    wire new_AGEMA_signal_29586 ;
    wire new_AGEMA_signal_29587 ;
    wire new_AGEMA_signal_29588 ;
    wire new_AGEMA_signal_29589 ;
    wire new_AGEMA_signal_29590 ;
    wire new_AGEMA_signal_29591 ;
    wire new_AGEMA_signal_29592 ;
    wire new_AGEMA_signal_29593 ;
    wire new_AGEMA_signal_29594 ;
    wire new_AGEMA_signal_29595 ;
    wire new_AGEMA_signal_29596 ;
    wire new_AGEMA_signal_29597 ;
    wire new_AGEMA_signal_29598 ;
    wire new_AGEMA_signal_29599 ;
    wire new_AGEMA_signal_29600 ;
    wire new_AGEMA_signal_29601 ;
    wire new_AGEMA_signal_29602 ;
    wire new_AGEMA_signal_29603 ;
    wire new_AGEMA_signal_29604 ;
    wire new_AGEMA_signal_29605 ;
    wire new_AGEMA_signal_29606 ;
    wire new_AGEMA_signal_29607 ;
    wire new_AGEMA_signal_29608 ;
    wire new_AGEMA_signal_29609 ;
    wire new_AGEMA_signal_29610 ;
    wire new_AGEMA_signal_29611 ;
    wire new_AGEMA_signal_29612 ;
    wire new_AGEMA_signal_29613 ;
    wire new_AGEMA_signal_29614 ;
    wire new_AGEMA_signal_29615 ;
    wire new_AGEMA_signal_29616 ;
    wire new_AGEMA_signal_29617 ;
    wire new_AGEMA_signal_29618 ;
    wire new_AGEMA_signal_29619 ;
    wire new_AGEMA_signal_29620 ;
    wire new_AGEMA_signal_29621 ;
    wire new_AGEMA_signal_29622 ;
    wire new_AGEMA_signal_29623 ;
    wire new_AGEMA_signal_29624 ;
    wire new_AGEMA_signal_29625 ;
    wire new_AGEMA_signal_29626 ;
    wire new_AGEMA_signal_29627 ;
    wire new_AGEMA_signal_29628 ;
    wire new_AGEMA_signal_29629 ;
    wire new_AGEMA_signal_29630 ;
    wire new_AGEMA_signal_29631 ;
    wire new_AGEMA_signal_29632 ;
    wire new_AGEMA_signal_29633 ;
    wire new_AGEMA_signal_29634 ;
    wire new_AGEMA_signal_29635 ;
    wire new_AGEMA_signal_29636 ;
    wire new_AGEMA_signal_29637 ;
    wire new_AGEMA_signal_29638 ;
    wire new_AGEMA_signal_29639 ;
    wire new_AGEMA_signal_29640 ;
    wire new_AGEMA_signal_29641 ;
    wire new_AGEMA_signal_29642 ;
    wire new_AGEMA_signal_29643 ;
    wire new_AGEMA_signal_29644 ;
    wire new_AGEMA_signal_29645 ;
    wire new_AGEMA_signal_29646 ;
    wire new_AGEMA_signal_29647 ;
    wire new_AGEMA_signal_29648 ;
    wire new_AGEMA_signal_29649 ;
    wire new_AGEMA_signal_29650 ;
    wire new_AGEMA_signal_29651 ;
    wire new_AGEMA_signal_29652 ;
    wire new_AGEMA_signal_29653 ;
    wire new_AGEMA_signal_29654 ;
    wire new_AGEMA_signal_29655 ;
    wire new_AGEMA_signal_29656 ;
    wire new_AGEMA_signal_29657 ;
    wire new_AGEMA_signal_29658 ;
    wire new_AGEMA_signal_29659 ;
    wire new_AGEMA_signal_29660 ;
    wire new_AGEMA_signal_29661 ;
    wire new_AGEMA_signal_29662 ;
    wire new_AGEMA_signal_29663 ;
    wire new_AGEMA_signal_29664 ;
    wire new_AGEMA_signal_29665 ;
    wire new_AGEMA_signal_29666 ;
    wire new_AGEMA_signal_29667 ;
    wire new_AGEMA_signal_29668 ;
    wire new_AGEMA_signal_29669 ;
    wire new_AGEMA_signal_29670 ;
    wire new_AGEMA_signal_29671 ;
    wire new_AGEMA_signal_29672 ;
    wire new_AGEMA_signal_29673 ;
    wire new_AGEMA_signal_29674 ;
    wire new_AGEMA_signal_29675 ;
    wire new_AGEMA_signal_29676 ;
    wire new_AGEMA_signal_29677 ;
    wire new_AGEMA_signal_29678 ;
    wire new_AGEMA_signal_29679 ;
    wire new_AGEMA_signal_29680 ;
    wire new_AGEMA_signal_29681 ;
    wire new_AGEMA_signal_29682 ;
    wire new_AGEMA_signal_29683 ;
    wire new_AGEMA_signal_29684 ;
    wire new_AGEMA_signal_29685 ;
    wire new_AGEMA_signal_29686 ;
    wire new_AGEMA_signal_29687 ;
    wire new_AGEMA_signal_29688 ;
    wire new_AGEMA_signal_29689 ;
    wire new_AGEMA_signal_29690 ;
    wire new_AGEMA_signal_29691 ;
    wire new_AGEMA_signal_29692 ;
    wire new_AGEMA_signal_29693 ;
    wire new_AGEMA_signal_29694 ;
    wire new_AGEMA_signal_29695 ;
    wire new_AGEMA_signal_29696 ;
    wire new_AGEMA_signal_29697 ;
    wire new_AGEMA_signal_29698 ;
    wire new_AGEMA_signal_29699 ;
    wire new_AGEMA_signal_29700 ;
    wire new_AGEMA_signal_29701 ;
    wire new_AGEMA_signal_29702 ;
    wire new_AGEMA_signal_29703 ;
    wire new_AGEMA_signal_29704 ;
    wire new_AGEMA_signal_29705 ;
    wire new_AGEMA_signal_29706 ;
    wire new_AGEMA_signal_29707 ;
    wire new_AGEMA_signal_29708 ;
    wire new_AGEMA_signal_29709 ;
    wire new_AGEMA_signal_29710 ;
    wire new_AGEMA_signal_29711 ;
    wire new_AGEMA_signal_29712 ;
    wire new_AGEMA_signal_29713 ;
    wire new_AGEMA_signal_29714 ;
    wire new_AGEMA_signal_29715 ;
    wire new_AGEMA_signal_29716 ;
    wire new_AGEMA_signal_29717 ;
    wire new_AGEMA_signal_29718 ;
    wire new_AGEMA_signal_29719 ;
    wire new_AGEMA_signal_29720 ;
    wire new_AGEMA_signal_29721 ;
    wire new_AGEMA_signal_29722 ;
    wire new_AGEMA_signal_29723 ;
    wire new_AGEMA_signal_29724 ;
    wire new_AGEMA_signal_29725 ;
    wire new_AGEMA_signal_29726 ;
    wire new_AGEMA_signal_29727 ;
    wire new_AGEMA_signal_29728 ;
    wire new_AGEMA_signal_29729 ;
    wire new_AGEMA_signal_29730 ;
    wire new_AGEMA_signal_29731 ;
    wire new_AGEMA_signal_29732 ;
    wire new_AGEMA_signal_29733 ;
    wire new_AGEMA_signal_29734 ;
    wire new_AGEMA_signal_29735 ;
    wire new_AGEMA_signal_29736 ;
    wire new_AGEMA_signal_29737 ;
    wire new_AGEMA_signal_29738 ;
    wire new_AGEMA_signal_29739 ;
    wire new_AGEMA_signal_29740 ;
    wire new_AGEMA_signal_29741 ;
    wire new_AGEMA_signal_29742 ;
    wire new_AGEMA_signal_29743 ;
    wire new_AGEMA_signal_29744 ;
    wire new_AGEMA_signal_29745 ;
    wire new_AGEMA_signal_29746 ;
    wire new_AGEMA_signal_29747 ;
    wire new_AGEMA_signal_29748 ;
    wire new_AGEMA_signal_29749 ;
    wire new_AGEMA_signal_29750 ;
    wire new_AGEMA_signal_29751 ;
    wire new_AGEMA_signal_29752 ;
    wire new_AGEMA_signal_29753 ;
    wire new_AGEMA_signal_29754 ;
    wire new_AGEMA_signal_29755 ;
    wire new_AGEMA_signal_29756 ;
    wire new_AGEMA_signal_29757 ;
    wire new_AGEMA_signal_29758 ;
    wire new_AGEMA_signal_29759 ;
    wire new_AGEMA_signal_29760 ;
    wire new_AGEMA_signal_29761 ;
    wire new_AGEMA_signal_29762 ;
    wire new_AGEMA_signal_29763 ;
    wire new_AGEMA_signal_29764 ;
    wire new_AGEMA_signal_29765 ;
    wire new_AGEMA_signal_29766 ;
    wire new_AGEMA_signal_29767 ;
    wire new_AGEMA_signal_29768 ;
    wire new_AGEMA_signal_29769 ;
    wire new_AGEMA_signal_29770 ;
    wire new_AGEMA_signal_29771 ;
    wire new_AGEMA_signal_29772 ;
    wire new_AGEMA_signal_29773 ;
    wire new_AGEMA_signal_29774 ;
    wire new_AGEMA_signal_29775 ;
    wire new_AGEMA_signal_29776 ;
    wire new_AGEMA_signal_29777 ;
    wire new_AGEMA_signal_29778 ;
    wire new_AGEMA_signal_29779 ;
    wire new_AGEMA_signal_29780 ;
    wire new_AGEMA_signal_29781 ;
    wire new_AGEMA_signal_29782 ;
    wire new_AGEMA_signal_29783 ;
    wire new_AGEMA_signal_29784 ;
    wire new_AGEMA_signal_29785 ;
    wire new_AGEMA_signal_29786 ;
    wire new_AGEMA_signal_29787 ;
    wire new_AGEMA_signal_29788 ;
    wire new_AGEMA_signal_29789 ;
    wire new_AGEMA_signal_29790 ;
    wire new_AGEMA_signal_29791 ;
    wire new_AGEMA_signal_29792 ;
    wire new_AGEMA_signal_29793 ;
    wire new_AGEMA_signal_29794 ;
    wire new_AGEMA_signal_29795 ;
    wire new_AGEMA_signal_29796 ;
    wire new_AGEMA_signal_29797 ;
    wire new_AGEMA_signal_29798 ;
    wire new_AGEMA_signal_29799 ;
    wire new_AGEMA_signal_29800 ;
    wire new_AGEMA_signal_29801 ;
    wire new_AGEMA_signal_29802 ;
    wire new_AGEMA_signal_29803 ;
    wire new_AGEMA_signal_29804 ;
    wire new_AGEMA_signal_29805 ;
    wire new_AGEMA_signal_29806 ;
    wire new_AGEMA_signal_29807 ;
    wire new_AGEMA_signal_29808 ;
    wire new_AGEMA_signal_29809 ;
    wire new_AGEMA_signal_29810 ;
    wire new_AGEMA_signal_29811 ;
    wire new_AGEMA_signal_29812 ;
    wire new_AGEMA_signal_29813 ;
    wire new_AGEMA_signal_29814 ;
    wire new_AGEMA_signal_29815 ;
    wire new_AGEMA_signal_29816 ;
    wire new_AGEMA_signal_29817 ;
    wire new_AGEMA_signal_29818 ;
    wire new_AGEMA_signal_29819 ;
    wire new_AGEMA_signal_29820 ;
    wire new_AGEMA_signal_29821 ;
    wire new_AGEMA_signal_29822 ;
    wire new_AGEMA_signal_29823 ;
    wire new_AGEMA_signal_29824 ;
    wire new_AGEMA_signal_29825 ;
    wire new_AGEMA_signal_29826 ;
    wire new_AGEMA_signal_29827 ;
    wire new_AGEMA_signal_29828 ;
    wire new_AGEMA_signal_29829 ;
    wire new_AGEMA_signal_29830 ;
    wire new_AGEMA_signal_29831 ;
    wire new_AGEMA_signal_29832 ;
    wire new_AGEMA_signal_29833 ;
    wire new_AGEMA_signal_29834 ;
    wire new_AGEMA_signal_29835 ;
    wire new_AGEMA_signal_29836 ;
    wire new_AGEMA_signal_29837 ;
    wire new_AGEMA_signal_29838 ;
    wire new_AGEMA_signal_29839 ;
    wire new_AGEMA_signal_29840 ;
    wire new_AGEMA_signal_29841 ;
    wire new_AGEMA_signal_29842 ;
    wire new_AGEMA_signal_29843 ;
    wire new_AGEMA_signal_29844 ;
    wire new_AGEMA_signal_29845 ;
    wire new_AGEMA_signal_29846 ;
    wire new_AGEMA_signal_29847 ;
    wire new_AGEMA_signal_29848 ;
    wire new_AGEMA_signal_29849 ;
    wire new_AGEMA_signal_29850 ;
    wire new_AGEMA_signal_29851 ;
    wire new_AGEMA_signal_29852 ;
    wire new_AGEMA_signal_29853 ;
    wire new_AGEMA_signal_29854 ;
    wire new_AGEMA_signal_29855 ;
    wire new_AGEMA_signal_29856 ;
    wire new_AGEMA_signal_29857 ;
    wire new_AGEMA_signal_29858 ;
    wire new_AGEMA_signal_29859 ;
    wire new_AGEMA_signal_29860 ;
    wire new_AGEMA_signal_29861 ;
    wire new_AGEMA_signal_29862 ;
    wire new_AGEMA_signal_29863 ;
    wire new_AGEMA_signal_29864 ;
    wire new_AGEMA_signal_29865 ;
    wire new_AGEMA_signal_29866 ;
    wire new_AGEMA_signal_29867 ;
    wire new_AGEMA_signal_29868 ;
    wire new_AGEMA_signal_29869 ;
    wire new_AGEMA_signal_29870 ;
    wire new_AGEMA_signal_29871 ;
    wire new_AGEMA_signal_29872 ;
    wire new_AGEMA_signal_29873 ;
    wire new_AGEMA_signal_29874 ;
    wire new_AGEMA_signal_29875 ;
    wire new_AGEMA_signal_29876 ;
    wire new_AGEMA_signal_29877 ;
    wire new_AGEMA_signal_29878 ;
    wire new_AGEMA_signal_29879 ;
    wire new_AGEMA_signal_29880 ;
    wire new_AGEMA_signal_29881 ;
    wire new_AGEMA_signal_29882 ;
    wire new_AGEMA_signal_29883 ;
    wire new_AGEMA_signal_29884 ;
    wire new_AGEMA_signal_29885 ;
    wire new_AGEMA_signal_29886 ;
    wire new_AGEMA_signal_29887 ;
    wire new_AGEMA_signal_29888 ;
    wire new_AGEMA_signal_29889 ;
    wire new_AGEMA_signal_29890 ;
    wire new_AGEMA_signal_29891 ;
    wire new_AGEMA_signal_29892 ;
    wire new_AGEMA_signal_29893 ;
    wire new_AGEMA_signal_29894 ;
    wire new_AGEMA_signal_29895 ;
    wire new_AGEMA_signal_29896 ;
    wire new_AGEMA_signal_29897 ;
    wire new_AGEMA_signal_29898 ;
    wire new_AGEMA_signal_29899 ;
    wire new_AGEMA_signal_29900 ;
    wire new_AGEMA_signal_29901 ;
    wire new_AGEMA_signal_29902 ;
    wire new_AGEMA_signal_29903 ;
    wire new_AGEMA_signal_29904 ;
    wire new_AGEMA_signal_29905 ;
    wire new_AGEMA_signal_29906 ;
    wire new_AGEMA_signal_29907 ;
    wire new_AGEMA_signal_29908 ;
    wire new_AGEMA_signal_29909 ;
    wire new_AGEMA_signal_29910 ;
    wire new_AGEMA_signal_29911 ;
    wire new_AGEMA_signal_29912 ;
    wire new_AGEMA_signal_29913 ;
    wire new_AGEMA_signal_29914 ;
    wire new_AGEMA_signal_29915 ;
    wire new_AGEMA_signal_29916 ;
    wire new_AGEMA_signal_29917 ;
    wire new_AGEMA_signal_29918 ;
    wire new_AGEMA_signal_29919 ;
    wire new_AGEMA_signal_29920 ;
    wire new_AGEMA_signal_29921 ;
    wire new_AGEMA_signal_29922 ;
    wire new_AGEMA_signal_29923 ;
    wire new_AGEMA_signal_29924 ;
    wire new_AGEMA_signal_29925 ;
    wire new_AGEMA_signal_29926 ;
    wire new_AGEMA_signal_29927 ;
    wire new_AGEMA_signal_29928 ;
    wire new_AGEMA_signal_29929 ;
    wire new_AGEMA_signal_29930 ;
    wire new_AGEMA_signal_29931 ;
    wire new_AGEMA_signal_29932 ;
    wire new_AGEMA_signal_29933 ;
    wire new_AGEMA_signal_29934 ;
    wire new_AGEMA_signal_29935 ;
    wire new_AGEMA_signal_29936 ;
    wire new_AGEMA_signal_29937 ;
    wire new_AGEMA_signal_29938 ;
    wire new_AGEMA_signal_29939 ;
    wire new_AGEMA_signal_29940 ;
    wire new_AGEMA_signal_29941 ;
    wire new_AGEMA_signal_29942 ;
    wire new_AGEMA_signal_29943 ;
    wire new_AGEMA_signal_29944 ;
    wire new_AGEMA_signal_29945 ;
    wire new_AGEMA_signal_29946 ;
    wire new_AGEMA_signal_29947 ;
    wire new_AGEMA_signal_29948 ;
    wire new_AGEMA_signal_29949 ;
    wire new_AGEMA_signal_29950 ;
    wire new_AGEMA_signal_29951 ;
    wire new_AGEMA_signal_29952 ;
    wire new_AGEMA_signal_29953 ;
    wire new_AGEMA_signal_29954 ;
    wire new_AGEMA_signal_29955 ;
    wire new_AGEMA_signal_29956 ;
    wire new_AGEMA_signal_29957 ;
    wire new_AGEMA_signal_29958 ;
    wire new_AGEMA_signal_29959 ;
    wire new_AGEMA_signal_29960 ;
    wire new_AGEMA_signal_29961 ;
    wire new_AGEMA_signal_29962 ;
    wire new_AGEMA_signal_29963 ;
    wire new_AGEMA_signal_29964 ;
    wire new_AGEMA_signal_29965 ;
    wire new_AGEMA_signal_29966 ;
    wire new_AGEMA_signal_29967 ;
    wire new_AGEMA_signal_29968 ;
    wire new_AGEMA_signal_29969 ;
    wire new_AGEMA_signal_29970 ;
    wire new_AGEMA_signal_29971 ;
    wire new_AGEMA_signal_29972 ;
    wire new_AGEMA_signal_29973 ;
    wire new_AGEMA_signal_29974 ;
    wire new_AGEMA_signal_29975 ;
    wire new_AGEMA_signal_29976 ;
    wire new_AGEMA_signal_29977 ;
    wire new_AGEMA_signal_29978 ;
    wire new_AGEMA_signal_29979 ;
    wire new_AGEMA_signal_29980 ;
    wire new_AGEMA_signal_29981 ;
    wire new_AGEMA_signal_29982 ;
    wire new_AGEMA_signal_29983 ;
    wire new_AGEMA_signal_29984 ;
    wire new_AGEMA_signal_29985 ;
    wire new_AGEMA_signal_29986 ;
    wire new_AGEMA_signal_29987 ;
    wire new_AGEMA_signal_29988 ;
    wire new_AGEMA_signal_29989 ;
    wire new_AGEMA_signal_29990 ;
    wire new_AGEMA_signal_29991 ;
    wire new_AGEMA_signal_29992 ;
    wire new_AGEMA_signal_29993 ;
    wire new_AGEMA_signal_29994 ;
    wire new_AGEMA_signal_29995 ;
    wire new_AGEMA_signal_29996 ;
    wire new_AGEMA_signal_29997 ;
    wire new_AGEMA_signal_29998 ;
    wire new_AGEMA_signal_29999 ;
    wire new_AGEMA_signal_30000 ;
    wire new_AGEMA_signal_30001 ;
    wire new_AGEMA_signal_30002 ;
    wire new_AGEMA_signal_30003 ;
    wire new_AGEMA_signal_30004 ;
    wire new_AGEMA_signal_30005 ;
    wire new_AGEMA_signal_30006 ;
    wire new_AGEMA_signal_30007 ;
    wire new_AGEMA_signal_30008 ;
    wire new_AGEMA_signal_30009 ;
    wire new_AGEMA_signal_30010 ;
    wire new_AGEMA_signal_30011 ;
    wire new_AGEMA_signal_30012 ;
    wire new_AGEMA_signal_30013 ;
    wire new_AGEMA_signal_30014 ;
    wire new_AGEMA_signal_30015 ;
    wire new_AGEMA_signal_30016 ;
    wire new_AGEMA_signal_30017 ;
    wire new_AGEMA_signal_30018 ;
    wire new_AGEMA_signal_30019 ;
    wire new_AGEMA_signal_30020 ;
    wire new_AGEMA_signal_30021 ;
    wire new_AGEMA_signal_30022 ;
    wire new_AGEMA_signal_30023 ;
    wire new_AGEMA_signal_30024 ;
    wire new_AGEMA_signal_30025 ;
    wire new_AGEMA_signal_30026 ;
    wire new_AGEMA_signal_30027 ;
    wire new_AGEMA_signal_30028 ;
    wire new_AGEMA_signal_30029 ;
    wire new_AGEMA_signal_30030 ;
    wire new_AGEMA_signal_30031 ;
    wire new_AGEMA_signal_30032 ;
    wire new_AGEMA_signal_30033 ;
    wire new_AGEMA_signal_30034 ;
    wire new_AGEMA_signal_30035 ;
    wire new_AGEMA_signal_30036 ;
    wire new_AGEMA_signal_30037 ;
    wire new_AGEMA_signal_30038 ;
    wire new_AGEMA_signal_30039 ;
    wire new_AGEMA_signal_30040 ;
    wire new_AGEMA_signal_30041 ;
    wire new_AGEMA_signal_30042 ;
    wire new_AGEMA_signal_30043 ;
    wire new_AGEMA_signal_30044 ;
    wire new_AGEMA_signal_30045 ;
    wire new_AGEMA_signal_30046 ;
    wire new_AGEMA_signal_30047 ;
    wire new_AGEMA_signal_30048 ;
    wire new_AGEMA_signal_30049 ;
    wire new_AGEMA_signal_30050 ;
    wire new_AGEMA_signal_30051 ;
    wire new_AGEMA_signal_30052 ;
    wire new_AGEMA_signal_30053 ;
    wire new_AGEMA_signal_30054 ;
    wire new_AGEMA_signal_30055 ;
    wire new_AGEMA_signal_30056 ;
    wire new_AGEMA_signal_30057 ;
    wire new_AGEMA_signal_30058 ;
    wire new_AGEMA_signal_30059 ;
    wire new_AGEMA_signal_30060 ;
    wire new_AGEMA_signal_30061 ;
    wire new_AGEMA_signal_30062 ;
    wire new_AGEMA_signal_30063 ;
    wire new_AGEMA_signal_30064 ;
    wire new_AGEMA_signal_30065 ;
    wire new_AGEMA_signal_30066 ;
    wire new_AGEMA_signal_30067 ;
    wire new_AGEMA_signal_30068 ;
    wire new_AGEMA_signal_30069 ;
    wire new_AGEMA_signal_30070 ;
    wire new_AGEMA_signal_30071 ;
    wire new_AGEMA_signal_30072 ;
    wire new_AGEMA_signal_30073 ;
    wire new_AGEMA_signal_30074 ;
    wire new_AGEMA_signal_30075 ;
    wire new_AGEMA_signal_30076 ;
    wire new_AGEMA_signal_30077 ;
    wire new_AGEMA_signal_30078 ;
    wire new_AGEMA_signal_30079 ;
    wire new_AGEMA_signal_30080 ;
    wire new_AGEMA_signal_30081 ;
    wire new_AGEMA_signal_30082 ;
    wire new_AGEMA_signal_30083 ;
    wire new_AGEMA_signal_30084 ;
    wire new_AGEMA_signal_30085 ;
    wire new_AGEMA_signal_30086 ;
    wire new_AGEMA_signal_30087 ;
    wire new_AGEMA_signal_30088 ;
    wire new_AGEMA_signal_30089 ;
    wire new_AGEMA_signal_30090 ;
    wire new_AGEMA_signal_30091 ;
    wire new_AGEMA_signal_30092 ;
    wire new_AGEMA_signal_30093 ;
    wire new_AGEMA_signal_30094 ;
    wire new_AGEMA_signal_30095 ;
    wire new_AGEMA_signal_30096 ;
    wire new_AGEMA_signal_30097 ;
    wire new_AGEMA_signal_30098 ;
    wire new_AGEMA_signal_30099 ;
    wire new_AGEMA_signal_30100 ;
    wire new_AGEMA_signal_30101 ;
    wire new_AGEMA_signal_30102 ;
    wire new_AGEMA_signal_30103 ;
    wire new_AGEMA_signal_30104 ;
    wire new_AGEMA_signal_30105 ;
    wire new_AGEMA_signal_30106 ;
    wire new_AGEMA_signal_30107 ;
    wire new_AGEMA_signal_30108 ;
    wire new_AGEMA_signal_30109 ;
    wire new_AGEMA_signal_30110 ;
    wire new_AGEMA_signal_30111 ;
    wire new_AGEMA_signal_30112 ;
    wire new_AGEMA_signal_30113 ;
    wire new_AGEMA_signal_30114 ;
    wire new_AGEMA_signal_30115 ;
    wire new_AGEMA_signal_30116 ;
    wire new_AGEMA_signal_30117 ;
    wire new_AGEMA_signal_30118 ;
    wire new_AGEMA_signal_30119 ;
    wire new_AGEMA_signal_30120 ;
    wire new_AGEMA_signal_30121 ;
    wire new_AGEMA_signal_30122 ;
    wire new_AGEMA_signal_30123 ;
    wire new_AGEMA_signal_30124 ;
    wire new_AGEMA_signal_30125 ;
    wire new_AGEMA_signal_30126 ;
    wire new_AGEMA_signal_30127 ;
    wire new_AGEMA_signal_30128 ;
    wire new_AGEMA_signal_30129 ;
    wire new_AGEMA_signal_30130 ;
    wire new_AGEMA_signal_30131 ;
    wire new_AGEMA_signal_30132 ;
    wire new_AGEMA_signal_30133 ;
    wire new_AGEMA_signal_30134 ;
    wire new_AGEMA_signal_30135 ;
    wire new_AGEMA_signal_30136 ;
    wire new_AGEMA_signal_30137 ;
    wire new_AGEMA_signal_30138 ;
    wire new_AGEMA_signal_30139 ;
    wire new_AGEMA_signal_30140 ;
    wire new_AGEMA_signal_30141 ;
    wire new_AGEMA_signal_30142 ;
    wire new_AGEMA_signal_30143 ;
    wire new_AGEMA_signal_30144 ;
    wire new_AGEMA_signal_30145 ;
    wire new_AGEMA_signal_30146 ;
    wire new_AGEMA_signal_30147 ;
    wire new_AGEMA_signal_30148 ;
    wire new_AGEMA_signal_30149 ;
    wire new_AGEMA_signal_30150 ;
    wire new_AGEMA_signal_30151 ;
    wire new_AGEMA_signal_30152 ;
    wire new_AGEMA_signal_30153 ;
    wire new_AGEMA_signal_30154 ;
    wire new_AGEMA_signal_30155 ;
    wire new_AGEMA_signal_30156 ;
    wire new_AGEMA_signal_30157 ;
    wire new_AGEMA_signal_30158 ;
    wire new_AGEMA_signal_30159 ;
    wire new_AGEMA_signal_30160 ;
    wire new_AGEMA_signal_30161 ;
    wire new_AGEMA_signal_30162 ;
    wire new_AGEMA_signal_30163 ;
    wire new_AGEMA_signal_30164 ;
    wire new_AGEMA_signal_30165 ;
    wire new_AGEMA_signal_30166 ;
    wire new_AGEMA_signal_30167 ;
    wire new_AGEMA_signal_30168 ;
    wire new_AGEMA_signal_30169 ;
    wire new_AGEMA_signal_30170 ;
    wire new_AGEMA_signal_30171 ;
    wire new_AGEMA_signal_30172 ;
    wire new_AGEMA_signal_30173 ;
    wire new_AGEMA_signal_30174 ;
    wire new_AGEMA_signal_30175 ;
    wire new_AGEMA_signal_30176 ;
    wire new_AGEMA_signal_30177 ;
    wire new_AGEMA_signal_30178 ;
    wire new_AGEMA_signal_30179 ;
    wire new_AGEMA_signal_30180 ;
    wire new_AGEMA_signal_30181 ;
    wire new_AGEMA_signal_30182 ;
    wire new_AGEMA_signal_30183 ;
    wire new_AGEMA_signal_30184 ;
    wire new_AGEMA_signal_30185 ;
    wire new_AGEMA_signal_30186 ;
    wire new_AGEMA_signal_30187 ;
    wire new_AGEMA_signal_30188 ;
    wire new_AGEMA_signal_30189 ;
    wire new_AGEMA_signal_30190 ;
    wire new_AGEMA_signal_30191 ;
    wire new_AGEMA_signal_30192 ;
    wire new_AGEMA_signal_30193 ;
    wire new_AGEMA_signal_30194 ;
    wire new_AGEMA_signal_30195 ;
    wire new_AGEMA_signal_30196 ;
    wire new_AGEMA_signal_30197 ;
    wire new_AGEMA_signal_30198 ;
    wire new_AGEMA_signal_30199 ;
    wire new_AGEMA_signal_30200 ;
    wire new_AGEMA_signal_30201 ;
    wire new_AGEMA_signal_30202 ;
    wire new_AGEMA_signal_30203 ;
    wire new_AGEMA_signal_30204 ;
    wire new_AGEMA_signal_30205 ;
    wire new_AGEMA_signal_30206 ;
    wire new_AGEMA_signal_30207 ;
    wire new_AGEMA_signal_30208 ;
    wire new_AGEMA_signal_30209 ;
    wire new_AGEMA_signal_30210 ;
    wire new_AGEMA_signal_30211 ;
    wire new_AGEMA_signal_30212 ;
    wire new_AGEMA_signal_30213 ;
    wire new_AGEMA_signal_30214 ;
    wire new_AGEMA_signal_30215 ;
    wire new_AGEMA_signal_30216 ;
    wire new_AGEMA_signal_30217 ;
    wire new_AGEMA_signal_30218 ;
    wire new_AGEMA_signal_30219 ;
    wire new_AGEMA_signal_30220 ;
    wire new_AGEMA_signal_30221 ;
    wire new_AGEMA_signal_30222 ;
    wire new_AGEMA_signal_30223 ;
    wire new_AGEMA_signal_30224 ;
    wire new_AGEMA_signal_30225 ;
    wire new_AGEMA_signal_30226 ;
    wire new_AGEMA_signal_30227 ;
    wire new_AGEMA_signal_30228 ;
    wire new_AGEMA_signal_30229 ;
    wire new_AGEMA_signal_30230 ;
    wire new_AGEMA_signal_30231 ;
    wire new_AGEMA_signal_30232 ;
    wire new_AGEMA_signal_30233 ;
    wire new_AGEMA_signal_30234 ;
    wire new_AGEMA_signal_30235 ;
    wire new_AGEMA_signal_30236 ;
    wire new_AGEMA_signal_30237 ;
    wire new_AGEMA_signal_30238 ;
    wire new_AGEMA_signal_30239 ;
    wire new_AGEMA_signal_30240 ;
    wire new_AGEMA_signal_30241 ;
    wire new_AGEMA_signal_30242 ;
    wire new_AGEMA_signal_30243 ;
    wire new_AGEMA_signal_30244 ;
    wire new_AGEMA_signal_30245 ;
    wire new_AGEMA_signal_30246 ;
    wire new_AGEMA_signal_30247 ;
    wire new_AGEMA_signal_30248 ;
    wire new_AGEMA_signal_30249 ;
    wire new_AGEMA_signal_30250 ;
    wire new_AGEMA_signal_30251 ;
    wire new_AGEMA_signal_30252 ;
    wire new_AGEMA_signal_30253 ;
    wire new_AGEMA_signal_30254 ;
    wire new_AGEMA_signal_30255 ;
    wire new_AGEMA_signal_30256 ;
    wire new_AGEMA_signal_30257 ;
    wire new_AGEMA_signal_30258 ;
    wire new_AGEMA_signal_30259 ;
    wire new_AGEMA_signal_30260 ;
    wire new_AGEMA_signal_30261 ;
    wire new_AGEMA_signal_30262 ;
    wire new_AGEMA_signal_30263 ;
    wire new_AGEMA_signal_30264 ;
    wire new_AGEMA_signal_30265 ;
    wire new_AGEMA_signal_30266 ;
    wire new_AGEMA_signal_30267 ;
    wire new_AGEMA_signal_30268 ;
    wire new_AGEMA_signal_30269 ;
    wire new_AGEMA_signal_30270 ;
    wire new_AGEMA_signal_30271 ;
    wire new_AGEMA_signal_30272 ;
    wire new_AGEMA_signal_30273 ;
    wire new_AGEMA_signal_30274 ;
    wire new_AGEMA_signal_30275 ;
    wire new_AGEMA_signal_30276 ;
    wire new_AGEMA_signal_30277 ;
    wire new_AGEMA_signal_30278 ;
    wire new_AGEMA_signal_30279 ;
    wire new_AGEMA_signal_30280 ;
    wire new_AGEMA_signal_30281 ;
    wire new_AGEMA_signal_30282 ;
    wire new_AGEMA_signal_30283 ;
    wire new_AGEMA_signal_30284 ;
    wire new_AGEMA_signal_30285 ;
    wire new_AGEMA_signal_30286 ;
    wire new_AGEMA_signal_30287 ;
    wire new_AGEMA_signal_30288 ;
    wire new_AGEMA_signal_30289 ;
    wire new_AGEMA_signal_30290 ;
    wire new_AGEMA_signal_30291 ;
    wire new_AGEMA_signal_30292 ;
    wire new_AGEMA_signal_30293 ;
    wire new_AGEMA_signal_30294 ;
    wire new_AGEMA_signal_30295 ;
    wire new_AGEMA_signal_30296 ;
    wire new_AGEMA_signal_30297 ;
    wire new_AGEMA_signal_30298 ;
    wire new_AGEMA_signal_30299 ;
    wire new_AGEMA_signal_30300 ;
    wire new_AGEMA_signal_30301 ;
    wire new_AGEMA_signal_30302 ;
    wire new_AGEMA_signal_30303 ;
    wire new_AGEMA_signal_30304 ;
    wire new_AGEMA_signal_30305 ;
    wire new_AGEMA_signal_30306 ;
    wire new_AGEMA_signal_30307 ;
    wire new_AGEMA_signal_30308 ;
    wire new_AGEMA_signal_30309 ;
    wire new_AGEMA_signal_30310 ;
    wire new_AGEMA_signal_30311 ;
    wire new_AGEMA_signal_30312 ;
    wire new_AGEMA_signal_30313 ;
    wire new_AGEMA_signal_30314 ;
    wire new_AGEMA_signal_30315 ;
    wire new_AGEMA_signal_30316 ;
    wire new_AGEMA_signal_30317 ;
    wire new_AGEMA_signal_30318 ;
    wire new_AGEMA_signal_30319 ;
    wire new_AGEMA_signal_30320 ;
    wire new_AGEMA_signal_30321 ;
    wire new_AGEMA_signal_30322 ;
    wire new_AGEMA_signal_30323 ;
    wire new_AGEMA_signal_30324 ;
    wire new_AGEMA_signal_30325 ;
    wire new_AGEMA_signal_30326 ;
    wire new_AGEMA_signal_30327 ;
    wire new_AGEMA_signal_30328 ;
    wire new_AGEMA_signal_30329 ;
    wire new_AGEMA_signal_30330 ;
    wire new_AGEMA_signal_30331 ;
    wire new_AGEMA_signal_30332 ;
    wire new_AGEMA_signal_30333 ;
    wire new_AGEMA_signal_30334 ;
    wire new_AGEMA_signal_30335 ;
    wire new_AGEMA_signal_30336 ;
    wire new_AGEMA_signal_30337 ;
    wire new_AGEMA_signal_30338 ;
    wire new_AGEMA_signal_30339 ;
    wire new_AGEMA_signal_30340 ;
    wire new_AGEMA_signal_30341 ;
    wire new_AGEMA_signal_30342 ;
    wire new_AGEMA_signal_30343 ;
    wire new_AGEMA_signal_30344 ;
    wire new_AGEMA_signal_30345 ;
    wire new_AGEMA_signal_30346 ;
    wire new_AGEMA_signal_30347 ;
    wire new_AGEMA_signal_30348 ;
    wire new_AGEMA_signal_30349 ;
    wire new_AGEMA_signal_30350 ;
    wire new_AGEMA_signal_30351 ;
    wire new_AGEMA_signal_30352 ;
    wire new_AGEMA_signal_30353 ;
    wire new_AGEMA_signal_30354 ;
    wire new_AGEMA_signal_30355 ;
    wire new_AGEMA_signal_30356 ;
    wire new_AGEMA_signal_30357 ;
    wire new_AGEMA_signal_30358 ;
    wire new_AGEMA_signal_30359 ;
    wire new_AGEMA_signal_30360 ;
    wire new_AGEMA_signal_30361 ;
    wire new_AGEMA_signal_30362 ;
    wire new_AGEMA_signal_30363 ;
    wire new_AGEMA_signal_30364 ;
    wire new_AGEMA_signal_30365 ;
    wire new_AGEMA_signal_30366 ;
    wire new_AGEMA_signal_30367 ;
    wire new_AGEMA_signal_30368 ;
    wire new_AGEMA_signal_30369 ;
    wire new_AGEMA_signal_30370 ;
    wire new_AGEMA_signal_30371 ;
    wire new_AGEMA_signal_30372 ;
    wire new_AGEMA_signal_30373 ;
    wire new_AGEMA_signal_30374 ;
    wire new_AGEMA_signal_30375 ;
    wire new_AGEMA_signal_30376 ;
    wire new_AGEMA_signal_30377 ;
    wire new_AGEMA_signal_30378 ;
    wire new_AGEMA_signal_30379 ;
    wire new_AGEMA_signal_30380 ;
    wire new_AGEMA_signal_30381 ;
    wire new_AGEMA_signal_30382 ;
    wire new_AGEMA_signal_30383 ;
    wire new_AGEMA_signal_30384 ;
    wire new_AGEMA_signal_30385 ;
    wire new_AGEMA_signal_30386 ;
    wire new_AGEMA_signal_30387 ;
    wire new_AGEMA_signal_30388 ;
    wire new_AGEMA_signal_30389 ;
    wire new_AGEMA_signal_30390 ;
    wire new_AGEMA_signal_30391 ;
    wire new_AGEMA_signal_30392 ;
    wire new_AGEMA_signal_30393 ;
    wire new_AGEMA_signal_30394 ;
    wire new_AGEMA_signal_30395 ;
    wire new_AGEMA_signal_30396 ;
    wire new_AGEMA_signal_30397 ;
    wire new_AGEMA_signal_30398 ;
    wire new_AGEMA_signal_30399 ;
    wire new_AGEMA_signal_30400 ;
    wire new_AGEMA_signal_30401 ;
    wire new_AGEMA_signal_30402 ;
    wire new_AGEMA_signal_30403 ;
    wire new_AGEMA_signal_30404 ;
    wire new_AGEMA_signal_30405 ;
    wire new_AGEMA_signal_30406 ;
    wire new_AGEMA_signal_30407 ;
    wire new_AGEMA_signal_30408 ;
    wire new_AGEMA_signal_30409 ;
    wire new_AGEMA_signal_30410 ;
    wire new_AGEMA_signal_30411 ;
    wire new_AGEMA_signal_30412 ;
    wire new_AGEMA_signal_30413 ;
    wire new_AGEMA_signal_30414 ;
    wire new_AGEMA_signal_30415 ;
    wire new_AGEMA_signal_30416 ;
    wire new_AGEMA_signal_30417 ;
    wire new_AGEMA_signal_30418 ;
    wire new_AGEMA_signal_30419 ;
    wire new_AGEMA_signal_30420 ;
    wire new_AGEMA_signal_30421 ;
    wire new_AGEMA_signal_30422 ;
    wire new_AGEMA_signal_30423 ;
    wire new_AGEMA_signal_30424 ;
    wire new_AGEMA_signal_30425 ;
    wire new_AGEMA_signal_30426 ;
    wire new_AGEMA_signal_30427 ;
    wire new_AGEMA_signal_30428 ;
    wire new_AGEMA_signal_30429 ;
    wire new_AGEMA_signal_30430 ;
    wire new_AGEMA_signal_30431 ;
    wire new_AGEMA_signal_30432 ;
    wire new_AGEMA_signal_30433 ;
    wire new_AGEMA_signal_30434 ;
    wire new_AGEMA_signal_30435 ;
    wire new_AGEMA_signal_30436 ;
    wire new_AGEMA_signal_30437 ;
    wire new_AGEMA_signal_30438 ;
    wire new_AGEMA_signal_30439 ;
    wire new_AGEMA_signal_30440 ;
    wire new_AGEMA_signal_30441 ;
    wire new_AGEMA_signal_30442 ;
    wire new_AGEMA_signal_30443 ;
    wire new_AGEMA_signal_30444 ;
    wire new_AGEMA_signal_30445 ;
    wire new_AGEMA_signal_30446 ;
    wire new_AGEMA_signal_30447 ;
    wire new_AGEMA_signal_30448 ;
    wire new_AGEMA_signal_30449 ;
    wire new_AGEMA_signal_30450 ;
    wire new_AGEMA_signal_30451 ;
    wire new_AGEMA_signal_30452 ;
    wire new_AGEMA_signal_30453 ;
    wire new_AGEMA_signal_30454 ;
    wire new_AGEMA_signal_30455 ;
    wire new_AGEMA_signal_30456 ;
    wire new_AGEMA_signal_30457 ;
    wire new_AGEMA_signal_30458 ;
    wire new_AGEMA_signal_30459 ;
    wire new_AGEMA_signal_30460 ;
    wire new_AGEMA_signal_30461 ;
    wire new_AGEMA_signal_30462 ;
    wire new_AGEMA_signal_30463 ;
    wire new_AGEMA_signal_30464 ;
    wire new_AGEMA_signal_30465 ;
    wire new_AGEMA_signal_30466 ;
    wire new_AGEMA_signal_30467 ;
    wire new_AGEMA_signal_30468 ;
    wire new_AGEMA_signal_30469 ;
    wire new_AGEMA_signal_30470 ;
    wire new_AGEMA_signal_30471 ;
    wire new_AGEMA_signal_30472 ;
    wire new_AGEMA_signal_30473 ;
    wire new_AGEMA_signal_30474 ;
    wire new_AGEMA_signal_30475 ;
    wire new_AGEMA_signal_30476 ;
    wire new_AGEMA_signal_30477 ;
    wire new_AGEMA_signal_30478 ;
    wire new_AGEMA_signal_30479 ;
    wire new_AGEMA_signal_30480 ;
    wire new_AGEMA_signal_30481 ;
    wire new_AGEMA_signal_30482 ;
    wire new_AGEMA_signal_30483 ;
    wire new_AGEMA_signal_30484 ;
    wire new_AGEMA_signal_30485 ;
    wire new_AGEMA_signal_30486 ;
    wire new_AGEMA_signal_30487 ;
    wire new_AGEMA_signal_30488 ;
    wire new_AGEMA_signal_30489 ;
    wire new_AGEMA_signal_30490 ;
    wire new_AGEMA_signal_30491 ;
    wire new_AGEMA_signal_30492 ;
    wire new_AGEMA_signal_30493 ;
    wire new_AGEMA_signal_30494 ;
    wire new_AGEMA_signal_30495 ;
    wire new_AGEMA_signal_30496 ;
    wire new_AGEMA_signal_30497 ;
    wire new_AGEMA_signal_30498 ;
    wire new_AGEMA_signal_30499 ;
    wire new_AGEMA_signal_30500 ;
    wire new_AGEMA_signal_30501 ;
    wire new_AGEMA_signal_30502 ;
    wire new_AGEMA_signal_30503 ;
    wire new_AGEMA_signal_30504 ;
    wire new_AGEMA_signal_30505 ;
    wire new_AGEMA_signal_30506 ;
    wire new_AGEMA_signal_30507 ;
    wire new_AGEMA_signal_30508 ;
    wire new_AGEMA_signal_30509 ;
    wire new_AGEMA_signal_30510 ;
    wire new_AGEMA_signal_30511 ;
    wire new_AGEMA_signal_30512 ;
    wire new_AGEMA_signal_30513 ;
    wire new_AGEMA_signal_30514 ;
    wire new_AGEMA_signal_30515 ;
    wire new_AGEMA_signal_30516 ;
    wire new_AGEMA_signal_30517 ;
    wire new_AGEMA_signal_30518 ;
    wire new_AGEMA_signal_30519 ;
    wire new_AGEMA_signal_30520 ;
    wire new_AGEMA_signal_30521 ;
    wire new_AGEMA_signal_30522 ;
    wire new_AGEMA_signal_30523 ;
    wire new_AGEMA_signal_30524 ;
    wire new_AGEMA_signal_30525 ;
    wire new_AGEMA_signal_30526 ;
    wire new_AGEMA_signal_30527 ;
    wire new_AGEMA_signal_30528 ;
    wire new_AGEMA_signal_30529 ;
    wire new_AGEMA_signal_30530 ;
    wire new_AGEMA_signal_30531 ;
    wire new_AGEMA_signal_30532 ;
    wire new_AGEMA_signal_30533 ;
    wire new_AGEMA_signal_30534 ;
    wire new_AGEMA_signal_30535 ;
    wire new_AGEMA_signal_30536 ;
    wire new_AGEMA_signal_30537 ;
    wire new_AGEMA_signal_30538 ;
    wire new_AGEMA_signal_30539 ;
    wire new_AGEMA_signal_30540 ;
    wire new_AGEMA_signal_30541 ;
    wire new_AGEMA_signal_30542 ;
    wire new_AGEMA_signal_30543 ;
    wire new_AGEMA_signal_30544 ;
    wire new_AGEMA_signal_30545 ;
    wire new_AGEMA_signal_30546 ;
    wire new_AGEMA_signal_30547 ;
    wire new_AGEMA_signal_30548 ;
    wire new_AGEMA_signal_30549 ;
    wire new_AGEMA_signal_30550 ;
    wire new_AGEMA_signal_30551 ;
    wire new_AGEMA_signal_30552 ;
    wire new_AGEMA_signal_30553 ;
    wire new_AGEMA_signal_30554 ;
    wire new_AGEMA_signal_30555 ;
    wire new_AGEMA_signal_30556 ;
    wire new_AGEMA_signal_30557 ;
    wire new_AGEMA_signal_30558 ;
    wire new_AGEMA_signal_30559 ;
    wire new_AGEMA_signal_30560 ;
    wire new_AGEMA_signal_30561 ;
    wire new_AGEMA_signal_30562 ;
    wire new_AGEMA_signal_30563 ;
    wire new_AGEMA_signal_30564 ;
    wire new_AGEMA_signal_30565 ;
    wire new_AGEMA_signal_30566 ;
    wire new_AGEMA_signal_30567 ;
    wire new_AGEMA_signal_30568 ;
    wire new_AGEMA_signal_30569 ;
    wire new_AGEMA_signal_30570 ;
    wire new_AGEMA_signal_30571 ;
    wire new_AGEMA_signal_30572 ;
    wire new_AGEMA_signal_30573 ;
    wire new_AGEMA_signal_30574 ;
    wire new_AGEMA_signal_30575 ;
    wire new_AGEMA_signal_30576 ;
    wire new_AGEMA_signal_30577 ;
    wire new_AGEMA_signal_30578 ;
    wire new_AGEMA_signal_30579 ;
    wire new_AGEMA_signal_30580 ;
    wire new_AGEMA_signal_30581 ;
    wire new_AGEMA_signal_30582 ;
    wire new_AGEMA_signal_30583 ;
    wire new_AGEMA_signal_30584 ;
    wire new_AGEMA_signal_30585 ;
    wire new_AGEMA_signal_30586 ;
    wire new_AGEMA_signal_30587 ;
    wire new_AGEMA_signal_30588 ;
    wire new_AGEMA_signal_30589 ;
    wire new_AGEMA_signal_30590 ;
    wire new_AGEMA_signal_30591 ;
    wire new_AGEMA_signal_30592 ;
    wire new_AGEMA_signal_30593 ;
    wire new_AGEMA_signal_30594 ;
    wire new_AGEMA_signal_30595 ;
    wire new_AGEMA_signal_30596 ;
    wire new_AGEMA_signal_30597 ;
    wire new_AGEMA_signal_30598 ;
    wire new_AGEMA_signal_30599 ;
    wire new_AGEMA_signal_30600 ;
    wire new_AGEMA_signal_30601 ;
    wire new_AGEMA_signal_30602 ;
    wire new_AGEMA_signal_30603 ;
    wire new_AGEMA_signal_30604 ;
    wire new_AGEMA_signal_30605 ;
    wire new_AGEMA_signal_30606 ;
    wire new_AGEMA_signal_30607 ;
    wire new_AGEMA_signal_30608 ;
    wire new_AGEMA_signal_30609 ;
    wire new_AGEMA_signal_30610 ;
    wire new_AGEMA_signal_30611 ;
    wire new_AGEMA_signal_30612 ;
    wire new_AGEMA_signal_30613 ;
    wire new_AGEMA_signal_30614 ;
    wire new_AGEMA_signal_30615 ;
    wire new_AGEMA_signal_30616 ;
    wire new_AGEMA_signal_30617 ;
    wire new_AGEMA_signal_30618 ;
    wire new_AGEMA_signal_30619 ;
    wire new_AGEMA_signal_30620 ;
    wire new_AGEMA_signal_30621 ;
    wire new_AGEMA_signal_30622 ;
    wire new_AGEMA_signal_30623 ;
    wire new_AGEMA_signal_30624 ;
    wire new_AGEMA_signal_30625 ;
    wire new_AGEMA_signal_30626 ;
    wire new_AGEMA_signal_30627 ;
    wire new_AGEMA_signal_30628 ;
    wire new_AGEMA_signal_30629 ;
    wire new_AGEMA_signal_30630 ;
    wire new_AGEMA_signal_30631 ;
    wire new_AGEMA_signal_30632 ;
    wire new_AGEMA_signal_30633 ;
    wire new_AGEMA_signal_30634 ;
    wire new_AGEMA_signal_30635 ;
    wire new_AGEMA_signal_30636 ;
    wire new_AGEMA_signal_30637 ;
    wire new_AGEMA_signal_30638 ;
    wire new_AGEMA_signal_30639 ;
    wire new_AGEMA_signal_30640 ;
    wire new_AGEMA_signal_30641 ;
    wire new_AGEMA_signal_30642 ;
    wire new_AGEMA_signal_30643 ;
    wire new_AGEMA_signal_30644 ;
    wire new_AGEMA_signal_30645 ;
    wire new_AGEMA_signal_30646 ;
    wire new_AGEMA_signal_30647 ;
    wire new_AGEMA_signal_30648 ;
    wire new_AGEMA_signal_30649 ;
    wire new_AGEMA_signal_30650 ;
    wire new_AGEMA_signal_30651 ;
    wire new_AGEMA_signal_30652 ;
    wire new_AGEMA_signal_30653 ;
    wire new_AGEMA_signal_30654 ;
    wire new_AGEMA_signal_30655 ;
    wire new_AGEMA_signal_30656 ;
    wire new_AGEMA_signal_30657 ;
    wire new_AGEMA_signal_30658 ;
    wire new_AGEMA_signal_30659 ;
    wire new_AGEMA_signal_30660 ;
    wire new_AGEMA_signal_30661 ;
    wire new_AGEMA_signal_30662 ;
    wire new_AGEMA_signal_30663 ;
    wire new_AGEMA_signal_30664 ;
    wire new_AGEMA_signal_30665 ;
    wire new_AGEMA_signal_30666 ;
    wire new_AGEMA_signal_30667 ;
    wire new_AGEMA_signal_30668 ;
    wire new_AGEMA_signal_30669 ;
    wire new_AGEMA_signal_30670 ;
    wire new_AGEMA_signal_30671 ;
    wire new_AGEMA_signal_30672 ;
    wire new_AGEMA_signal_30673 ;
    wire new_AGEMA_signal_30674 ;
    wire new_AGEMA_signal_30675 ;
    wire new_AGEMA_signal_30676 ;
    wire new_AGEMA_signal_30677 ;
    wire new_AGEMA_signal_30678 ;
    wire new_AGEMA_signal_30679 ;
    wire new_AGEMA_signal_30680 ;
    wire new_AGEMA_signal_30681 ;
    wire new_AGEMA_signal_30682 ;
    wire new_AGEMA_signal_30683 ;
    wire new_AGEMA_signal_30684 ;
    wire new_AGEMA_signal_30685 ;
    wire new_AGEMA_signal_30686 ;
    wire new_AGEMA_signal_30687 ;
    wire new_AGEMA_signal_30688 ;
    wire new_AGEMA_signal_30689 ;
    wire new_AGEMA_signal_30690 ;
    wire new_AGEMA_signal_30691 ;
    wire new_AGEMA_signal_30692 ;
    wire new_AGEMA_signal_30693 ;
    wire new_AGEMA_signal_30694 ;
    wire new_AGEMA_signal_30695 ;
    wire new_AGEMA_signal_30696 ;
    wire new_AGEMA_signal_30697 ;
    wire new_AGEMA_signal_30698 ;
    wire new_AGEMA_signal_30699 ;
    wire new_AGEMA_signal_30700 ;
    wire new_AGEMA_signal_30701 ;
    wire new_AGEMA_signal_30702 ;
    wire new_AGEMA_signal_30703 ;
    wire new_AGEMA_signal_30704 ;
    wire new_AGEMA_signal_30705 ;
    wire new_AGEMA_signal_30706 ;
    wire new_AGEMA_signal_30707 ;
    wire new_AGEMA_signal_30708 ;
    wire new_AGEMA_signal_30709 ;
    wire new_AGEMA_signal_30710 ;
    wire new_AGEMA_signal_30711 ;
    wire new_AGEMA_signal_30712 ;
    wire new_AGEMA_signal_30713 ;
    wire new_AGEMA_signal_30714 ;
    wire new_AGEMA_signal_30715 ;
    wire new_AGEMA_signal_30716 ;
    wire new_AGEMA_signal_30717 ;
    wire new_AGEMA_signal_30718 ;
    wire new_AGEMA_signal_30719 ;
    wire new_AGEMA_signal_30720 ;
    wire new_AGEMA_signal_30721 ;
    wire new_AGEMA_signal_30722 ;
    wire new_AGEMA_signal_30723 ;
    wire new_AGEMA_signal_30724 ;
    wire new_AGEMA_signal_30725 ;
    wire new_AGEMA_signal_30726 ;
    wire new_AGEMA_signal_30727 ;
    wire new_AGEMA_signal_30728 ;
    wire new_AGEMA_signal_30729 ;
    wire new_AGEMA_signal_30730 ;
    wire new_AGEMA_signal_30731 ;
    wire new_AGEMA_signal_30732 ;
    wire new_AGEMA_signal_30733 ;
    wire new_AGEMA_signal_30734 ;
    wire new_AGEMA_signal_30735 ;
    wire new_AGEMA_signal_30736 ;
    wire new_AGEMA_signal_30737 ;
    wire new_AGEMA_signal_30738 ;
    wire new_AGEMA_signal_30739 ;
    wire new_AGEMA_signal_30740 ;
    wire new_AGEMA_signal_30741 ;
    wire new_AGEMA_signal_30742 ;
    wire new_AGEMA_signal_30743 ;
    wire new_AGEMA_signal_30744 ;
    wire new_AGEMA_signal_30745 ;
    wire new_AGEMA_signal_30746 ;
    wire new_AGEMA_signal_30747 ;
    wire new_AGEMA_signal_30748 ;
    wire new_AGEMA_signal_30749 ;
    wire new_AGEMA_signal_30750 ;
    wire new_AGEMA_signal_30751 ;
    wire new_AGEMA_signal_30752 ;
    wire new_AGEMA_signal_30753 ;
    wire new_AGEMA_signal_30754 ;
    wire new_AGEMA_signal_30755 ;
    wire new_AGEMA_signal_30756 ;
    wire new_AGEMA_signal_30757 ;
    wire new_AGEMA_signal_30758 ;
    wire new_AGEMA_signal_30759 ;
    wire new_AGEMA_signal_30760 ;
    wire new_AGEMA_signal_30761 ;
    wire new_AGEMA_signal_30762 ;
    wire new_AGEMA_signal_30763 ;
    wire new_AGEMA_signal_30764 ;
    wire new_AGEMA_signal_30765 ;
    wire new_AGEMA_signal_30766 ;
    wire new_AGEMA_signal_30767 ;
    wire new_AGEMA_signal_30768 ;
    wire new_AGEMA_signal_30769 ;
    wire new_AGEMA_signal_30770 ;
    wire new_AGEMA_signal_30771 ;
    wire new_AGEMA_signal_30772 ;
    wire new_AGEMA_signal_30773 ;
    wire new_AGEMA_signal_30774 ;
    wire new_AGEMA_signal_30775 ;
    wire new_AGEMA_signal_30776 ;
    wire new_AGEMA_signal_30777 ;
    wire new_AGEMA_signal_30778 ;
    wire new_AGEMA_signal_30779 ;
    wire new_AGEMA_signal_30780 ;
    wire new_AGEMA_signal_30781 ;
    wire new_AGEMA_signal_30782 ;
    wire new_AGEMA_signal_30783 ;
    wire new_AGEMA_signal_30784 ;
    wire new_AGEMA_signal_30785 ;
    wire new_AGEMA_signal_30786 ;
    wire new_AGEMA_signal_30787 ;
    wire new_AGEMA_signal_30788 ;
    wire new_AGEMA_signal_30789 ;
    wire new_AGEMA_signal_30790 ;
    wire new_AGEMA_signal_30791 ;
    wire new_AGEMA_signal_30792 ;
    wire new_AGEMA_signal_30793 ;
    wire new_AGEMA_signal_30794 ;
    wire new_AGEMA_signal_30795 ;
    wire new_AGEMA_signal_30796 ;
    wire new_AGEMA_signal_30797 ;
    wire new_AGEMA_signal_30798 ;
    wire new_AGEMA_signal_30799 ;
    wire new_AGEMA_signal_30800 ;
    wire new_AGEMA_signal_30801 ;
    wire new_AGEMA_signal_30802 ;
    wire new_AGEMA_signal_30803 ;
    wire new_AGEMA_signal_30804 ;
    wire new_AGEMA_signal_30805 ;
    wire new_AGEMA_signal_30806 ;
    wire new_AGEMA_signal_30807 ;
    wire new_AGEMA_signal_30808 ;
    wire new_AGEMA_signal_30809 ;
    wire new_AGEMA_signal_30810 ;
    wire new_AGEMA_signal_30811 ;
    wire new_AGEMA_signal_30812 ;
    wire new_AGEMA_signal_30813 ;
    wire new_AGEMA_signal_30814 ;
    wire new_AGEMA_signal_30815 ;
    wire new_AGEMA_signal_30816 ;
    wire new_AGEMA_signal_30817 ;
    wire new_AGEMA_signal_30818 ;
    wire new_AGEMA_signal_30819 ;
    wire new_AGEMA_signal_30820 ;
    wire new_AGEMA_signal_30821 ;
    wire new_AGEMA_signal_30822 ;
    wire new_AGEMA_signal_30823 ;
    wire new_AGEMA_signal_30824 ;
    wire new_AGEMA_signal_30825 ;
    wire new_AGEMA_signal_30826 ;
    wire new_AGEMA_signal_30827 ;
    wire new_AGEMA_signal_30828 ;
    wire new_AGEMA_signal_30829 ;
    wire new_AGEMA_signal_30830 ;
    wire new_AGEMA_signal_30831 ;
    wire new_AGEMA_signal_30832 ;
    wire new_AGEMA_signal_30833 ;
    wire new_AGEMA_signal_30834 ;
    wire new_AGEMA_signal_30835 ;
    wire new_AGEMA_signal_30836 ;
    wire new_AGEMA_signal_30837 ;
    wire new_AGEMA_signal_30838 ;
    wire new_AGEMA_signal_30839 ;
    wire new_AGEMA_signal_30840 ;
    wire new_AGEMA_signal_30841 ;
    wire new_AGEMA_signal_30842 ;
    wire new_AGEMA_signal_30843 ;
    wire new_AGEMA_signal_30844 ;
    wire new_AGEMA_signal_30845 ;
    wire new_AGEMA_signal_30846 ;
    wire new_AGEMA_signal_30847 ;
    wire new_AGEMA_signal_30848 ;
    wire new_AGEMA_signal_30849 ;
    wire new_AGEMA_signal_30850 ;
    wire new_AGEMA_signal_30851 ;
    wire new_AGEMA_signal_30852 ;
    wire new_AGEMA_signal_30853 ;
    wire new_AGEMA_signal_30854 ;
    wire new_AGEMA_signal_30855 ;
    wire new_AGEMA_signal_30856 ;
    wire new_AGEMA_signal_30857 ;
    wire new_AGEMA_signal_30858 ;
    wire new_AGEMA_signal_30859 ;
    wire new_AGEMA_signal_30860 ;
    wire new_AGEMA_signal_30861 ;
    wire new_AGEMA_signal_30862 ;
    wire new_AGEMA_signal_30863 ;
    wire new_AGEMA_signal_30864 ;
    wire new_AGEMA_signal_30865 ;
    wire new_AGEMA_signal_30866 ;
    wire new_AGEMA_signal_30867 ;
    wire new_AGEMA_signal_30868 ;
    wire new_AGEMA_signal_30869 ;
    wire new_AGEMA_signal_30870 ;
    wire new_AGEMA_signal_30871 ;
    wire new_AGEMA_signal_30872 ;
    wire new_AGEMA_signal_30873 ;
    wire new_AGEMA_signal_30874 ;
    wire new_AGEMA_signal_30875 ;
    wire new_AGEMA_signal_30876 ;
    wire new_AGEMA_signal_30877 ;
    wire new_AGEMA_signal_30878 ;
    wire new_AGEMA_signal_30879 ;
    wire new_AGEMA_signal_30880 ;
    wire new_AGEMA_signal_30881 ;
    wire new_AGEMA_signal_30882 ;
    wire new_AGEMA_signal_30883 ;
    wire new_AGEMA_signal_30884 ;
    wire new_AGEMA_signal_30885 ;
    wire new_AGEMA_signal_30886 ;
    wire new_AGEMA_signal_30887 ;
    wire new_AGEMA_signal_30888 ;
    wire new_AGEMA_signal_30889 ;
    wire new_AGEMA_signal_30890 ;
    wire new_AGEMA_signal_30891 ;
    wire new_AGEMA_signal_30892 ;
    wire new_AGEMA_signal_30893 ;
    wire new_AGEMA_signal_30894 ;
    wire new_AGEMA_signal_30895 ;
    wire new_AGEMA_signal_30896 ;
    wire new_AGEMA_signal_30897 ;
    wire new_AGEMA_signal_30898 ;
    wire new_AGEMA_signal_30899 ;
    wire new_AGEMA_signal_30900 ;
    wire new_AGEMA_signal_30901 ;
    wire new_AGEMA_signal_30902 ;
    wire new_AGEMA_signal_30903 ;
    wire new_AGEMA_signal_30904 ;
    wire new_AGEMA_signal_30905 ;
    wire new_AGEMA_signal_30906 ;
    wire new_AGEMA_signal_30907 ;
    wire new_AGEMA_signal_30908 ;
    wire new_AGEMA_signal_30909 ;
    wire new_AGEMA_signal_30910 ;
    wire new_AGEMA_signal_30911 ;
    wire new_AGEMA_signal_30912 ;
    wire new_AGEMA_signal_30913 ;
    wire new_AGEMA_signal_30914 ;
    wire new_AGEMA_signal_30915 ;
    wire new_AGEMA_signal_30916 ;
    wire new_AGEMA_signal_30917 ;
    wire new_AGEMA_signal_30918 ;
    wire new_AGEMA_signal_30919 ;
    wire new_AGEMA_signal_30920 ;
    wire new_AGEMA_signal_30921 ;
    wire new_AGEMA_signal_30922 ;
    wire new_AGEMA_signal_30923 ;
    wire new_AGEMA_signal_30924 ;
    wire new_AGEMA_signal_30925 ;
    wire new_AGEMA_signal_30926 ;
    wire new_AGEMA_signal_30927 ;
    wire new_AGEMA_signal_30928 ;
    wire new_AGEMA_signal_30929 ;
    wire new_AGEMA_signal_30930 ;
    wire new_AGEMA_signal_30931 ;
    wire new_AGEMA_signal_30932 ;
    wire new_AGEMA_signal_30933 ;
    wire new_AGEMA_signal_30934 ;
    wire new_AGEMA_signal_30935 ;
    wire new_AGEMA_signal_30936 ;
    wire new_AGEMA_signal_30937 ;
    wire new_AGEMA_signal_30938 ;
    wire new_AGEMA_signal_30939 ;
    wire new_AGEMA_signal_30940 ;
    wire new_AGEMA_signal_30941 ;
    wire new_AGEMA_signal_30942 ;
    wire new_AGEMA_signal_30943 ;
    wire new_AGEMA_signal_30944 ;
    wire new_AGEMA_signal_30945 ;
    wire new_AGEMA_signal_30946 ;
    wire new_AGEMA_signal_30947 ;
    wire new_AGEMA_signal_30948 ;
    wire new_AGEMA_signal_30949 ;
    wire new_AGEMA_signal_30950 ;
    wire new_AGEMA_signal_30951 ;
    wire new_AGEMA_signal_30952 ;
    wire new_AGEMA_signal_30953 ;
    wire new_AGEMA_signal_30954 ;
    wire new_AGEMA_signal_30955 ;
    wire new_AGEMA_signal_30956 ;
    wire new_AGEMA_signal_30957 ;
    wire new_AGEMA_signal_30958 ;
    wire new_AGEMA_signal_30959 ;
    wire new_AGEMA_signal_30960 ;
    wire new_AGEMA_signal_30961 ;
    wire new_AGEMA_signal_30962 ;
    wire new_AGEMA_signal_30963 ;
    wire new_AGEMA_signal_30964 ;
    wire new_AGEMA_signal_30965 ;
    wire new_AGEMA_signal_30966 ;
    wire new_AGEMA_signal_30967 ;
    wire new_AGEMA_signal_30968 ;
    wire new_AGEMA_signal_30969 ;
    wire new_AGEMA_signal_30970 ;
    wire new_AGEMA_signal_30971 ;
    wire new_AGEMA_signal_30972 ;
    wire new_AGEMA_signal_30973 ;
    wire new_AGEMA_signal_30974 ;
    wire new_AGEMA_signal_30975 ;
    wire new_AGEMA_signal_30976 ;
    wire new_AGEMA_signal_30977 ;
    wire new_AGEMA_signal_30978 ;
    wire new_AGEMA_signal_30979 ;
    wire new_AGEMA_signal_30980 ;
    wire new_AGEMA_signal_30981 ;
    wire new_AGEMA_signal_30982 ;
    wire new_AGEMA_signal_30983 ;
    wire new_AGEMA_signal_30984 ;
    wire new_AGEMA_signal_30985 ;
    wire new_AGEMA_signal_30986 ;
    wire new_AGEMA_signal_30987 ;
    wire new_AGEMA_signal_30988 ;
    wire new_AGEMA_signal_30989 ;
    wire new_AGEMA_signal_30990 ;
    wire new_AGEMA_signal_30991 ;
    wire new_AGEMA_signal_30992 ;
    wire new_AGEMA_signal_30993 ;
    wire new_AGEMA_signal_30994 ;
    wire new_AGEMA_signal_30995 ;
    wire new_AGEMA_signal_30996 ;
    wire new_AGEMA_signal_30997 ;
    wire new_AGEMA_signal_30998 ;
    wire new_AGEMA_signal_30999 ;
    wire new_AGEMA_signal_31000 ;
    wire new_AGEMA_signal_31001 ;
    wire new_AGEMA_signal_31002 ;
    wire new_AGEMA_signal_31003 ;
    wire new_AGEMA_signal_31004 ;
    wire new_AGEMA_signal_31005 ;
    wire new_AGEMA_signal_31006 ;
    wire new_AGEMA_signal_31007 ;
    wire new_AGEMA_signal_31008 ;
    wire new_AGEMA_signal_31009 ;
    wire new_AGEMA_signal_31010 ;
    wire new_AGEMA_signal_31011 ;
    wire new_AGEMA_signal_31012 ;
    wire new_AGEMA_signal_31013 ;
    wire new_AGEMA_signal_31014 ;
    wire new_AGEMA_signal_31015 ;
    wire new_AGEMA_signal_31016 ;
    wire new_AGEMA_signal_31017 ;
    wire new_AGEMA_signal_31018 ;
    wire new_AGEMA_signal_31019 ;
    wire new_AGEMA_signal_31020 ;
    wire new_AGEMA_signal_31021 ;
    wire new_AGEMA_signal_31022 ;
    wire new_AGEMA_signal_31023 ;
    wire new_AGEMA_signal_31024 ;
    wire new_AGEMA_signal_31025 ;
    wire new_AGEMA_signal_31026 ;
    wire new_AGEMA_signal_31027 ;
    wire new_AGEMA_signal_31028 ;
    wire new_AGEMA_signal_31029 ;
    wire new_AGEMA_signal_31030 ;
    wire new_AGEMA_signal_31031 ;
    wire new_AGEMA_signal_31032 ;
    wire new_AGEMA_signal_31033 ;
    wire new_AGEMA_signal_31034 ;
    wire new_AGEMA_signal_31035 ;
    wire new_AGEMA_signal_31036 ;
    wire new_AGEMA_signal_31037 ;
    wire new_AGEMA_signal_31038 ;
    wire new_AGEMA_signal_31039 ;
    wire new_AGEMA_signal_31040 ;
    wire new_AGEMA_signal_31041 ;
    wire new_AGEMA_signal_31042 ;
    wire new_AGEMA_signal_31043 ;
    wire new_AGEMA_signal_31044 ;
    wire new_AGEMA_signal_31045 ;
    wire new_AGEMA_signal_31046 ;
    wire new_AGEMA_signal_31047 ;
    wire new_AGEMA_signal_31048 ;
    wire new_AGEMA_signal_31049 ;
    wire new_AGEMA_signal_31050 ;
    wire new_AGEMA_signal_31051 ;
    wire new_AGEMA_signal_31052 ;
    wire new_AGEMA_signal_31053 ;
    wire new_AGEMA_signal_31054 ;
    wire new_AGEMA_signal_31055 ;
    wire new_AGEMA_signal_31056 ;
    wire new_AGEMA_signal_31057 ;
    wire new_AGEMA_signal_31058 ;
    wire new_AGEMA_signal_31059 ;
    wire new_AGEMA_signal_31060 ;
    wire new_AGEMA_signal_31061 ;
    wire new_AGEMA_signal_31062 ;
    wire new_AGEMA_signal_31063 ;
    wire new_AGEMA_signal_31064 ;
    wire new_AGEMA_signal_31065 ;
    wire new_AGEMA_signal_31066 ;
    wire new_AGEMA_signal_31067 ;
    wire new_AGEMA_signal_31068 ;
    wire new_AGEMA_signal_31069 ;
    wire new_AGEMA_signal_31070 ;
    wire new_AGEMA_signal_31071 ;
    wire new_AGEMA_signal_31072 ;
    wire new_AGEMA_signal_31073 ;
    wire new_AGEMA_signal_31074 ;
    wire new_AGEMA_signal_31075 ;
    wire new_AGEMA_signal_31076 ;
    wire new_AGEMA_signal_31077 ;
    wire new_AGEMA_signal_31078 ;
    wire new_AGEMA_signal_31079 ;
    wire new_AGEMA_signal_31080 ;
    wire new_AGEMA_signal_31081 ;
    wire new_AGEMA_signal_31082 ;
    wire new_AGEMA_signal_31083 ;
    wire new_AGEMA_signal_31084 ;
    wire new_AGEMA_signal_31085 ;
    wire new_AGEMA_signal_31086 ;
    wire new_AGEMA_signal_31087 ;
    wire new_AGEMA_signal_31088 ;
    wire new_AGEMA_signal_31089 ;
    wire new_AGEMA_signal_31090 ;
    wire new_AGEMA_signal_31091 ;
    wire new_AGEMA_signal_31092 ;
    wire new_AGEMA_signal_31093 ;
    wire new_AGEMA_signal_31094 ;
    wire new_AGEMA_signal_31095 ;
    wire new_AGEMA_signal_31096 ;
    wire new_AGEMA_signal_31097 ;
    wire new_AGEMA_signal_31098 ;
    wire new_AGEMA_signal_31099 ;
    wire new_AGEMA_signal_31100 ;
    wire new_AGEMA_signal_31101 ;
    wire new_AGEMA_signal_31102 ;
    wire new_AGEMA_signal_31103 ;
    wire new_AGEMA_signal_31104 ;
    wire new_AGEMA_signal_31105 ;
    wire new_AGEMA_signal_31106 ;
    wire new_AGEMA_signal_31107 ;
    wire new_AGEMA_signal_31108 ;
    wire new_AGEMA_signal_31109 ;
    wire new_AGEMA_signal_31110 ;
    wire new_AGEMA_signal_31111 ;
    wire new_AGEMA_signal_31112 ;
    wire new_AGEMA_signal_31113 ;
    wire new_AGEMA_signal_31114 ;
    wire new_AGEMA_signal_31115 ;
    wire new_AGEMA_signal_31116 ;
    wire new_AGEMA_signal_31117 ;
    wire new_AGEMA_signal_31118 ;
    wire new_AGEMA_signal_31119 ;
    wire new_AGEMA_signal_31120 ;
    wire new_AGEMA_signal_31121 ;
    wire new_AGEMA_signal_31122 ;
    wire new_AGEMA_signal_31123 ;
    wire new_AGEMA_signal_31124 ;
    wire new_AGEMA_signal_31125 ;
    wire new_AGEMA_signal_31126 ;
    wire new_AGEMA_signal_31127 ;
    wire new_AGEMA_signal_31128 ;
    wire new_AGEMA_signal_31129 ;
    wire new_AGEMA_signal_31130 ;
    wire new_AGEMA_signal_31131 ;
    wire new_AGEMA_signal_31132 ;
    wire new_AGEMA_signal_31133 ;
    wire new_AGEMA_signal_31134 ;
    wire new_AGEMA_signal_31135 ;
    wire new_AGEMA_signal_31136 ;
    wire new_AGEMA_signal_31137 ;
    wire new_AGEMA_signal_31138 ;
    wire new_AGEMA_signal_31139 ;
    wire new_AGEMA_signal_31140 ;
    wire new_AGEMA_signal_31141 ;
    wire new_AGEMA_signal_31142 ;
    wire new_AGEMA_signal_31143 ;
    wire new_AGEMA_signal_31144 ;
    wire new_AGEMA_signal_31145 ;
    wire new_AGEMA_signal_31146 ;
    wire new_AGEMA_signal_31147 ;
    wire new_AGEMA_signal_31148 ;
    wire new_AGEMA_signal_31149 ;
    wire new_AGEMA_signal_31150 ;
    wire new_AGEMA_signal_31151 ;
    wire new_AGEMA_signal_31152 ;
    wire new_AGEMA_signal_31153 ;
    wire new_AGEMA_signal_31154 ;
    wire new_AGEMA_signal_31155 ;
    wire new_AGEMA_signal_31156 ;
    wire new_AGEMA_signal_31157 ;
    wire new_AGEMA_signal_31158 ;
    wire new_AGEMA_signal_31159 ;
    wire new_AGEMA_signal_31160 ;
    wire new_AGEMA_signal_31161 ;
    wire new_AGEMA_signal_31162 ;
    wire new_AGEMA_signal_31163 ;
    wire new_AGEMA_signal_31164 ;
    wire new_AGEMA_signal_31165 ;
    wire new_AGEMA_signal_31166 ;
    wire new_AGEMA_signal_31167 ;
    wire new_AGEMA_signal_31168 ;
    wire new_AGEMA_signal_31169 ;
    wire new_AGEMA_signal_31170 ;
    wire new_AGEMA_signal_31171 ;
    wire new_AGEMA_signal_31172 ;
    wire new_AGEMA_signal_31173 ;
    wire new_AGEMA_signal_31174 ;
    wire new_AGEMA_signal_31175 ;
    wire new_AGEMA_signal_31176 ;
    wire new_AGEMA_signal_31177 ;
    wire new_AGEMA_signal_31178 ;
    wire new_AGEMA_signal_31179 ;
    wire new_AGEMA_signal_31180 ;
    wire new_AGEMA_signal_31181 ;
    wire new_AGEMA_signal_31182 ;
    wire new_AGEMA_signal_31183 ;
    wire new_AGEMA_signal_31184 ;
    wire new_AGEMA_signal_31185 ;
    wire new_AGEMA_signal_31186 ;
    wire new_AGEMA_signal_31187 ;
    wire new_AGEMA_signal_31188 ;
    wire new_AGEMA_signal_31189 ;
    wire new_AGEMA_signal_31190 ;
    wire new_AGEMA_signal_31191 ;
    wire new_AGEMA_signal_31192 ;
    wire new_AGEMA_signal_31193 ;
    wire new_AGEMA_signal_31194 ;
    wire new_AGEMA_signal_31195 ;
    wire new_AGEMA_signal_31196 ;
    wire new_AGEMA_signal_31197 ;
    wire new_AGEMA_signal_31198 ;
    wire new_AGEMA_signal_31199 ;
    wire new_AGEMA_signal_31200 ;
    wire new_AGEMA_signal_31201 ;
    wire new_AGEMA_signal_31202 ;
    wire new_AGEMA_signal_31203 ;
    wire new_AGEMA_signal_31204 ;
    wire new_AGEMA_signal_31205 ;
    wire new_AGEMA_signal_31206 ;
    wire new_AGEMA_signal_31207 ;
    wire new_AGEMA_signal_31208 ;
    wire new_AGEMA_signal_31209 ;
    wire new_AGEMA_signal_31210 ;
    wire new_AGEMA_signal_31211 ;
    wire new_AGEMA_signal_31212 ;
    wire new_AGEMA_signal_31213 ;
    wire new_AGEMA_signal_31214 ;
    wire new_AGEMA_signal_31215 ;
    wire new_AGEMA_signal_31216 ;
    wire new_AGEMA_signal_31217 ;
    wire new_AGEMA_signal_31218 ;
    wire new_AGEMA_signal_31219 ;
    wire new_AGEMA_signal_31220 ;
    wire new_AGEMA_signal_31221 ;
    wire new_AGEMA_signal_31222 ;
    wire new_AGEMA_signal_31223 ;
    wire new_AGEMA_signal_31224 ;
    wire new_AGEMA_signal_31225 ;
    wire new_AGEMA_signal_31226 ;
    wire new_AGEMA_signal_31227 ;
    wire new_AGEMA_signal_31228 ;
    wire new_AGEMA_signal_31229 ;
    wire new_AGEMA_signal_31230 ;
    wire new_AGEMA_signal_31231 ;
    wire new_AGEMA_signal_31232 ;
    wire new_AGEMA_signal_31233 ;
    wire new_AGEMA_signal_31234 ;
    wire new_AGEMA_signal_31235 ;
    wire new_AGEMA_signal_31236 ;
    wire new_AGEMA_signal_31237 ;
    wire new_AGEMA_signal_31238 ;
    wire new_AGEMA_signal_31239 ;
    wire new_AGEMA_signal_31240 ;
    wire new_AGEMA_signal_31241 ;
    wire new_AGEMA_signal_31242 ;
    wire new_AGEMA_signal_31243 ;
    wire new_AGEMA_signal_31244 ;
    wire new_AGEMA_signal_31245 ;
    wire new_AGEMA_signal_31246 ;
    wire new_AGEMA_signal_31247 ;
    wire new_AGEMA_signal_31248 ;
    wire new_AGEMA_signal_31249 ;
    wire new_AGEMA_signal_31250 ;
    wire new_AGEMA_signal_31251 ;
    wire new_AGEMA_signal_31252 ;
    wire new_AGEMA_signal_31253 ;
    wire new_AGEMA_signal_31254 ;
    wire new_AGEMA_signal_31255 ;
    wire new_AGEMA_signal_31256 ;
    wire new_AGEMA_signal_31257 ;
    wire new_AGEMA_signal_31258 ;
    wire new_AGEMA_signal_31259 ;
    wire new_AGEMA_signal_31260 ;
    wire new_AGEMA_signal_31261 ;
    wire new_AGEMA_signal_31262 ;
    wire new_AGEMA_signal_31263 ;
    wire new_AGEMA_signal_31264 ;
    wire new_AGEMA_signal_31265 ;
    wire new_AGEMA_signal_31266 ;
    wire new_AGEMA_signal_31267 ;
    wire new_AGEMA_signal_31268 ;
    wire new_AGEMA_signal_31269 ;
    wire new_AGEMA_signal_31270 ;
    wire new_AGEMA_signal_31271 ;
    wire new_AGEMA_signal_31272 ;
    wire new_AGEMA_signal_31273 ;
    wire new_AGEMA_signal_31274 ;
    wire new_AGEMA_signal_31275 ;
    wire new_AGEMA_signal_31276 ;
    wire new_AGEMA_signal_31277 ;
    wire new_AGEMA_signal_31278 ;
    wire new_AGEMA_signal_31279 ;
    wire new_AGEMA_signal_31280 ;
    wire new_AGEMA_signal_31281 ;
    wire new_AGEMA_signal_31282 ;
    wire new_AGEMA_signal_31283 ;
    wire new_AGEMA_signal_31284 ;
    wire new_AGEMA_signal_31285 ;
    wire new_AGEMA_signal_31286 ;
    wire new_AGEMA_signal_31287 ;
    wire new_AGEMA_signal_31288 ;
    wire new_AGEMA_signal_31289 ;
    wire new_AGEMA_signal_31290 ;
    wire new_AGEMA_signal_31291 ;
    wire new_AGEMA_signal_31292 ;
    wire new_AGEMA_signal_31293 ;
    wire new_AGEMA_signal_31294 ;
    wire new_AGEMA_signal_31295 ;
    wire new_AGEMA_signal_31296 ;
    wire new_AGEMA_signal_31297 ;
    wire new_AGEMA_signal_31298 ;
    wire new_AGEMA_signal_31299 ;
    wire new_AGEMA_signal_31300 ;
    wire new_AGEMA_signal_31301 ;
    wire new_AGEMA_signal_31302 ;
    wire new_AGEMA_signal_31303 ;
    wire new_AGEMA_signal_31304 ;
    wire new_AGEMA_signal_31305 ;
    wire new_AGEMA_signal_31306 ;
    wire new_AGEMA_signal_31307 ;
    wire new_AGEMA_signal_31308 ;
    wire new_AGEMA_signal_31309 ;
    wire new_AGEMA_signal_31310 ;
    wire new_AGEMA_signal_31311 ;
    wire new_AGEMA_signal_31312 ;
    wire new_AGEMA_signal_31313 ;
    wire new_AGEMA_signal_31314 ;
    wire new_AGEMA_signal_31315 ;
    wire new_AGEMA_signal_31316 ;
    wire new_AGEMA_signal_31317 ;
    wire new_AGEMA_signal_31318 ;
    wire new_AGEMA_signal_31319 ;
    wire new_AGEMA_signal_31320 ;
    wire new_AGEMA_signal_31321 ;
    wire new_AGEMA_signal_31322 ;
    wire new_AGEMA_signal_31323 ;
    wire new_AGEMA_signal_31324 ;
    wire new_AGEMA_signal_31325 ;
    wire new_AGEMA_signal_31326 ;
    wire new_AGEMA_signal_31327 ;
    wire new_AGEMA_signal_31328 ;
    wire new_AGEMA_signal_31329 ;
    wire new_AGEMA_signal_31330 ;
    wire new_AGEMA_signal_31331 ;
    wire new_AGEMA_signal_31332 ;
    wire new_AGEMA_signal_31333 ;
    wire new_AGEMA_signal_31334 ;
    wire new_AGEMA_signal_31335 ;
    wire new_AGEMA_signal_31336 ;
    wire new_AGEMA_signal_31337 ;
    wire new_AGEMA_signal_31338 ;
    wire new_AGEMA_signal_31339 ;
    wire new_AGEMA_signal_31340 ;
    wire new_AGEMA_signal_31341 ;
    wire new_AGEMA_signal_31342 ;
    wire new_AGEMA_signal_31343 ;
    wire new_AGEMA_signal_31344 ;
    wire new_AGEMA_signal_31345 ;
    wire new_AGEMA_signal_31346 ;
    wire new_AGEMA_signal_31347 ;
    wire new_AGEMA_signal_31348 ;
    wire new_AGEMA_signal_31349 ;
    wire new_AGEMA_signal_31350 ;
    wire new_AGEMA_signal_31351 ;
    wire new_AGEMA_signal_31352 ;
    wire new_AGEMA_signal_31353 ;
    wire new_AGEMA_signal_31354 ;
    wire new_AGEMA_signal_31355 ;
    wire new_AGEMA_signal_31356 ;
    wire new_AGEMA_signal_31357 ;
    wire new_AGEMA_signal_31358 ;
    wire new_AGEMA_signal_31359 ;
    wire new_AGEMA_signal_31360 ;
    wire new_AGEMA_signal_31361 ;
    wire new_AGEMA_signal_31362 ;
    wire new_AGEMA_signal_31363 ;
    wire new_AGEMA_signal_31364 ;
    wire new_AGEMA_signal_31365 ;
    wire new_AGEMA_signal_31366 ;
    wire new_AGEMA_signal_31367 ;
    wire new_AGEMA_signal_31368 ;
    wire new_AGEMA_signal_31369 ;
    wire new_AGEMA_signal_31370 ;
    wire new_AGEMA_signal_31371 ;
    wire new_AGEMA_signal_31372 ;
    wire new_AGEMA_signal_31373 ;
    wire new_AGEMA_signal_31374 ;
    wire new_AGEMA_signal_31375 ;
    wire new_AGEMA_signal_31376 ;
    wire new_AGEMA_signal_31377 ;
    wire new_AGEMA_signal_31378 ;
    wire new_AGEMA_signal_31379 ;
    wire new_AGEMA_signal_31380 ;
    wire new_AGEMA_signal_31381 ;
    wire new_AGEMA_signal_31382 ;
    wire new_AGEMA_signal_31383 ;
    wire new_AGEMA_signal_31384 ;
    wire new_AGEMA_signal_31385 ;
    wire new_AGEMA_signal_31386 ;
    wire new_AGEMA_signal_31387 ;
    wire new_AGEMA_signal_31388 ;
    wire new_AGEMA_signal_31389 ;
    wire new_AGEMA_signal_31390 ;
    wire new_AGEMA_signal_31391 ;
    wire new_AGEMA_signal_31392 ;
    wire new_AGEMA_signal_31393 ;
    wire new_AGEMA_signal_31394 ;
    wire new_AGEMA_signal_31395 ;
    wire new_AGEMA_signal_31396 ;
    wire new_AGEMA_signal_31397 ;
    wire new_AGEMA_signal_31398 ;
    wire new_AGEMA_signal_31399 ;
    wire new_AGEMA_signal_31400 ;
    wire new_AGEMA_signal_31401 ;
    wire new_AGEMA_signal_31402 ;
    wire new_AGEMA_signal_31403 ;
    wire new_AGEMA_signal_31404 ;
    wire new_AGEMA_signal_31405 ;
    wire new_AGEMA_signal_31406 ;
    wire new_AGEMA_signal_31407 ;
    wire new_AGEMA_signal_31408 ;
    wire new_AGEMA_signal_31409 ;
    wire new_AGEMA_signal_31410 ;
    wire new_AGEMA_signal_31411 ;
    wire new_AGEMA_signal_31412 ;
    wire new_AGEMA_signal_31413 ;
    wire new_AGEMA_signal_31414 ;
    wire new_AGEMA_signal_31415 ;
    wire new_AGEMA_signal_31416 ;
    wire new_AGEMA_signal_31417 ;
    wire new_AGEMA_signal_31418 ;
    wire new_AGEMA_signal_31419 ;
    wire new_AGEMA_signal_31420 ;
    wire new_AGEMA_signal_31421 ;
    wire new_AGEMA_signal_31422 ;
    wire new_AGEMA_signal_31423 ;
    wire new_AGEMA_signal_31424 ;
    wire new_AGEMA_signal_31425 ;
    wire new_AGEMA_signal_31426 ;
    wire new_AGEMA_signal_31427 ;
    wire new_AGEMA_signal_31428 ;
    wire new_AGEMA_signal_31429 ;
    wire new_AGEMA_signal_31430 ;
    wire new_AGEMA_signal_31431 ;
    wire new_AGEMA_signal_31432 ;
    wire new_AGEMA_signal_31433 ;
    wire new_AGEMA_signal_31434 ;
    wire new_AGEMA_signal_31435 ;
    wire new_AGEMA_signal_31436 ;
    wire new_AGEMA_signal_31437 ;
    wire new_AGEMA_signal_31438 ;
    wire new_AGEMA_signal_31439 ;
    wire new_AGEMA_signal_31440 ;
    wire new_AGEMA_signal_31441 ;
    wire new_AGEMA_signal_31442 ;
    wire new_AGEMA_signal_31443 ;
    wire new_AGEMA_signal_31444 ;
    wire new_AGEMA_signal_31445 ;
    wire new_AGEMA_signal_31446 ;
    wire new_AGEMA_signal_31447 ;
    wire new_AGEMA_signal_31448 ;
    wire new_AGEMA_signal_31449 ;
    wire new_AGEMA_signal_31450 ;
    wire new_AGEMA_signal_31451 ;
    wire new_AGEMA_signal_31452 ;
    wire new_AGEMA_signal_31453 ;
    wire new_AGEMA_signal_31454 ;
    wire new_AGEMA_signal_31455 ;
    wire new_AGEMA_signal_31456 ;
    wire new_AGEMA_signal_31457 ;
    wire new_AGEMA_signal_31458 ;
    wire new_AGEMA_signal_31459 ;
    wire new_AGEMA_signal_31460 ;
    wire new_AGEMA_signal_31461 ;
    wire new_AGEMA_signal_31462 ;
    wire new_AGEMA_signal_31463 ;
    wire new_AGEMA_signal_31464 ;
    wire new_AGEMA_signal_31465 ;
    wire new_AGEMA_signal_31466 ;
    wire new_AGEMA_signal_31467 ;
    wire new_AGEMA_signal_31468 ;
    wire new_AGEMA_signal_31469 ;
    wire new_AGEMA_signal_31470 ;
    wire new_AGEMA_signal_31471 ;
    wire new_AGEMA_signal_31472 ;
    wire new_AGEMA_signal_31473 ;
    wire new_AGEMA_signal_31474 ;
    wire new_AGEMA_signal_31475 ;
    wire new_AGEMA_signal_31476 ;
    wire new_AGEMA_signal_31477 ;
    wire new_AGEMA_signal_31478 ;
    wire new_AGEMA_signal_31479 ;
    wire new_AGEMA_signal_31480 ;
    wire new_AGEMA_signal_31481 ;
    wire new_AGEMA_signal_31482 ;
    wire new_AGEMA_signal_31483 ;
    wire new_AGEMA_signal_31484 ;
    wire new_AGEMA_signal_31485 ;
    wire new_AGEMA_signal_31486 ;
    wire new_AGEMA_signal_31487 ;
    wire new_AGEMA_signal_31488 ;
    wire new_AGEMA_signal_31489 ;
    wire new_AGEMA_signal_31490 ;
    wire new_AGEMA_signal_31491 ;
    wire new_AGEMA_signal_31492 ;
    wire new_AGEMA_signal_31493 ;
    wire new_AGEMA_signal_31494 ;
    wire new_AGEMA_signal_31495 ;
    wire new_AGEMA_signal_31496 ;
    wire new_AGEMA_signal_31497 ;
    wire new_AGEMA_signal_31498 ;
    wire new_AGEMA_signal_31499 ;
    wire new_AGEMA_signal_31500 ;
    wire new_AGEMA_signal_31501 ;
    wire new_AGEMA_signal_31502 ;
    wire new_AGEMA_signal_31503 ;
    wire new_AGEMA_signal_31504 ;
    wire new_AGEMA_signal_31505 ;
    wire new_AGEMA_signal_31506 ;
    wire new_AGEMA_signal_31507 ;
    wire new_AGEMA_signal_31508 ;
    wire new_AGEMA_signal_31509 ;
    wire new_AGEMA_signal_31510 ;
    wire new_AGEMA_signal_31511 ;
    wire new_AGEMA_signal_31512 ;
    wire new_AGEMA_signal_31513 ;
    wire new_AGEMA_signal_31514 ;
    wire new_AGEMA_signal_31515 ;
    wire new_AGEMA_signal_31516 ;
    wire new_AGEMA_signal_31517 ;
    wire new_AGEMA_signal_31518 ;
    wire new_AGEMA_signal_31519 ;
    wire new_AGEMA_signal_31520 ;
    wire new_AGEMA_signal_31521 ;
    wire new_AGEMA_signal_31522 ;
    wire new_AGEMA_signal_31523 ;
    wire new_AGEMA_signal_31524 ;
    wire new_AGEMA_signal_31525 ;
    wire new_AGEMA_signal_31526 ;
    wire new_AGEMA_signal_31527 ;
    wire new_AGEMA_signal_31528 ;
    wire new_AGEMA_signal_31529 ;
    wire new_AGEMA_signal_31530 ;
    wire new_AGEMA_signal_31531 ;
    wire new_AGEMA_signal_31532 ;
    wire new_AGEMA_signal_31533 ;
    wire new_AGEMA_signal_31534 ;
    wire new_AGEMA_signal_31535 ;
    wire new_AGEMA_signal_31536 ;
    wire new_AGEMA_signal_31537 ;
    wire new_AGEMA_signal_31538 ;
    wire new_AGEMA_signal_31539 ;
    wire new_AGEMA_signal_31540 ;
    wire new_AGEMA_signal_31541 ;
    wire new_AGEMA_signal_31542 ;
    wire new_AGEMA_signal_31543 ;
    wire new_AGEMA_signal_31544 ;
    wire new_AGEMA_signal_31545 ;
    wire new_AGEMA_signal_31546 ;
    wire new_AGEMA_signal_31547 ;
    wire new_AGEMA_signal_31548 ;
    wire new_AGEMA_signal_31549 ;
    wire new_AGEMA_signal_31550 ;
    wire new_AGEMA_signal_31551 ;
    wire new_AGEMA_signal_31552 ;
    wire new_AGEMA_signal_31553 ;
    wire new_AGEMA_signal_31554 ;
    wire new_AGEMA_signal_31555 ;
    wire new_AGEMA_signal_31556 ;
    wire new_AGEMA_signal_31557 ;
    wire new_AGEMA_signal_31558 ;
    wire new_AGEMA_signal_31559 ;
    wire new_AGEMA_signal_31560 ;
    wire new_AGEMA_signal_31561 ;
    wire new_AGEMA_signal_31562 ;
    wire new_AGEMA_signal_31563 ;
    wire new_AGEMA_signal_31564 ;
    wire new_AGEMA_signal_31565 ;
    wire new_AGEMA_signal_31566 ;
    wire new_AGEMA_signal_31567 ;
    wire new_AGEMA_signal_31568 ;
    wire new_AGEMA_signal_31569 ;
    wire new_AGEMA_signal_31570 ;
    wire new_AGEMA_signal_31571 ;
    wire new_AGEMA_signal_31572 ;
    wire new_AGEMA_signal_31573 ;
    wire new_AGEMA_signal_31574 ;
    wire new_AGEMA_signal_31575 ;
    wire new_AGEMA_signal_31576 ;
    wire new_AGEMA_signal_31577 ;
    wire new_AGEMA_signal_31578 ;
    wire new_AGEMA_signal_31579 ;
    wire new_AGEMA_signal_31580 ;
    wire new_AGEMA_signal_31581 ;
    wire new_AGEMA_signal_31582 ;
    wire new_AGEMA_signal_31583 ;
    wire new_AGEMA_signal_31584 ;
    wire new_AGEMA_signal_31585 ;
    wire new_AGEMA_signal_31586 ;
    wire new_AGEMA_signal_31587 ;
    wire new_AGEMA_signal_31588 ;
    wire new_AGEMA_signal_31589 ;
    wire new_AGEMA_signal_31590 ;
    wire new_AGEMA_signal_31591 ;
    wire new_AGEMA_signal_31592 ;
    wire new_AGEMA_signal_31593 ;
    wire new_AGEMA_signal_31594 ;
    wire new_AGEMA_signal_31595 ;
    wire new_AGEMA_signal_31596 ;
    wire new_AGEMA_signal_31597 ;
    wire new_AGEMA_signal_31598 ;
    wire new_AGEMA_signal_31599 ;
    wire new_AGEMA_signal_31600 ;
    wire new_AGEMA_signal_31601 ;
    wire new_AGEMA_signal_31602 ;
    wire new_AGEMA_signal_31603 ;
    wire new_AGEMA_signal_31604 ;
    wire new_AGEMA_signal_31605 ;
    wire new_AGEMA_signal_31606 ;
    wire new_AGEMA_signal_31607 ;
    wire new_AGEMA_signal_31608 ;
    wire new_AGEMA_signal_31609 ;
    wire new_AGEMA_signal_31610 ;
    wire new_AGEMA_signal_31611 ;
    wire new_AGEMA_signal_31612 ;
    wire new_AGEMA_signal_31613 ;
    wire new_AGEMA_signal_31614 ;
    wire new_AGEMA_signal_31615 ;
    wire new_AGEMA_signal_31616 ;
    wire new_AGEMA_signal_31617 ;
    wire new_AGEMA_signal_31618 ;
    wire new_AGEMA_signal_31619 ;
    wire new_AGEMA_signal_31620 ;
    wire new_AGEMA_signal_31621 ;
    wire new_AGEMA_signal_31622 ;
    wire new_AGEMA_signal_31623 ;
    wire new_AGEMA_signal_31624 ;
    wire new_AGEMA_signal_31625 ;
    wire new_AGEMA_signal_31626 ;
    wire new_AGEMA_signal_31627 ;
    wire new_AGEMA_signal_31628 ;
    wire new_AGEMA_signal_31629 ;
    wire new_AGEMA_signal_31630 ;
    wire new_AGEMA_signal_31631 ;
    wire new_AGEMA_signal_31632 ;
    wire new_AGEMA_signal_31633 ;
    wire new_AGEMA_signal_31634 ;
    wire new_AGEMA_signal_31635 ;
    wire new_AGEMA_signal_31636 ;
    wire new_AGEMA_signal_31637 ;
    wire new_AGEMA_signal_31638 ;
    wire new_AGEMA_signal_31639 ;
    wire new_AGEMA_signal_31640 ;
    wire new_AGEMA_signal_31641 ;
    wire new_AGEMA_signal_31642 ;
    wire new_AGEMA_signal_31643 ;
    wire new_AGEMA_signal_31644 ;
    wire new_AGEMA_signal_31645 ;
    wire new_AGEMA_signal_31646 ;
    wire new_AGEMA_signal_31647 ;
    wire new_AGEMA_signal_31648 ;
    wire new_AGEMA_signal_31649 ;
    wire new_AGEMA_signal_31650 ;
    wire new_AGEMA_signal_31651 ;
    wire new_AGEMA_signal_31652 ;
    wire new_AGEMA_signal_31653 ;
    wire new_AGEMA_signal_31654 ;
    wire new_AGEMA_signal_31655 ;
    wire new_AGEMA_signal_31656 ;
    wire new_AGEMA_signal_31657 ;
    wire new_AGEMA_signal_31658 ;
    wire new_AGEMA_signal_31659 ;
    wire new_AGEMA_signal_31660 ;
    wire new_AGEMA_signal_31661 ;
    wire new_AGEMA_signal_31662 ;
    wire new_AGEMA_signal_31663 ;
    wire new_AGEMA_signal_31664 ;
    wire new_AGEMA_signal_31665 ;
    wire new_AGEMA_signal_31666 ;
    wire new_AGEMA_signal_31667 ;
    wire new_AGEMA_signal_31668 ;
    wire new_AGEMA_signal_31669 ;
    wire new_AGEMA_signal_31670 ;
    wire new_AGEMA_signal_31671 ;
    wire new_AGEMA_signal_31672 ;
    wire new_AGEMA_signal_31673 ;
    wire new_AGEMA_signal_31674 ;
    wire new_AGEMA_signal_31675 ;
    wire new_AGEMA_signal_31676 ;
    wire new_AGEMA_signal_31677 ;
    wire new_AGEMA_signal_31678 ;
    wire new_AGEMA_signal_31679 ;
    wire new_AGEMA_signal_31680 ;
    wire new_AGEMA_signal_31681 ;
    wire new_AGEMA_signal_31682 ;
    wire new_AGEMA_signal_31683 ;
    wire new_AGEMA_signal_31684 ;
    wire new_AGEMA_signal_31685 ;
    wire new_AGEMA_signal_31686 ;
    wire new_AGEMA_signal_31687 ;
    wire new_AGEMA_signal_31688 ;
    wire new_AGEMA_signal_31689 ;
    wire new_AGEMA_signal_31690 ;
    wire new_AGEMA_signal_31691 ;
    wire new_AGEMA_signal_31692 ;
    wire new_AGEMA_signal_31693 ;
    wire new_AGEMA_signal_31694 ;
    wire new_AGEMA_signal_31695 ;
    wire new_AGEMA_signal_31696 ;
    wire new_AGEMA_signal_31697 ;
    wire new_AGEMA_signal_31698 ;
    wire new_AGEMA_signal_31699 ;
    wire new_AGEMA_signal_31700 ;
    wire new_AGEMA_signal_31701 ;
    wire new_AGEMA_signal_31702 ;
    wire new_AGEMA_signal_31703 ;
    wire new_AGEMA_signal_31704 ;
    wire new_AGEMA_signal_31705 ;
    wire new_AGEMA_signal_31706 ;
    wire new_AGEMA_signal_31707 ;
    wire new_AGEMA_signal_31708 ;
    wire new_AGEMA_signal_31709 ;
    wire new_AGEMA_signal_31710 ;
    wire new_AGEMA_signal_31711 ;
    wire new_AGEMA_signal_31712 ;
    wire new_AGEMA_signal_31713 ;
    wire new_AGEMA_signal_31714 ;
    wire new_AGEMA_signal_31715 ;
    wire new_AGEMA_signal_31716 ;
    wire new_AGEMA_signal_31717 ;
    wire new_AGEMA_signal_31718 ;
    wire new_AGEMA_signal_31719 ;
    wire new_AGEMA_signal_31720 ;
    wire new_AGEMA_signal_31721 ;
    wire new_AGEMA_signal_31722 ;
    wire new_AGEMA_signal_31723 ;
    wire new_AGEMA_signal_31724 ;
    wire new_AGEMA_signal_31725 ;
    wire new_AGEMA_signal_31726 ;
    wire new_AGEMA_signal_31727 ;
    wire new_AGEMA_signal_31728 ;
    wire new_AGEMA_signal_31729 ;
    wire new_AGEMA_signal_31730 ;
    wire new_AGEMA_signal_31731 ;
    wire new_AGEMA_signal_31732 ;
    wire new_AGEMA_signal_31733 ;
    wire new_AGEMA_signal_31734 ;
    wire new_AGEMA_signal_31735 ;
    wire new_AGEMA_signal_31736 ;
    wire new_AGEMA_signal_31737 ;
    wire new_AGEMA_signal_31738 ;
    wire new_AGEMA_signal_31739 ;
    wire new_AGEMA_signal_31740 ;
    wire new_AGEMA_signal_31741 ;
    wire new_AGEMA_signal_31742 ;
    wire new_AGEMA_signal_31743 ;
    wire new_AGEMA_signal_31744 ;
    wire new_AGEMA_signal_31745 ;
    wire new_AGEMA_signal_31746 ;
    wire new_AGEMA_signal_31747 ;
    wire new_AGEMA_signal_31748 ;
    wire new_AGEMA_signal_31749 ;
    wire new_AGEMA_signal_31750 ;
    wire new_AGEMA_signal_31751 ;
    wire new_AGEMA_signal_31752 ;
    wire new_AGEMA_signal_31753 ;
    wire new_AGEMA_signal_31754 ;
    wire new_AGEMA_signal_31755 ;
    wire new_AGEMA_signal_31756 ;
    wire new_AGEMA_signal_31757 ;
    wire new_AGEMA_signal_31758 ;
    wire new_AGEMA_signal_31759 ;
    wire new_AGEMA_signal_31760 ;
    wire new_AGEMA_signal_31761 ;
    wire new_AGEMA_signal_31762 ;
    wire new_AGEMA_signal_31763 ;
    wire new_AGEMA_signal_31764 ;
    wire new_AGEMA_signal_31765 ;
    wire new_AGEMA_signal_31766 ;
    wire new_AGEMA_signal_31767 ;
    wire new_AGEMA_signal_31768 ;
    wire new_AGEMA_signal_31769 ;
    wire new_AGEMA_signal_31770 ;
    wire new_AGEMA_signal_31771 ;
    wire new_AGEMA_signal_31772 ;
    wire new_AGEMA_signal_31773 ;
    wire new_AGEMA_signal_31774 ;
    wire new_AGEMA_signal_31775 ;
    wire new_AGEMA_signal_31776 ;
    wire new_AGEMA_signal_31777 ;
    wire new_AGEMA_signal_31778 ;
    wire new_AGEMA_signal_31779 ;
    wire new_AGEMA_signal_31780 ;
    wire new_AGEMA_signal_31781 ;
    wire new_AGEMA_signal_31782 ;
    wire new_AGEMA_signal_31783 ;
    wire new_AGEMA_signal_31784 ;
    wire new_AGEMA_signal_31785 ;
    wire new_AGEMA_signal_31786 ;
    wire new_AGEMA_signal_31787 ;
    wire new_AGEMA_signal_31788 ;
    wire new_AGEMA_signal_31789 ;
    wire new_AGEMA_signal_31790 ;
    wire new_AGEMA_signal_31791 ;
    wire new_AGEMA_signal_31792 ;
    wire new_AGEMA_signal_31793 ;
    wire new_AGEMA_signal_31794 ;
    wire new_AGEMA_signal_31795 ;
    wire new_AGEMA_signal_31796 ;
    wire new_AGEMA_signal_31797 ;
    wire new_AGEMA_signal_31798 ;
    wire new_AGEMA_signal_31799 ;
    wire new_AGEMA_signal_31800 ;
    wire new_AGEMA_signal_31801 ;
    wire new_AGEMA_signal_31802 ;
    wire new_AGEMA_signal_31803 ;
    wire new_AGEMA_signal_31804 ;
    wire new_AGEMA_signal_31805 ;
    wire new_AGEMA_signal_31806 ;
    wire new_AGEMA_signal_31807 ;
    wire new_AGEMA_signal_31808 ;
    wire new_AGEMA_signal_31809 ;
    wire new_AGEMA_signal_31810 ;
    wire new_AGEMA_signal_31811 ;
    wire new_AGEMA_signal_31812 ;
    wire new_AGEMA_signal_31813 ;
    wire new_AGEMA_signal_31814 ;
    wire new_AGEMA_signal_31815 ;
    wire new_AGEMA_signal_31816 ;
    wire new_AGEMA_signal_31817 ;
    wire new_AGEMA_signal_31818 ;
    wire new_AGEMA_signal_31819 ;
    wire new_AGEMA_signal_31820 ;
    wire new_AGEMA_signal_31821 ;
    wire new_AGEMA_signal_31822 ;
    wire new_AGEMA_signal_31823 ;
    wire new_AGEMA_signal_31824 ;
    wire new_AGEMA_signal_31825 ;
    wire new_AGEMA_signal_31826 ;
    wire new_AGEMA_signal_31827 ;
    wire new_AGEMA_signal_31828 ;
    wire new_AGEMA_signal_31829 ;
    wire new_AGEMA_signal_31830 ;
    wire new_AGEMA_signal_31831 ;
    wire new_AGEMA_signal_31832 ;
    wire new_AGEMA_signal_31833 ;
    wire new_AGEMA_signal_31834 ;
    wire new_AGEMA_signal_31835 ;
    wire new_AGEMA_signal_31836 ;
    wire new_AGEMA_signal_31837 ;
    wire new_AGEMA_signal_31838 ;
    wire new_AGEMA_signal_31839 ;
    wire new_AGEMA_signal_31840 ;
    wire new_AGEMA_signal_31841 ;
    wire new_AGEMA_signal_31842 ;
    wire new_AGEMA_signal_31843 ;
    wire new_AGEMA_signal_31844 ;
    wire new_AGEMA_signal_31845 ;
    wire new_AGEMA_signal_31846 ;
    wire new_AGEMA_signal_31847 ;
    wire new_AGEMA_signal_31848 ;
    wire new_AGEMA_signal_31849 ;
    wire new_AGEMA_signal_31850 ;
    wire new_AGEMA_signal_31851 ;
    wire new_AGEMA_signal_31852 ;
    wire new_AGEMA_signal_31853 ;
    wire new_AGEMA_signal_31854 ;
    wire new_AGEMA_signal_31855 ;
    wire new_AGEMA_signal_31856 ;
    wire new_AGEMA_signal_31857 ;
    wire new_AGEMA_signal_31858 ;
    wire new_AGEMA_signal_31859 ;
    wire new_AGEMA_signal_31860 ;
    wire new_AGEMA_signal_31861 ;
    wire new_AGEMA_signal_31862 ;
    wire new_AGEMA_signal_31863 ;
    wire new_AGEMA_signal_31864 ;
    wire new_AGEMA_signal_31865 ;
    wire new_AGEMA_signal_31866 ;
    wire new_AGEMA_signal_31867 ;
    wire new_AGEMA_signal_31868 ;
    wire new_AGEMA_signal_31869 ;
    wire new_AGEMA_signal_31870 ;
    wire new_AGEMA_signal_31871 ;
    wire new_AGEMA_signal_31872 ;
    wire new_AGEMA_signal_31873 ;
    wire new_AGEMA_signal_31874 ;
    wire new_AGEMA_signal_31875 ;
    wire new_AGEMA_signal_31876 ;
    wire new_AGEMA_signal_31877 ;
    wire new_AGEMA_signal_31878 ;
    wire new_AGEMA_signal_31879 ;
    wire new_AGEMA_signal_31880 ;
    wire new_AGEMA_signal_31881 ;
    wire new_AGEMA_signal_31882 ;
    wire new_AGEMA_signal_31883 ;
    wire new_AGEMA_signal_31884 ;
    wire new_AGEMA_signal_31885 ;
    wire new_AGEMA_signal_31886 ;
    wire new_AGEMA_signal_31887 ;
    wire new_AGEMA_signal_31888 ;
    wire new_AGEMA_signal_31889 ;
    wire new_AGEMA_signal_31890 ;
    wire new_AGEMA_signal_31891 ;
    wire new_AGEMA_signal_31892 ;
    wire new_AGEMA_signal_31893 ;
    wire new_AGEMA_signal_31894 ;
    wire new_AGEMA_signal_31895 ;
    wire new_AGEMA_signal_31896 ;
    wire new_AGEMA_signal_31897 ;
    wire new_AGEMA_signal_31898 ;
    wire new_AGEMA_signal_31899 ;
    wire new_AGEMA_signal_31900 ;
    wire new_AGEMA_signal_31901 ;
    wire new_AGEMA_signal_31902 ;
    wire new_AGEMA_signal_31903 ;
    wire new_AGEMA_signal_31904 ;
    wire new_AGEMA_signal_31905 ;
    wire new_AGEMA_signal_31906 ;
    wire new_AGEMA_signal_31907 ;
    wire new_AGEMA_signal_31908 ;
    wire new_AGEMA_signal_31909 ;
    wire new_AGEMA_signal_31910 ;
    wire new_AGEMA_signal_31911 ;
    wire new_AGEMA_signal_31912 ;
    wire new_AGEMA_signal_31913 ;
    wire new_AGEMA_signal_31914 ;
    wire new_AGEMA_signal_31915 ;
    wire new_AGEMA_signal_31916 ;
    wire new_AGEMA_signal_31917 ;
    wire new_AGEMA_signal_31918 ;
    wire new_AGEMA_signal_31919 ;
    wire new_AGEMA_signal_31920 ;
    wire new_AGEMA_signal_31921 ;
    wire new_AGEMA_signal_31922 ;
    wire new_AGEMA_signal_31923 ;
    wire new_AGEMA_signal_31924 ;
    wire new_AGEMA_signal_31925 ;
    wire new_AGEMA_signal_31926 ;
    wire new_AGEMA_signal_31927 ;
    wire new_AGEMA_signal_31928 ;
    wire new_AGEMA_signal_31929 ;
    wire new_AGEMA_signal_31930 ;
    wire new_AGEMA_signal_31931 ;
    wire new_AGEMA_signal_31932 ;
    wire new_AGEMA_signal_31933 ;
    wire new_AGEMA_signal_31934 ;
    wire new_AGEMA_signal_31935 ;
    wire new_AGEMA_signal_31936 ;
    wire new_AGEMA_signal_31937 ;
    wire new_AGEMA_signal_31938 ;
    wire new_AGEMA_signal_31939 ;
    wire new_AGEMA_signal_31940 ;
    wire new_AGEMA_signal_31941 ;
    wire new_AGEMA_signal_31942 ;
    wire new_AGEMA_signal_31943 ;
    wire new_AGEMA_signal_31944 ;
    wire new_AGEMA_signal_31945 ;
    wire new_AGEMA_signal_31946 ;
    wire new_AGEMA_signal_31947 ;
    wire new_AGEMA_signal_31948 ;
    wire new_AGEMA_signal_31949 ;
    wire new_AGEMA_signal_31950 ;
    wire new_AGEMA_signal_31951 ;
    wire new_AGEMA_signal_31952 ;
    wire new_AGEMA_signal_31953 ;
    wire new_AGEMA_signal_31954 ;
    wire new_AGEMA_signal_31955 ;
    wire new_AGEMA_signal_31956 ;
    wire new_AGEMA_signal_31957 ;
    wire new_AGEMA_signal_31958 ;
    wire new_AGEMA_signal_31959 ;
    wire new_AGEMA_signal_31960 ;
    wire new_AGEMA_signal_31961 ;
    wire new_AGEMA_signal_31962 ;
    wire new_AGEMA_signal_31963 ;
    wire new_AGEMA_signal_31964 ;
    wire new_AGEMA_signal_31965 ;
    wire new_AGEMA_signal_31966 ;
    wire new_AGEMA_signal_31967 ;
    wire new_AGEMA_signal_31968 ;
    wire new_AGEMA_signal_31969 ;
    wire new_AGEMA_signal_31970 ;
    wire new_AGEMA_signal_31971 ;
    wire new_AGEMA_signal_31972 ;
    wire new_AGEMA_signal_31973 ;
    wire new_AGEMA_signal_31974 ;
    wire new_AGEMA_signal_31975 ;
    wire new_AGEMA_signal_31976 ;
    wire new_AGEMA_signal_31977 ;
    wire new_AGEMA_signal_31978 ;
    wire new_AGEMA_signal_31979 ;
    wire new_AGEMA_signal_31980 ;
    wire new_AGEMA_signal_31981 ;
    wire new_AGEMA_signal_31982 ;
    wire new_AGEMA_signal_31983 ;
    wire new_AGEMA_signal_31984 ;
    wire new_AGEMA_signal_31985 ;
    wire new_AGEMA_signal_31986 ;
    wire new_AGEMA_signal_31987 ;
    wire new_AGEMA_signal_31988 ;
    wire new_AGEMA_signal_31989 ;
    wire new_AGEMA_signal_31990 ;
    wire new_AGEMA_signal_31991 ;
    wire new_AGEMA_signal_31992 ;
    wire new_AGEMA_signal_31993 ;
    wire new_AGEMA_signal_31994 ;
    wire new_AGEMA_signal_31995 ;
    wire new_AGEMA_signal_31996 ;
    wire new_AGEMA_signal_31997 ;
    wire new_AGEMA_signal_31998 ;
    wire new_AGEMA_signal_31999 ;
    wire new_AGEMA_signal_32000 ;
    wire new_AGEMA_signal_32001 ;
    wire new_AGEMA_signal_32002 ;
    wire new_AGEMA_signal_32003 ;
    wire new_AGEMA_signal_32004 ;
    wire new_AGEMA_signal_32005 ;
    wire new_AGEMA_signal_32006 ;
    wire new_AGEMA_signal_32007 ;
    wire new_AGEMA_signal_32008 ;
    wire new_AGEMA_signal_32009 ;
    wire new_AGEMA_signal_32010 ;
    wire new_AGEMA_signal_32011 ;
    wire new_AGEMA_signal_32012 ;
    wire new_AGEMA_signal_32013 ;
    wire new_AGEMA_signal_32014 ;
    wire new_AGEMA_signal_32015 ;
    wire new_AGEMA_signal_32016 ;
    wire new_AGEMA_signal_32017 ;
    wire new_AGEMA_signal_32018 ;
    wire new_AGEMA_signal_32019 ;
    wire new_AGEMA_signal_32020 ;
    wire new_AGEMA_signal_32021 ;
    wire new_AGEMA_signal_32022 ;
    wire new_AGEMA_signal_32023 ;
    wire new_AGEMA_signal_32024 ;
    wire new_AGEMA_signal_32025 ;
    wire new_AGEMA_signal_32026 ;
    wire new_AGEMA_signal_32027 ;
    wire new_AGEMA_signal_32028 ;
    wire new_AGEMA_signal_32029 ;
    wire new_AGEMA_signal_32030 ;
    wire new_AGEMA_signal_32031 ;
    wire new_AGEMA_signal_32032 ;
    wire new_AGEMA_signal_32033 ;
    wire new_AGEMA_signal_32034 ;
    wire new_AGEMA_signal_32035 ;
    wire new_AGEMA_signal_32036 ;
    wire new_AGEMA_signal_32037 ;
    wire new_AGEMA_signal_32038 ;
    wire new_AGEMA_signal_32039 ;
    wire new_AGEMA_signal_32040 ;
    wire new_AGEMA_signal_32041 ;
    wire new_AGEMA_signal_32042 ;
    wire new_AGEMA_signal_32043 ;
    wire new_AGEMA_signal_32044 ;
    wire new_AGEMA_signal_32045 ;
    wire new_AGEMA_signal_32046 ;
    wire new_AGEMA_signal_32047 ;
    wire new_AGEMA_signal_32048 ;
    wire new_AGEMA_signal_32049 ;
    wire new_AGEMA_signal_32050 ;
    wire new_AGEMA_signal_32051 ;
    wire new_AGEMA_signal_32052 ;
    wire new_AGEMA_signal_32053 ;
    wire new_AGEMA_signal_32054 ;
    wire new_AGEMA_signal_32055 ;
    wire new_AGEMA_signal_32056 ;
    wire new_AGEMA_signal_32057 ;
    wire new_AGEMA_signal_32058 ;
    wire new_AGEMA_signal_32059 ;
    wire new_AGEMA_signal_32060 ;
    wire new_AGEMA_signal_32061 ;
    wire new_AGEMA_signal_32062 ;
    wire new_AGEMA_signal_32063 ;
    wire new_AGEMA_signal_32064 ;
    wire new_AGEMA_signal_32065 ;
    wire new_AGEMA_signal_32066 ;
    wire new_AGEMA_signal_32067 ;
    wire new_AGEMA_signal_32068 ;
    wire new_AGEMA_signal_32069 ;
    wire new_AGEMA_signal_32070 ;
    wire new_AGEMA_signal_32071 ;
    wire new_AGEMA_signal_32072 ;
    wire new_AGEMA_signal_32073 ;
    wire new_AGEMA_signal_32074 ;
    wire new_AGEMA_signal_32075 ;
    wire new_AGEMA_signal_32076 ;
    wire new_AGEMA_signal_32077 ;
    wire new_AGEMA_signal_32078 ;
    wire new_AGEMA_signal_32079 ;
    wire new_AGEMA_signal_32080 ;
    wire new_AGEMA_signal_32081 ;
    wire new_AGEMA_signal_32082 ;
    wire new_AGEMA_signal_32083 ;
    wire new_AGEMA_signal_32084 ;
    wire new_AGEMA_signal_32085 ;
    wire new_AGEMA_signal_32086 ;
    wire new_AGEMA_signal_32087 ;
    wire new_AGEMA_signal_32088 ;
    wire new_AGEMA_signal_32089 ;
    wire new_AGEMA_signal_32090 ;
    wire new_AGEMA_signal_32091 ;
    wire new_AGEMA_signal_32092 ;
    wire new_AGEMA_signal_32093 ;
    wire new_AGEMA_signal_32094 ;
    wire new_AGEMA_signal_32095 ;
    wire new_AGEMA_signal_32096 ;
    wire new_AGEMA_signal_32097 ;
    wire new_AGEMA_signal_32098 ;
    wire new_AGEMA_signal_32099 ;
    wire new_AGEMA_signal_32100 ;
    wire new_AGEMA_signal_32101 ;
    wire new_AGEMA_signal_32102 ;
    wire new_AGEMA_signal_32103 ;
    wire new_AGEMA_signal_32104 ;
    wire new_AGEMA_signal_32105 ;
    wire new_AGEMA_signal_32106 ;
    wire new_AGEMA_signal_32107 ;
    wire new_AGEMA_signal_32108 ;
    wire new_AGEMA_signal_32109 ;
    wire new_AGEMA_signal_32110 ;
    wire new_AGEMA_signal_32111 ;
    wire new_AGEMA_signal_32112 ;
    wire new_AGEMA_signal_32113 ;
    wire new_AGEMA_signal_32114 ;
    wire new_AGEMA_signal_32115 ;
    wire new_AGEMA_signal_32116 ;
    wire new_AGEMA_signal_32117 ;
    wire new_AGEMA_signal_32118 ;
    wire new_AGEMA_signal_32119 ;
    wire new_AGEMA_signal_32120 ;
    wire new_AGEMA_signal_32121 ;
    wire new_AGEMA_signal_32122 ;
    wire new_AGEMA_signal_32123 ;
    wire new_AGEMA_signal_32124 ;
    wire new_AGEMA_signal_32125 ;
    wire new_AGEMA_signal_32126 ;
    wire new_AGEMA_signal_32127 ;
    wire new_AGEMA_signal_32128 ;
    wire new_AGEMA_signal_32129 ;
    wire new_AGEMA_signal_32130 ;
    wire new_AGEMA_signal_32131 ;
    wire new_AGEMA_signal_32132 ;
    wire new_AGEMA_signal_32133 ;
    wire new_AGEMA_signal_32134 ;
    wire new_AGEMA_signal_32135 ;
    wire new_AGEMA_signal_32136 ;
    wire new_AGEMA_signal_32137 ;
    wire new_AGEMA_signal_32138 ;
    wire new_AGEMA_signal_32139 ;
    wire new_AGEMA_signal_32140 ;
    wire new_AGEMA_signal_32141 ;
    wire new_AGEMA_signal_32142 ;
    wire new_AGEMA_signal_32143 ;
    wire new_AGEMA_signal_32144 ;
    wire new_AGEMA_signal_32145 ;
    wire new_AGEMA_signal_32146 ;
    wire new_AGEMA_signal_32147 ;
    wire new_AGEMA_signal_32148 ;
    wire new_AGEMA_signal_32149 ;
    wire new_AGEMA_signal_32150 ;
    wire new_AGEMA_signal_32151 ;
    wire new_AGEMA_signal_32152 ;
    wire new_AGEMA_signal_32153 ;
    wire new_AGEMA_signal_32154 ;
    wire new_AGEMA_signal_32155 ;
    wire new_AGEMA_signal_32156 ;
    wire new_AGEMA_signal_32157 ;
    wire new_AGEMA_signal_32158 ;
    wire new_AGEMA_signal_32159 ;
    wire new_AGEMA_signal_32160 ;
    wire new_AGEMA_signal_32161 ;
    wire new_AGEMA_signal_32162 ;
    wire new_AGEMA_signal_32163 ;
    wire new_AGEMA_signal_32164 ;
    wire new_AGEMA_signal_32165 ;
    wire new_AGEMA_signal_32166 ;
    wire new_AGEMA_signal_32167 ;
    wire new_AGEMA_signal_32168 ;
    wire new_AGEMA_signal_32169 ;
    wire new_AGEMA_signal_32170 ;
    wire new_AGEMA_signal_32171 ;
    wire new_AGEMA_signal_32172 ;
    wire new_AGEMA_signal_32173 ;
    wire new_AGEMA_signal_32174 ;
    wire new_AGEMA_signal_32175 ;
    wire new_AGEMA_signal_32176 ;
    wire new_AGEMA_signal_32177 ;
    wire new_AGEMA_signal_32178 ;
    wire new_AGEMA_signal_32179 ;
    wire new_AGEMA_signal_32180 ;
    wire new_AGEMA_signal_32181 ;
    wire new_AGEMA_signal_32182 ;
    wire new_AGEMA_signal_32183 ;
    wire new_AGEMA_signal_32184 ;
    wire new_AGEMA_signal_32185 ;
    wire new_AGEMA_signal_32186 ;
    wire new_AGEMA_signal_32187 ;
    wire new_AGEMA_signal_32188 ;
    wire new_AGEMA_signal_32189 ;
    wire new_AGEMA_signal_32190 ;
    wire new_AGEMA_signal_32191 ;
    wire new_AGEMA_signal_32192 ;
    wire new_AGEMA_signal_32193 ;
    wire new_AGEMA_signal_32194 ;
    wire new_AGEMA_signal_32195 ;
    wire new_AGEMA_signal_32196 ;
    wire new_AGEMA_signal_32197 ;
    wire new_AGEMA_signal_32198 ;
    wire new_AGEMA_signal_32199 ;
    wire new_AGEMA_signal_32200 ;
    wire new_AGEMA_signal_32201 ;
    wire new_AGEMA_signal_32202 ;
    wire new_AGEMA_signal_32203 ;
    wire new_AGEMA_signal_32204 ;
    wire new_AGEMA_signal_32205 ;
    wire new_AGEMA_signal_32206 ;
    wire new_AGEMA_signal_32207 ;
    wire new_AGEMA_signal_32208 ;
    wire new_AGEMA_signal_32209 ;
    wire new_AGEMA_signal_32210 ;
    wire new_AGEMA_signal_32211 ;
    wire new_AGEMA_signal_32212 ;
    wire new_AGEMA_signal_32213 ;
    wire new_AGEMA_signal_32214 ;
    wire new_AGEMA_signal_32215 ;
    wire new_AGEMA_signal_32216 ;
    wire new_AGEMA_signal_32217 ;
    wire new_AGEMA_signal_32218 ;
    wire new_AGEMA_signal_32219 ;
    wire new_AGEMA_signal_32220 ;
    wire new_AGEMA_signal_32221 ;
    wire new_AGEMA_signal_32222 ;
    wire new_AGEMA_signal_32223 ;
    wire new_AGEMA_signal_32224 ;
    wire new_AGEMA_signal_32225 ;
    wire new_AGEMA_signal_32226 ;
    wire new_AGEMA_signal_32227 ;
    wire new_AGEMA_signal_32228 ;
    wire new_AGEMA_signal_32229 ;
    wire new_AGEMA_signal_32230 ;
    wire new_AGEMA_signal_32231 ;
    wire new_AGEMA_signal_32232 ;
    wire new_AGEMA_signal_32233 ;
    wire new_AGEMA_signal_32234 ;
    wire new_AGEMA_signal_32235 ;
    wire new_AGEMA_signal_32236 ;
    wire new_AGEMA_signal_32237 ;
    wire new_AGEMA_signal_32238 ;
    wire new_AGEMA_signal_32239 ;
    wire new_AGEMA_signal_32240 ;
    wire new_AGEMA_signal_32241 ;
    wire new_AGEMA_signal_32242 ;
    wire new_AGEMA_signal_32243 ;
    wire new_AGEMA_signal_32244 ;
    wire new_AGEMA_signal_32245 ;
    wire new_AGEMA_signal_32246 ;
    wire new_AGEMA_signal_32247 ;
    wire new_AGEMA_signal_32248 ;
    wire new_AGEMA_signal_32249 ;
    wire new_AGEMA_signal_32250 ;
    wire new_AGEMA_signal_32251 ;
    wire new_AGEMA_signal_32252 ;
    wire new_AGEMA_signal_32253 ;
    wire new_AGEMA_signal_32254 ;
    wire new_AGEMA_signal_32255 ;
    wire new_AGEMA_signal_32256 ;
    wire new_AGEMA_signal_32257 ;
    wire new_AGEMA_signal_32258 ;
    wire new_AGEMA_signal_32259 ;
    wire new_AGEMA_signal_32260 ;
    wire new_AGEMA_signal_32261 ;
    wire new_AGEMA_signal_32262 ;
    wire new_AGEMA_signal_32263 ;
    wire new_AGEMA_signal_32264 ;
    wire new_AGEMA_signal_32265 ;
    wire new_AGEMA_signal_32266 ;
    wire new_AGEMA_signal_32267 ;
    wire new_AGEMA_signal_32268 ;
    wire new_AGEMA_signal_32269 ;
    wire new_AGEMA_signal_32270 ;
    wire new_AGEMA_signal_32271 ;
    wire new_AGEMA_signal_32272 ;
    wire new_AGEMA_signal_32273 ;
    wire new_AGEMA_signal_32274 ;
    wire new_AGEMA_signal_32275 ;
    wire new_AGEMA_signal_32276 ;
    wire new_AGEMA_signal_32277 ;
    wire new_AGEMA_signal_32278 ;
    wire new_AGEMA_signal_32279 ;
    wire new_AGEMA_signal_32280 ;
    wire new_AGEMA_signal_32281 ;
    wire new_AGEMA_signal_32282 ;
    wire new_AGEMA_signal_32283 ;
    wire new_AGEMA_signal_32284 ;
    wire new_AGEMA_signal_32285 ;
    wire new_AGEMA_signal_32286 ;
    wire new_AGEMA_signal_32287 ;
    wire new_AGEMA_signal_32288 ;
    wire new_AGEMA_signal_32289 ;
    wire new_AGEMA_signal_32290 ;
    wire new_AGEMA_signal_32291 ;
    wire new_AGEMA_signal_32292 ;
    wire new_AGEMA_signal_32293 ;
    wire new_AGEMA_signal_32294 ;
    wire new_AGEMA_signal_32295 ;
    wire new_AGEMA_signal_32296 ;
    wire new_AGEMA_signal_32297 ;
    wire new_AGEMA_signal_32298 ;
    wire new_AGEMA_signal_32299 ;
    wire new_AGEMA_signal_32300 ;
    wire new_AGEMA_signal_32301 ;
    wire new_AGEMA_signal_32302 ;
    wire new_AGEMA_signal_32303 ;
    wire new_AGEMA_signal_32304 ;
    wire new_AGEMA_signal_32305 ;
    wire new_AGEMA_signal_32306 ;
    wire new_AGEMA_signal_32307 ;
    wire new_AGEMA_signal_32308 ;
    wire new_AGEMA_signal_32309 ;
    wire new_AGEMA_signal_32310 ;
    wire new_AGEMA_signal_32311 ;
    wire new_AGEMA_signal_32312 ;
    wire new_AGEMA_signal_32313 ;
    wire new_AGEMA_signal_32314 ;
    wire new_AGEMA_signal_32315 ;
    wire new_AGEMA_signal_32316 ;
    wire new_AGEMA_signal_32317 ;
    wire new_AGEMA_signal_32318 ;
    wire new_AGEMA_signal_32319 ;
    wire new_AGEMA_signal_32320 ;
    wire new_AGEMA_signal_32321 ;
    wire new_AGEMA_signal_32322 ;
    wire new_AGEMA_signal_32323 ;
    wire new_AGEMA_signal_32324 ;
    wire new_AGEMA_signal_32325 ;
    wire new_AGEMA_signal_32326 ;
    wire new_AGEMA_signal_32327 ;
    wire new_AGEMA_signal_32328 ;
    wire new_AGEMA_signal_32329 ;
    wire new_AGEMA_signal_32330 ;
    wire new_AGEMA_signal_32331 ;
    wire new_AGEMA_signal_32332 ;
    wire new_AGEMA_signal_32333 ;
    wire new_AGEMA_signal_32334 ;
    wire new_AGEMA_signal_32335 ;
    wire new_AGEMA_signal_32336 ;
    wire new_AGEMA_signal_32337 ;
    wire new_AGEMA_signal_32338 ;
    wire new_AGEMA_signal_32339 ;
    wire new_AGEMA_signal_32340 ;
    wire new_AGEMA_signal_32341 ;
    wire new_AGEMA_signal_32342 ;
    wire new_AGEMA_signal_32343 ;
    wire new_AGEMA_signal_32344 ;
    wire new_AGEMA_signal_32345 ;
    wire new_AGEMA_signal_32346 ;
    wire new_AGEMA_signal_32347 ;
    wire new_AGEMA_signal_32348 ;
    wire new_AGEMA_signal_32349 ;
    wire new_AGEMA_signal_32350 ;
    wire new_AGEMA_signal_32351 ;
    wire new_AGEMA_signal_32352 ;
    wire new_AGEMA_signal_32353 ;
    wire new_AGEMA_signal_32354 ;
    wire new_AGEMA_signal_32355 ;
    wire new_AGEMA_signal_32356 ;
    wire new_AGEMA_signal_32357 ;
    wire new_AGEMA_signal_32358 ;
    wire new_AGEMA_signal_32359 ;
    wire new_AGEMA_signal_32360 ;
    wire new_AGEMA_signal_32361 ;
    wire new_AGEMA_signal_32362 ;
    wire new_AGEMA_signal_32363 ;
    wire new_AGEMA_signal_32364 ;
    wire new_AGEMA_signal_32365 ;
    wire new_AGEMA_signal_32366 ;
    wire new_AGEMA_signal_32367 ;
    wire new_AGEMA_signal_32368 ;
    wire new_AGEMA_signal_32369 ;
    wire new_AGEMA_signal_32370 ;
    wire new_AGEMA_signal_32371 ;
    wire new_AGEMA_signal_32372 ;
    wire new_AGEMA_signal_32373 ;
    wire new_AGEMA_signal_32374 ;
    wire new_AGEMA_signal_32375 ;
    wire new_AGEMA_signal_32376 ;
    wire new_AGEMA_signal_32377 ;
    wire new_AGEMA_signal_32378 ;
    wire new_AGEMA_signal_32379 ;
    wire new_AGEMA_signal_32380 ;
    wire new_AGEMA_signal_32381 ;
    wire new_AGEMA_signal_32382 ;
    wire new_AGEMA_signal_32383 ;
    wire new_AGEMA_signal_32384 ;
    wire new_AGEMA_signal_32385 ;
    wire new_AGEMA_signal_32386 ;
    wire new_AGEMA_signal_32387 ;
    wire new_AGEMA_signal_32388 ;
    wire new_AGEMA_signal_32389 ;
    wire new_AGEMA_signal_32390 ;
    wire new_AGEMA_signal_32391 ;
    wire new_AGEMA_signal_32392 ;
    wire new_AGEMA_signal_32393 ;
    wire new_AGEMA_signal_32394 ;
    wire new_AGEMA_signal_32395 ;
    wire new_AGEMA_signal_32396 ;
    wire new_AGEMA_signal_32397 ;
    wire new_AGEMA_signal_32398 ;
    wire new_AGEMA_signal_32399 ;
    wire new_AGEMA_signal_32400 ;
    wire new_AGEMA_signal_32401 ;
    wire new_AGEMA_signal_32402 ;
    wire new_AGEMA_signal_32403 ;
    wire new_AGEMA_signal_32404 ;
    wire new_AGEMA_signal_32405 ;
    wire new_AGEMA_signal_32406 ;
    wire new_AGEMA_signal_32407 ;
    wire new_AGEMA_signal_32408 ;
    wire new_AGEMA_signal_32409 ;
    wire new_AGEMA_signal_32410 ;
    wire new_AGEMA_signal_32411 ;
    wire new_AGEMA_signal_32412 ;
    wire new_AGEMA_signal_32413 ;
    wire new_AGEMA_signal_32414 ;
    wire new_AGEMA_signal_32415 ;
    wire new_AGEMA_signal_32416 ;
    wire new_AGEMA_signal_32417 ;
    wire new_AGEMA_signal_32418 ;
    wire new_AGEMA_signal_32419 ;
    wire new_AGEMA_signal_32420 ;
    wire new_AGEMA_signal_32421 ;
    wire new_AGEMA_signal_32422 ;
    wire new_AGEMA_signal_32423 ;
    wire new_AGEMA_signal_32424 ;
    wire new_AGEMA_signal_32425 ;
    wire new_AGEMA_signal_32426 ;
    wire new_AGEMA_signal_32427 ;
    wire new_AGEMA_signal_32428 ;
    wire new_AGEMA_signal_32429 ;
    wire new_AGEMA_signal_32430 ;
    wire new_AGEMA_signal_32431 ;
    wire new_AGEMA_signal_32432 ;
    wire new_AGEMA_signal_32433 ;
    wire new_AGEMA_signal_32434 ;
    wire new_AGEMA_signal_32435 ;
    wire new_AGEMA_signal_32436 ;
    wire new_AGEMA_signal_32437 ;
    wire new_AGEMA_signal_32438 ;
    wire new_AGEMA_signal_32439 ;
    wire new_AGEMA_signal_32440 ;
    wire new_AGEMA_signal_32441 ;
    wire new_AGEMA_signal_32442 ;
    wire new_AGEMA_signal_32443 ;
    wire new_AGEMA_signal_32444 ;
    wire new_AGEMA_signal_32445 ;
    wire new_AGEMA_signal_32446 ;
    wire new_AGEMA_signal_32447 ;
    wire new_AGEMA_signal_32448 ;
    wire new_AGEMA_signal_32449 ;
    wire new_AGEMA_signal_32450 ;
    wire new_AGEMA_signal_32451 ;
    wire new_AGEMA_signal_32452 ;
    wire new_AGEMA_signal_32453 ;
    wire new_AGEMA_signal_32454 ;
    wire new_AGEMA_signal_32455 ;
    wire new_AGEMA_signal_32456 ;
    wire new_AGEMA_signal_32457 ;
    wire new_AGEMA_signal_32458 ;
    wire new_AGEMA_signal_32459 ;
    wire new_AGEMA_signal_32460 ;
    wire new_AGEMA_signal_32461 ;
    wire new_AGEMA_signal_32462 ;
    wire new_AGEMA_signal_32463 ;
    wire new_AGEMA_signal_32464 ;
    wire new_AGEMA_signal_32465 ;
    wire new_AGEMA_signal_32466 ;
    wire new_AGEMA_signal_32467 ;
    wire new_AGEMA_signal_32468 ;
    wire new_AGEMA_signal_32469 ;
    wire new_AGEMA_signal_32470 ;
    wire new_AGEMA_signal_32471 ;
    wire new_AGEMA_signal_32472 ;
    wire new_AGEMA_signal_32473 ;
    wire new_AGEMA_signal_32474 ;
    wire new_AGEMA_signal_32475 ;
    wire new_AGEMA_signal_32476 ;
    wire new_AGEMA_signal_32477 ;
    wire new_AGEMA_signal_32478 ;
    wire new_AGEMA_signal_32479 ;
    wire new_AGEMA_signal_32480 ;
    wire new_AGEMA_signal_32481 ;
    wire new_AGEMA_signal_32482 ;
    wire new_AGEMA_signal_32483 ;
    wire new_AGEMA_signal_32484 ;
    wire new_AGEMA_signal_32485 ;
    wire new_AGEMA_signal_32486 ;
    wire new_AGEMA_signal_32487 ;
    wire new_AGEMA_signal_32488 ;
    wire new_AGEMA_signal_32489 ;
    wire new_AGEMA_signal_32490 ;
    wire new_AGEMA_signal_32491 ;
    wire new_AGEMA_signal_32492 ;
    wire new_AGEMA_signal_32493 ;
    wire new_AGEMA_signal_32494 ;
    wire new_AGEMA_signal_32495 ;
    wire new_AGEMA_signal_32496 ;
    wire new_AGEMA_signal_32497 ;
    wire new_AGEMA_signal_32498 ;
    wire new_AGEMA_signal_32499 ;
    wire new_AGEMA_signal_32500 ;
    wire new_AGEMA_signal_32501 ;
    wire new_AGEMA_signal_32502 ;
    wire new_AGEMA_signal_32503 ;
    wire new_AGEMA_signal_32504 ;
    wire new_AGEMA_signal_32505 ;
    wire new_AGEMA_signal_32506 ;
    wire new_AGEMA_signal_32507 ;
    wire new_AGEMA_signal_32508 ;
    wire new_AGEMA_signal_32509 ;
    wire new_AGEMA_signal_32510 ;
    wire new_AGEMA_signal_32511 ;
    wire new_AGEMA_signal_32512 ;
    wire new_AGEMA_signal_32513 ;
    wire new_AGEMA_signal_32514 ;
    wire new_AGEMA_signal_32515 ;
    wire new_AGEMA_signal_32516 ;
    wire new_AGEMA_signal_32517 ;
    wire new_AGEMA_signal_32518 ;
    wire new_AGEMA_signal_32519 ;
    wire new_AGEMA_signal_32520 ;
    wire new_AGEMA_signal_32521 ;
    wire new_AGEMA_signal_32522 ;
    wire new_AGEMA_signal_32523 ;
    wire new_AGEMA_signal_32524 ;
    wire new_AGEMA_signal_32525 ;
    wire new_AGEMA_signal_32526 ;
    wire new_AGEMA_signal_32527 ;
    wire new_AGEMA_signal_32528 ;
    wire new_AGEMA_signal_32529 ;
    wire new_AGEMA_signal_32530 ;
    wire new_AGEMA_signal_32531 ;
    wire new_AGEMA_signal_32532 ;
    wire new_AGEMA_signal_32533 ;
    wire new_AGEMA_signal_32534 ;
    wire new_AGEMA_signal_32535 ;
    wire new_AGEMA_signal_32536 ;
    wire new_AGEMA_signal_32537 ;
    wire new_AGEMA_signal_32538 ;
    wire new_AGEMA_signal_32539 ;
    wire new_AGEMA_signal_32540 ;
    wire new_AGEMA_signal_32541 ;
    wire new_AGEMA_signal_32542 ;
    wire new_AGEMA_signal_32543 ;
    wire new_AGEMA_signal_32544 ;
    wire new_AGEMA_signal_32545 ;
    wire new_AGEMA_signal_32546 ;
    wire new_AGEMA_signal_32547 ;
    wire new_AGEMA_signal_32548 ;
    wire new_AGEMA_signal_32549 ;
    wire new_AGEMA_signal_32550 ;
    wire new_AGEMA_signal_32551 ;
    wire new_AGEMA_signal_32552 ;
    wire new_AGEMA_signal_32553 ;
    wire new_AGEMA_signal_32554 ;
    wire new_AGEMA_signal_32555 ;
    wire new_AGEMA_signal_32556 ;
    wire new_AGEMA_signal_32557 ;
    wire new_AGEMA_signal_32558 ;
    wire new_AGEMA_signal_32559 ;
    wire new_AGEMA_signal_32560 ;
    wire new_AGEMA_signal_32561 ;
    wire new_AGEMA_signal_32562 ;
    wire new_AGEMA_signal_32563 ;
    wire new_AGEMA_signal_32564 ;
    wire new_AGEMA_signal_32565 ;
    wire new_AGEMA_signal_32566 ;
    wire new_AGEMA_signal_32567 ;
    wire new_AGEMA_signal_32568 ;
    wire new_AGEMA_signal_32569 ;
    wire new_AGEMA_signal_32570 ;
    wire new_AGEMA_signal_32571 ;
    wire new_AGEMA_signal_32572 ;
    wire new_AGEMA_signal_32573 ;
    wire new_AGEMA_signal_32574 ;
    wire new_AGEMA_signal_32575 ;
    wire new_AGEMA_signal_32576 ;
    wire new_AGEMA_signal_32577 ;
    wire new_AGEMA_signal_32578 ;
    wire new_AGEMA_signal_32579 ;
    wire new_AGEMA_signal_32580 ;
    wire new_AGEMA_signal_32581 ;
    wire new_AGEMA_signal_32582 ;
    wire new_AGEMA_signal_32583 ;
    wire new_AGEMA_signal_32584 ;
    wire new_AGEMA_signal_32585 ;
    wire new_AGEMA_signal_32586 ;
    wire new_AGEMA_signal_32587 ;
    wire new_AGEMA_signal_32588 ;
    wire new_AGEMA_signal_32589 ;
    wire new_AGEMA_signal_32590 ;
    wire new_AGEMA_signal_32591 ;
    wire new_AGEMA_signal_32592 ;
    wire new_AGEMA_signal_32593 ;
    wire new_AGEMA_signal_32594 ;
    wire new_AGEMA_signal_32595 ;
    wire new_AGEMA_signal_32596 ;
    wire new_AGEMA_signal_32597 ;
    wire new_AGEMA_signal_32598 ;
    wire new_AGEMA_signal_32599 ;
    wire new_AGEMA_signal_32600 ;
    wire new_AGEMA_signal_32601 ;
    wire new_AGEMA_signal_32602 ;
    wire new_AGEMA_signal_32603 ;
    wire new_AGEMA_signal_32604 ;
    wire new_AGEMA_signal_32605 ;
    wire new_AGEMA_signal_32606 ;
    wire new_AGEMA_signal_32607 ;
    wire new_AGEMA_signal_32608 ;
    wire new_AGEMA_signal_32609 ;
    wire new_AGEMA_signal_32610 ;
    wire new_AGEMA_signal_32611 ;
    wire new_AGEMA_signal_32612 ;
    wire new_AGEMA_signal_32613 ;
    wire new_AGEMA_signal_32614 ;
    wire new_AGEMA_signal_32615 ;
    wire new_AGEMA_signal_32616 ;
    wire new_AGEMA_signal_32617 ;
    wire new_AGEMA_signal_32618 ;
    wire new_AGEMA_signal_32619 ;
    wire new_AGEMA_signal_32620 ;
    wire new_AGEMA_signal_32621 ;
    wire new_AGEMA_signal_32622 ;
    wire new_AGEMA_signal_32623 ;
    wire new_AGEMA_signal_32624 ;
    wire new_AGEMA_signal_32625 ;
    wire new_AGEMA_signal_32626 ;
    wire new_AGEMA_signal_32627 ;
    wire new_AGEMA_signal_32628 ;
    wire new_AGEMA_signal_32629 ;
    wire new_AGEMA_signal_32630 ;
    wire new_AGEMA_signal_32631 ;
    wire new_AGEMA_signal_32632 ;
    wire new_AGEMA_signal_32633 ;
    wire new_AGEMA_signal_32634 ;
    wire new_AGEMA_signal_32635 ;
    wire new_AGEMA_signal_32636 ;
    wire new_AGEMA_signal_32637 ;
    wire new_AGEMA_signal_32638 ;
    wire new_AGEMA_signal_32639 ;
    wire new_AGEMA_signal_32640 ;
    wire new_AGEMA_signal_32641 ;
    wire new_AGEMA_signal_32642 ;
    wire new_AGEMA_signal_32643 ;
    wire new_AGEMA_signal_32644 ;
    wire new_AGEMA_signal_32645 ;
    wire new_AGEMA_signal_32646 ;
    wire new_AGEMA_signal_32647 ;
    wire new_AGEMA_signal_32648 ;
    wire new_AGEMA_signal_32649 ;
    wire new_AGEMA_signal_32650 ;
    wire new_AGEMA_signal_32651 ;
    wire new_AGEMA_signal_32652 ;
    wire new_AGEMA_signal_32653 ;
    wire new_AGEMA_signal_32654 ;
    wire new_AGEMA_signal_32655 ;
    wire new_AGEMA_signal_32656 ;
    wire new_AGEMA_signal_32657 ;
    wire new_AGEMA_signal_32658 ;
    wire new_AGEMA_signal_32659 ;
    wire new_AGEMA_signal_32660 ;
    wire new_AGEMA_signal_32661 ;
    wire new_AGEMA_signal_32662 ;
    wire new_AGEMA_signal_32663 ;
    wire new_AGEMA_signal_32664 ;
    wire new_AGEMA_signal_32665 ;
    wire new_AGEMA_signal_32666 ;
    wire new_AGEMA_signal_32667 ;
    wire new_AGEMA_signal_32668 ;
    wire new_AGEMA_signal_32669 ;
    wire new_AGEMA_signal_32670 ;
    wire new_AGEMA_signal_32671 ;
    wire new_AGEMA_signal_32672 ;
    wire new_AGEMA_signal_32673 ;
    wire new_AGEMA_signal_32674 ;
    wire new_AGEMA_signal_32675 ;
    wire new_AGEMA_signal_32676 ;
    wire new_AGEMA_signal_32677 ;
    wire new_AGEMA_signal_32678 ;
    wire new_AGEMA_signal_32679 ;
    wire new_AGEMA_signal_32680 ;
    wire new_AGEMA_signal_32681 ;
    wire new_AGEMA_signal_32682 ;
    wire new_AGEMA_signal_32683 ;
    wire new_AGEMA_signal_32684 ;
    wire new_AGEMA_signal_32685 ;
    wire new_AGEMA_signal_32686 ;
    wire new_AGEMA_signal_32687 ;
    wire new_AGEMA_signal_32688 ;
    wire new_AGEMA_signal_32689 ;
    wire new_AGEMA_signal_32690 ;
    wire new_AGEMA_signal_32691 ;
    wire new_AGEMA_signal_32692 ;
    wire new_AGEMA_signal_32693 ;
    wire new_AGEMA_signal_32694 ;
    wire new_AGEMA_signal_32695 ;
    wire new_AGEMA_signal_32696 ;
    wire new_AGEMA_signal_32697 ;
    wire new_AGEMA_signal_32698 ;
    wire new_AGEMA_signal_32699 ;
    wire new_AGEMA_signal_32700 ;
    wire new_AGEMA_signal_32701 ;
    wire new_AGEMA_signal_32702 ;
    wire new_AGEMA_signal_32703 ;
    wire new_AGEMA_signal_32704 ;
    wire new_AGEMA_signal_32705 ;
    wire new_AGEMA_signal_32706 ;
    wire new_AGEMA_signal_32707 ;
    wire new_AGEMA_signal_32708 ;
    wire new_AGEMA_signal_32709 ;
    wire new_AGEMA_signal_32710 ;
    wire new_AGEMA_signal_32711 ;
    wire new_AGEMA_signal_32712 ;
    wire new_AGEMA_signal_32713 ;
    wire new_AGEMA_signal_32714 ;
    wire new_AGEMA_signal_32715 ;
    wire new_AGEMA_signal_32716 ;
    wire new_AGEMA_signal_32717 ;
    wire new_AGEMA_signal_32718 ;
    wire new_AGEMA_signal_32719 ;
    wire new_AGEMA_signal_32720 ;
    wire new_AGEMA_signal_32721 ;
    wire new_AGEMA_signal_32722 ;
    wire new_AGEMA_signal_32723 ;
    wire new_AGEMA_signal_32724 ;
    wire new_AGEMA_signal_32725 ;
    wire new_AGEMA_signal_32726 ;
    wire new_AGEMA_signal_32727 ;
    wire new_AGEMA_signal_32728 ;
    wire new_AGEMA_signal_32729 ;
    wire new_AGEMA_signal_32730 ;
    wire new_AGEMA_signal_32731 ;
    wire new_AGEMA_signal_32732 ;
    wire new_AGEMA_signal_32733 ;
    wire new_AGEMA_signal_32734 ;
    wire new_AGEMA_signal_32735 ;
    wire new_AGEMA_signal_32736 ;
    wire new_AGEMA_signal_32737 ;
    wire new_AGEMA_signal_32738 ;
    wire new_AGEMA_signal_32739 ;
    wire new_AGEMA_signal_32740 ;
    wire new_AGEMA_signal_32741 ;
    wire new_AGEMA_signal_32742 ;
    wire new_AGEMA_signal_32743 ;
    wire new_AGEMA_signal_32744 ;
    wire new_AGEMA_signal_32745 ;
    wire new_AGEMA_signal_32746 ;
    wire new_AGEMA_signal_32747 ;
    wire new_AGEMA_signal_32748 ;
    wire new_AGEMA_signal_32749 ;
    wire new_AGEMA_signal_32750 ;
    wire new_AGEMA_signal_32751 ;
    wire new_AGEMA_signal_32752 ;
    wire new_AGEMA_signal_32753 ;
    wire new_AGEMA_signal_32754 ;
    wire new_AGEMA_signal_32755 ;
    wire new_AGEMA_signal_32756 ;
    wire new_AGEMA_signal_32757 ;
    wire new_AGEMA_signal_32758 ;
    wire new_AGEMA_signal_32759 ;
    wire new_AGEMA_signal_32760 ;
    wire new_AGEMA_signal_32761 ;
    wire new_AGEMA_signal_32762 ;
    wire new_AGEMA_signal_32763 ;
    wire new_AGEMA_signal_32764 ;
    wire new_AGEMA_signal_32765 ;
    wire new_AGEMA_signal_32766 ;
    wire new_AGEMA_signal_32767 ;
    wire new_AGEMA_signal_32768 ;
    wire new_AGEMA_signal_32769 ;
    wire new_AGEMA_signal_32770 ;
    wire new_AGEMA_signal_32771 ;
    wire new_AGEMA_signal_32772 ;
    wire new_AGEMA_signal_32773 ;
    wire new_AGEMA_signal_32774 ;
    wire new_AGEMA_signal_32775 ;
    wire new_AGEMA_signal_32776 ;
    wire new_AGEMA_signal_32777 ;
    wire new_AGEMA_signal_32778 ;
    wire new_AGEMA_signal_32779 ;
    wire new_AGEMA_signal_32780 ;
    wire new_AGEMA_signal_32781 ;
    wire new_AGEMA_signal_32782 ;
    wire new_AGEMA_signal_32783 ;
    wire new_AGEMA_signal_32784 ;
    wire new_AGEMA_signal_32785 ;
    wire new_AGEMA_signal_32786 ;
    wire new_AGEMA_signal_32787 ;
    wire new_AGEMA_signal_32788 ;
    wire new_AGEMA_signal_32789 ;
    wire new_AGEMA_signal_32790 ;
    wire new_AGEMA_signal_32791 ;
    wire new_AGEMA_signal_32792 ;
    wire new_AGEMA_signal_32793 ;
    wire new_AGEMA_signal_32794 ;
    wire new_AGEMA_signal_32795 ;
    wire new_AGEMA_signal_32796 ;
    wire new_AGEMA_signal_32797 ;
    wire new_AGEMA_signal_32798 ;
    wire new_AGEMA_signal_32799 ;
    wire new_AGEMA_signal_32800 ;
    wire new_AGEMA_signal_32801 ;
    wire new_AGEMA_signal_32802 ;
    wire new_AGEMA_signal_32803 ;
    wire new_AGEMA_signal_32804 ;
    wire new_AGEMA_signal_32805 ;
    wire new_AGEMA_signal_32806 ;
    wire new_AGEMA_signal_32807 ;
    wire new_AGEMA_signal_32808 ;
    wire new_AGEMA_signal_32809 ;
    wire new_AGEMA_signal_32810 ;
    wire new_AGEMA_signal_32811 ;
    wire new_AGEMA_signal_32812 ;
    wire new_AGEMA_signal_32813 ;
    wire new_AGEMA_signal_32814 ;
    wire new_AGEMA_signal_32815 ;
    wire new_AGEMA_signal_32816 ;
    wire new_AGEMA_signal_32817 ;
    wire new_AGEMA_signal_32818 ;
    wire new_AGEMA_signal_32819 ;
    wire new_AGEMA_signal_32820 ;
    wire new_AGEMA_signal_32821 ;
    wire new_AGEMA_signal_32822 ;
    wire new_AGEMA_signal_32823 ;
    wire new_AGEMA_signal_32824 ;
    wire new_AGEMA_signal_32825 ;
    wire new_AGEMA_signal_32826 ;
    wire new_AGEMA_signal_32827 ;
    wire new_AGEMA_signal_32828 ;
    wire new_AGEMA_signal_32829 ;
    wire new_AGEMA_signal_32830 ;
    wire new_AGEMA_signal_32831 ;
    wire new_AGEMA_signal_32832 ;
    wire new_AGEMA_signal_32833 ;
    wire new_AGEMA_signal_32834 ;
    wire new_AGEMA_signal_32835 ;
    wire new_AGEMA_signal_32836 ;
    wire new_AGEMA_signal_32837 ;
    wire new_AGEMA_signal_32838 ;
    wire new_AGEMA_signal_32839 ;
    wire new_AGEMA_signal_32840 ;
    wire new_AGEMA_signal_32841 ;
    wire new_AGEMA_signal_32842 ;
    wire new_AGEMA_signal_32843 ;
    wire new_AGEMA_signal_32844 ;
    wire new_AGEMA_signal_32845 ;
    wire new_AGEMA_signal_32846 ;
    wire new_AGEMA_signal_32847 ;
    wire new_AGEMA_signal_32848 ;
    wire new_AGEMA_signal_32849 ;
    wire new_AGEMA_signal_32850 ;
    wire new_AGEMA_signal_32851 ;
    wire new_AGEMA_signal_32852 ;
    wire new_AGEMA_signal_32853 ;
    wire new_AGEMA_signal_32854 ;
    wire new_AGEMA_signal_32855 ;
    wire new_AGEMA_signal_32856 ;
    wire new_AGEMA_signal_32857 ;
    wire new_AGEMA_signal_32858 ;
    wire new_AGEMA_signal_32859 ;
    wire new_AGEMA_signal_32860 ;
    wire new_AGEMA_signal_32861 ;
    wire new_AGEMA_signal_32862 ;
    wire new_AGEMA_signal_32863 ;
    wire new_AGEMA_signal_32864 ;
    wire new_AGEMA_signal_32865 ;
    wire new_AGEMA_signal_32866 ;
    wire new_AGEMA_signal_32867 ;
    wire new_AGEMA_signal_32868 ;
    wire new_AGEMA_signal_32869 ;
    wire new_AGEMA_signal_32870 ;
    wire new_AGEMA_signal_32871 ;
    wire new_AGEMA_signal_32872 ;
    wire new_AGEMA_signal_32873 ;
    wire new_AGEMA_signal_32874 ;
    wire new_AGEMA_signal_32875 ;
    wire new_AGEMA_signal_32876 ;
    wire new_AGEMA_signal_32877 ;
    wire new_AGEMA_signal_32878 ;
    wire new_AGEMA_signal_32879 ;
    wire new_AGEMA_signal_32880 ;
    wire new_AGEMA_signal_32881 ;
    wire new_AGEMA_signal_32882 ;
    wire new_AGEMA_signal_32883 ;
    wire new_AGEMA_signal_32884 ;
    wire new_AGEMA_signal_32885 ;
    wire new_AGEMA_signal_32886 ;
    wire new_AGEMA_signal_32887 ;
    wire new_AGEMA_signal_32888 ;
    wire new_AGEMA_signal_32889 ;
    wire new_AGEMA_signal_32890 ;
    wire new_AGEMA_signal_32891 ;
    wire new_AGEMA_signal_32892 ;
    wire new_AGEMA_signal_32893 ;
    wire new_AGEMA_signal_32894 ;
    wire new_AGEMA_signal_32895 ;
    wire new_AGEMA_signal_32896 ;
    wire new_AGEMA_signal_32897 ;
    wire new_AGEMA_signal_32898 ;
    wire new_AGEMA_signal_32899 ;
    wire new_AGEMA_signal_32900 ;
    wire new_AGEMA_signal_32901 ;
    wire new_AGEMA_signal_32902 ;
    wire new_AGEMA_signal_32903 ;
    wire new_AGEMA_signal_32904 ;
    wire new_AGEMA_signal_32905 ;
    wire new_AGEMA_signal_32906 ;
    wire new_AGEMA_signal_32907 ;
    wire new_AGEMA_signal_32908 ;
    wire new_AGEMA_signal_32909 ;
    wire new_AGEMA_signal_32910 ;
    wire new_AGEMA_signal_32911 ;
    wire new_AGEMA_signal_32912 ;
    wire new_AGEMA_signal_32913 ;
    wire new_AGEMA_signal_32914 ;
    wire new_AGEMA_signal_32915 ;
    wire new_AGEMA_signal_32916 ;
    wire new_AGEMA_signal_32917 ;
    wire new_AGEMA_signal_32918 ;
    wire new_AGEMA_signal_32919 ;
    wire new_AGEMA_signal_32920 ;
    wire new_AGEMA_signal_32921 ;
    wire new_AGEMA_signal_32922 ;
    wire new_AGEMA_signal_32923 ;
    wire new_AGEMA_signal_32924 ;
    wire new_AGEMA_signal_32925 ;
    wire new_AGEMA_signal_32926 ;
    wire new_AGEMA_signal_32927 ;
    wire new_AGEMA_signal_32928 ;
    wire new_AGEMA_signal_32929 ;
    wire new_AGEMA_signal_32930 ;
    wire new_AGEMA_signal_32931 ;
    wire new_AGEMA_signal_32932 ;
    wire new_AGEMA_signal_32933 ;
    wire new_AGEMA_signal_32934 ;
    wire new_AGEMA_signal_32935 ;
    wire new_AGEMA_signal_32936 ;
    wire new_AGEMA_signal_32937 ;
    wire new_AGEMA_signal_32938 ;
    wire new_AGEMA_signal_32939 ;
    wire new_AGEMA_signal_32940 ;
    wire new_AGEMA_signal_32941 ;
    wire new_AGEMA_signal_32942 ;
    wire new_AGEMA_signal_32943 ;
    wire new_AGEMA_signal_32944 ;
    wire new_AGEMA_signal_32945 ;
    wire new_AGEMA_signal_32946 ;
    wire new_AGEMA_signal_32947 ;
    wire new_AGEMA_signal_32948 ;
    wire new_AGEMA_signal_32949 ;
    wire new_AGEMA_signal_32950 ;
    wire new_AGEMA_signal_32951 ;
    wire new_AGEMA_signal_32952 ;
    wire new_AGEMA_signal_32953 ;
    wire new_AGEMA_signal_32954 ;
    wire new_AGEMA_signal_32955 ;
    wire new_AGEMA_signal_32956 ;
    wire new_AGEMA_signal_32957 ;
    wire new_AGEMA_signal_32958 ;
    wire new_AGEMA_signal_32959 ;
    wire new_AGEMA_signal_32960 ;
    wire new_AGEMA_signal_32961 ;
    wire new_AGEMA_signal_32962 ;
    wire new_AGEMA_signal_32963 ;
    wire new_AGEMA_signal_32964 ;
    wire new_AGEMA_signal_32965 ;
    wire new_AGEMA_signal_32966 ;
    wire new_AGEMA_signal_32967 ;
    wire new_AGEMA_signal_32968 ;
    wire new_AGEMA_signal_32969 ;
    wire new_AGEMA_signal_32970 ;
    wire new_AGEMA_signal_32971 ;
    wire new_AGEMA_signal_32972 ;
    wire new_AGEMA_signal_32973 ;
    wire new_AGEMA_signal_32974 ;
    wire new_AGEMA_signal_32975 ;
    wire new_AGEMA_signal_32976 ;
    wire new_AGEMA_signal_32977 ;
    wire new_AGEMA_signal_32978 ;
    wire new_AGEMA_signal_32979 ;
    wire new_AGEMA_signal_32980 ;
    wire new_AGEMA_signal_32981 ;
    wire new_AGEMA_signal_32982 ;
    wire new_AGEMA_signal_32983 ;
    wire new_AGEMA_signal_32984 ;
    wire new_AGEMA_signal_32985 ;
    wire new_AGEMA_signal_32986 ;
    wire new_AGEMA_signal_32987 ;
    wire new_AGEMA_signal_32988 ;
    wire new_AGEMA_signal_32989 ;
    wire new_AGEMA_signal_32990 ;
    wire new_AGEMA_signal_32991 ;
    wire new_AGEMA_signal_32992 ;
    wire new_AGEMA_signal_32993 ;
    wire new_AGEMA_signal_32994 ;
    wire new_AGEMA_signal_32995 ;
    wire new_AGEMA_signal_32996 ;
    wire new_AGEMA_signal_32997 ;
    wire new_AGEMA_signal_32998 ;
    wire new_AGEMA_signal_32999 ;
    wire new_AGEMA_signal_33000 ;
    wire new_AGEMA_signal_33001 ;
    wire new_AGEMA_signal_33002 ;
    wire new_AGEMA_signal_33003 ;
    wire new_AGEMA_signal_33004 ;
    wire new_AGEMA_signal_33005 ;
    wire new_AGEMA_signal_33006 ;
    wire new_AGEMA_signal_33007 ;
    wire new_AGEMA_signal_33008 ;
    wire new_AGEMA_signal_33009 ;
    wire new_AGEMA_signal_33010 ;
    wire new_AGEMA_signal_33011 ;
    wire new_AGEMA_signal_33012 ;
    wire new_AGEMA_signal_33013 ;
    wire new_AGEMA_signal_33014 ;
    wire new_AGEMA_signal_33015 ;
    wire new_AGEMA_signal_33016 ;
    wire new_AGEMA_signal_33017 ;
    wire new_AGEMA_signal_33018 ;
    wire new_AGEMA_signal_33019 ;
    wire new_AGEMA_signal_33020 ;
    wire new_AGEMA_signal_33021 ;
    wire new_AGEMA_signal_33022 ;
    wire new_AGEMA_signal_33023 ;
    wire new_AGEMA_signal_33024 ;
    wire new_AGEMA_signal_33025 ;
    wire new_AGEMA_signal_33026 ;
    wire new_AGEMA_signal_33027 ;
    wire new_AGEMA_signal_33028 ;
    wire new_AGEMA_signal_33029 ;
    wire new_AGEMA_signal_33030 ;
    wire new_AGEMA_signal_33031 ;
    wire new_AGEMA_signal_33032 ;
    wire new_AGEMA_signal_33033 ;
    wire new_AGEMA_signal_33034 ;
    wire new_AGEMA_signal_33035 ;
    wire new_AGEMA_signal_33036 ;
    wire new_AGEMA_signal_33037 ;
    wire new_AGEMA_signal_33038 ;
    wire new_AGEMA_signal_33039 ;
    wire new_AGEMA_signal_33040 ;
    wire new_AGEMA_signal_33041 ;
    wire new_AGEMA_signal_33042 ;
    wire new_AGEMA_signal_33043 ;
    wire new_AGEMA_signal_33044 ;
    wire new_AGEMA_signal_33045 ;
    wire new_AGEMA_signal_33046 ;
    wire new_AGEMA_signal_33047 ;
    wire new_AGEMA_signal_33048 ;
    wire new_AGEMA_signal_33049 ;
    wire new_AGEMA_signal_33050 ;
    wire new_AGEMA_signal_33051 ;
    wire new_AGEMA_signal_33052 ;
    wire new_AGEMA_signal_33053 ;
    wire new_AGEMA_signal_33054 ;
    wire new_AGEMA_signal_33055 ;
    wire new_AGEMA_signal_33056 ;
    wire new_AGEMA_signal_33057 ;
    wire new_AGEMA_signal_33058 ;
    wire new_AGEMA_signal_33059 ;
    wire new_AGEMA_signal_33060 ;
    wire new_AGEMA_signal_33061 ;
    wire new_AGEMA_signal_33062 ;
    wire new_AGEMA_signal_33063 ;
    wire new_AGEMA_signal_33064 ;
    wire new_AGEMA_signal_33065 ;
    wire new_AGEMA_signal_33066 ;
    wire new_AGEMA_signal_33067 ;
    wire new_AGEMA_signal_33068 ;
    wire new_AGEMA_signal_33069 ;
    wire new_AGEMA_signal_33070 ;
    wire new_AGEMA_signal_33071 ;
    wire new_AGEMA_signal_33072 ;
    wire new_AGEMA_signal_33073 ;
    wire new_AGEMA_signal_33074 ;
    wire new_AGEMA_signal_33075 ;
    wire new_AGEMA_signal_33076 ;
    wire new_AGEMA_signal_33077 ;
    wire new_AGEMA_signal_33078 ;
    wire new_AGEMA_signal_33079 ;
    wire new_AGEMA_signal_33080 ;
    wire new_AGEMA_signal_33081 ;
    wire new_AGEMA_signal_33082 ;
    wire new_AGEMA_signal_33083 ;
    wire new_AGEMA_signal_33084 ;
    wire new_AGEMA_signal_33085 ;
    wire new_AGEMA_signal_33086 ;
    wire new_AGEMA_signal_33087 ;
    wire new_AGEMA_signal_33088 ;
    wire new_AGEMA_signal_33089 ;
    wire new_AGEMA_signal_33090 ;
    wire new_AGEMA_signal_33091 ;
    wire new_AGEMA_signal_33092 ;
    wire new_AGEMA_signal_33093 ;
    wire new_AGEMA_signal_33094 ;
    wire new_AGEMA_signal_33095 ;
    wire new_AGEMA_signal_33096 ;
    wire new_AGEMA_signal_33097 ;
    wire new_AGEMA_signal_33098 ;
    wire new_AGEMA_signal_33099 ;
    wire new_AGEMA_signal_33100 ;
    wire new_AGEMA_signal_33101 ;
    wire new_AGEMA_signal_33102 ;
    wire new_AGEMA_signal_33103 ;
    wire new_AGEMA_signal_33104 ;
    wire new_AGEMA_signal_33105 ;
    wire new_AGEMA_signal_33106 ;
    wire new_AGEMA_signal_33107 ;
    wire new_AGEMA_signal_33108 ;
    wire new_AGEMA_signal_33109 ;
    wire new_AGEMA_signal_33110 ;
    wire new_AGEMA_signal_33111 ;
    wire new_AGEMA_signal_33112 ;
    wire new_AGEMA_signal_33113 ;
    wire new_AGEMA_signal_33114 ;
    wire new_AGEMA_signal_33115 ;
    wire new_AGEMA_signal_33116 ;
    wire new_AGEMA_signal_33117 ;
    wire new_AGEMA_signal_33118 ;
    wire new_AGEMA_signal_33119 ;
    wire new_AGEMA_signal_33120 ;
    wire new_AGEMA_signal_33121 ;
    wire new_AGEMA_signal_33122 ;
    wire new_AGEMA_signal_33123 ;
    wire new_AGEMA_signal_33124 ;
    wire new_AGEMA_signal_33125 ;
    wire new_AGEMA_signal_33126 ;
    wire new_AGEMA_signal_33127 ;
    wire new_AGEMA_signal_33128 ;
    wire new_AGEMA_signal_33129 ;
    wire new_AGEMA_signal_33130 ;
    wire new_AGEMA_signal_33131 ;
    wire new_AGEMA_signal_33132 ;
    wire new_AGEMA_signal_33133 ;
    wire new_AGEMA_signal_33134 ;
    wire new_AGEMA_signal_33135 ;
    wire new_AGEMA_signal_33136 ;
    wire new_AGEMA_signal_33137 ;
    wire new_AGEMA_signal_33138 ;
    wire new_AGEMA_signal_33139 ;
    wire new_AGEMA_signal_33140 ;
    wire new_AGEMA_signal_33141 ;
    wire new_AGEMA_signal_33142 ;
    wire new_AGEMA_signal_33143 ;
    wire new_AGEMA_signal_33144 ;
    wire new_AGEMA_signal_33145 ;
    wire new_AGEMA_signal_33146 ;
    wire new_AGEMA_signal_33147 ;
    wire new_AGEMA_signal_33148 ;
    wire new_AGEMA_signal_33149 ;
    wire new_AGEMA_signal_33150 ;
    wire new_AGEMA_signal_33151 ;
    wire new_AGEMA_signal_33152 ;
    wire new_AGEMA_signal_33153 ;
    wire new_AGEMA_signal_33154 ;
    wire new_AGEMA_signal_33155 ;
    wire new_AGEMA_signal_33156 ;
    wire new_AGEMA_signal_33157 ;
    wire new_AGEMA_signal_33158 ;
    wire new_AGEMA_signal_33159 ;
    wire new_AGEMA_signal_33160 ;
    wire new_AGEMA_signal_33161 ;
    wire new_AGEMA_signal_33162 ;
    wire new_AGEMA_signal_33163 ;
    wire new_AGEMA_signal_33164 ;
    wire new_AGEMA_signal_33165 ;
    wire new_AGEMA_signal_33166 ;
    wire new_AGEMA_signal_33167 ;
    wire new_AGEMA_signal_33168 ;
    wire new_AGEMA_signal_33169 ;
    wire new_AGEMA_signal_33170 ;
    wire new_AGEMA_signal_33171 ;
    wire new_AGEMA_signal_33172 ;
    wire new_AGEMA_signal_33173 ;
    wire new_AGEMA_signal_33174 ;
    wire new_AGEMA_signal_33175 ;
    wire new_AGEMA_signal_33176 ;
    wire new_AGEMA_signal_33177 ;
    wire new_AGEMA_signal_33178 ;
    wire new_AGEMA_signal_33179 ;
    wire new_AGEMA_signal_33180 ;
    wire new_AGEMA_signal_33181 ;
    wire new_AGEMA_signal_33182 ;
    wire new_AGEMA_signal_33183 ;
    wire new_AGEMA_signal_33184 ;
    wire new_AGEMA_signal_33185 ;
    wire new_AGEMA_signal_33186 ;
    wire new_AGEMA_signal_33187 ;
    wire new_AGEMA_signal_33188 ;
    wire new_AGEMA_signal_33189 ;
    wire new_AGEMA_signal_33190 ;
    wire new_AGEMA_signal_33191 ;
    wire new_AGEMA_signal_33192 ;
    wire new_AGEMA_signal_33193 ;
    wire new_AGEMA_signal_33194 ;
    wire new_AGEMA_signal_33195 ;
    wire new_AGEMA_signal_33196 ;
    wire new_AGEMA_signal_33197 ;
    wire new_AGEMA_signal_33198 ;
    wire new_AGEMA_signal_33199 ;
    wire new_AGEMA_signal_33200 ;
    wire new_AGEMA_signal_33201 ;
    wire new_AGEMA_signal_33202 ;
    wire new_AGEMA_signal_33203 ;
    wire new_AGEMA_signal_33204 ;
    wire new_AGEMA_signal_33205 ;
    wire new_AGEMA_signal_33206 ;
    wire new_AGEMA_signal_33207 ;
    wire new_AGEMA_signal_33208 ;
    wire new_AGEMA_signal_33209 ;
    wire new_AGEMA_signal_33210 ;
    wire new_AGEMA_signal_33211 ;
    wire new_AGEMA_signal_33212 ;
    wire new_AGEMA_signal_33213 ;
    wire new_AGEMA_signal_33214 ;
    wire new_AGEMA_signal_33215 ;
    wire new_AGEMA_signal_33216 ;
    wire new_AGEMA_signal_33217 ;
    wire new_AGEMA_signal_33218 ;
    wire new_AGEMA_signal_33219 ;
    wire new_AGEMA_signal_33220 ;
    wire new_AGEMA_signal_33221 ;
    wire new_AGEMA_signal_33222 ;
    wire new_AGEMA_signal_33223 ;
    wire new_AGEMA_signal_33224 ;
    wire new_AGEMA_signal_33225 ;
    wire new_AGEMA_signal_33226 ;
    wire new_AGEMA_signal_33227 ;
    wire new_AGEMA_signal_33228 ;
    wire new_AGEMA_signal_33229 ;
    wire new_AGEMA_signal_33230 ;
    wire new_AGEMA_signal_33231 ;
    wire new_AGEMA_signal_33232 ;
    wire new_AGEMA_signal_33233 ;
    wire new_AGEMA_signal_33234 ;
    wire new_AGEMA_signal_33235 ;
    wire new_AGEMA_signal_33236 ;
    wire new_AGEMA_signal_33237 ;
    wire new_AGEMA_signal_33238 ;
    wire new_AGEMA_signal_33239 ;
    wire new_AGEMA_signal_33240 ;
    wire new_AGEMA_signal_33241 ;
    wire new_AGEMA_signal_33242 ;
    wire new_AGEMA_signal_33243 ;
    wire new_AGEMA_signal_33244 ;
    wire new_AGEMA_signal_33245 ;
    wire new_AGEMA_signal_33246 ;
    wire new_AGEMA_signal_33247 ;
    wire new_AGEMA_signal_33248 ;
    wire new_AGEMA_signal_33249 ;
    wire new_AGEMA_signal_33250 ;
    wire new_AGEMA_signal_33251 ;
    wire new_AGEMA_signal_33252 ;
    wire new_AGEMA_signal_33253 ;
    wire new_AGEMA_signal_33254 ;
    wire new_AGEMA_signal_33255 ;
    wire new_AGEMA_signal_33256 ;
    wire new_AGEMA_signal_33257 ;
    wire new_AGEMA_signal_33258 ;
    wire new_AGEMA_signal_33259 ;
    wire new_AGEMA_signal_33260 ;
    wire new_AGEMA_signal_33261 ;
    wire new_AGEMA_signal_33262 ;
    wire new_AGEMA_signal_33263 ;
    wire new_AGEMA_signal_33264 ;
    wire new_AGEMA_signal_33265 ;
    wire new_AGEMA_signal_33266 ;
    wire new_AGEMA_signal_33267 ;
    wire new_AGEMA_signal_33268 ;
    wire new_AGEMA_signal_33269 ;
    wire new_AGEMA_signal_33270 ;
    wire new_AGEMA_signal_33271 ;
    wire new_AGEMA_signal_33272 ;
    wire new_AGEMA_signal_33273 ;
    wire new_AGEMA_signal_33274 ;
    wire new_AGEMA_signal_33275 ;
    wire new_AGEMA_signal_33276 ;
    wire new_AGEMA_signal_33277 ;
    wire new_AGEMA_signal_33278 ;
    wire new_AGEMA_signal_33279 ;
    wire new_AGEMA_signal_33280 ;
    wire new_AGEMA_signal_33281 ;
    wire new_AGEMA_signal_33282 ;
    wire new_AGEMA_signal_33283 ;
    wire new_AGEMA_signal_33284 ;
    wire new_AGEMA_signal_33285 ;
    wire new_AGEMA_signal_33286 ;
    wire new_AGEMA_signal_33287 ;
    wire new_AGEMA_signal_33288 ;
    wire new_AGEMA_signal_33289 ;
    wire new_AGEMA_signal_33290 ;
    wire new_AGEMA_signal_33291 ;
    wire new_AGEMA_signal_33292 ;
    wire new_AGEMA_signal_33293 ;
    wire new_AGEMA_signal_33294 ;
    wire new_AGEMA_signal_33295 ;
    wire new_AGEMA_signal_33296 ;
    wire new_AGEMA_signal_33297 ;
    wire new_AGEMA_signal_33298 ;
    wire new_AGEMA_signal_33299 ;
    wire new_AGEMA_signal_33300 ;
    wire new_AGEMA_signal_33301 ;
    wire new_AGEMA_signal_33302 ;
    wire new_AGEMA_signal_33303 ;
    wire new_AGEMA_signal_33304 ;
    wire new_AGEMA_signal_33305 ;
    wire new_AGEMA_signal_33306 ;
    wire new_AGEMA_signal_33307 ;
    wire new_AGEMA_signal_33308 ;
    wire new_AGEMA_signal_33309 ;
    wire new_AGEMA_signal_33310 ;
    wire new_AGEMA_signal_33311 ;
    wire new_AGEMA_signal_33312 ;
    wire new_AGEMA_signal_33313 ;
    wire new_AGEMA_signal_33314 ;
    wire new_AGEMA_signal_33315 ;
    wire new_AGEMA_signal_33316 ;
    wire new_AGEMA_signal_33317 ;
    wire new_AGEMA_signal_33318 ;
    wire new_AGEMA_signal_33319 ;
    wire new_AGEMA_signal_33320 ;
    wire new_AGEMA_signal_33321 ;
    wire new_AGEMA_signal_33322 ;
    wire new_AGEMA_signal_33323 ;
    wire new_AGEMA_signal_33324 ;
    wire new_AGEMA_signal_33325 ;
    wire new_AGEMA_signal_33326 ;
    wire new_AGEMA_signal_33327 ;
    wire new_AGEMA_signal_33328 ;
    wire new_AGEMA_signal_33329 ;
    wire new_AGEMA_signal_33330 ;
    wire new_AGEMA_signal_33331 ;
    wire new_AGEMA_signal_33332 ;
    wire new_AGEMA_signal_33333 ;
    wire new_AGEMA_signal_33334 ;
    wire new_AGEMA_signal_33335 ;
    wire new_AGEMA_signal_33336 ;
    wire new_AGEMA_signal_33337 ;
    wire new_AGEMA_signal_33338 ;
    wire new_AGEMA_signal_33339 ;
    wire new_AGEMA_signal_33340 ;
    wire new_AGEMA_signal_33341 ;
    wire new_AGEMA_signal_33342 ;
    wire new_AGEMA_signal_33343 ;
    wire new_AGEMA_signal_33344 ;
    wire new_AGEMA_signal_33345 ;
    wire new_AGEMA_signal_33346 ;
    wire new_AGEMA_signal_33347 ;
    wire new_AGEMA_signal_33348 ;
    wire new_AGEMA_signal_33349 ;
    wire new_AGEMA_signal_33350 ;
    wire new_AGEMA_signal_33351 ;
    wire new_AGEMA_signal_33352 ;
    wire new_AGEMA_signal_33353 ;
    wire new_AGEMA_signal_33354 ;
    wire new_AGEMA_signal_33355 ;
    wire new_AGEMA_signal_33356 ;
    wire new_AGEMA_signal_33357 ;
    wire new_AGEMA_signal_33358 ;
    wire new_AGEMA_signal_33359 ;
    wire new_AGEMA_signal_33360 ;
    wire new_AGEMA_signal_33361 ;
    wire new_AGEMA_signal_33362 ;
    wire new_AGEMA_signal_33363 ;
    wire new_AGEMA_signal_33364 ;
    wire new_AGEMA_signal_33365 ;
    wire new_AGEMA_signal_33366 ;
    wire new_AGEMA_signal_33367 ;
    wire new_AGEMA_signal_33368 ;
    wire new_AGEMA_signal_33369 ;
    wire new_AGEMA_signal_33370 ;
    wire new_AGEMA_signal_33371 ;
    wire new_AGEMA_signal_33372 ;
    wire new_AGEMA_signal_33373 ;
    wire new_AGEMA_signal_33374 ;
    wire new_AGEMA_signal_33375 ;
    wire new_AGEMA_signal_33376 ;
    wire new_AGEMA_signal_33377 ;
    wire new_AGEMA_signal_33378 ;
    wire new_AGEMA_signal_33379 ;
    wire new_AGEMA_signal_33380 ;
    wire new_AGEMA_signal_33381 ;
    wire new_AGEMA_signal_33382 ;
    wire new_AGEMA_signal_33383 ;
    wire new_AGEMA_signal_33384 ;
    wire new_AGEMA_signal_33385 ;
    wire new_AGEMA_signal_33386 ;
    wire new_AGEMA_signal_33387 ;
    wire new_AGEMA_signal_33388 ;
    wire new_AGEMA_signal_33389 ;
    wire new_AGEMA_signal_33390 ;
    wire new_AGEMA_signal_33391 ;
    wire new_AGEMA_signal_33392 ;
    wire new_AGEMA_signal_33393 ;
    wire new_AGEMA_signal_33394 ;
    wire new_AGEMA_signal_33395 ;
    wire new_AGEMA_signal_33396 ;
    wire new_AGEMA_signal_33397 ;
    wire new_AGEMA_signal_33398 ;
    wire new_AGEMA_signal_33399 ;
    wire new_AGEMA_signal_33400 ;
    wire new_AGEMA_signal_33401 ;
    wire new_AGEMA_signal_33402 ;
    wire new_AGEMA_signal_33403 ;
    wire new_AGEMA_signal_33404 ;
    wire new_AGEMA_signal_33405 ;
    wire new_AGEMA_signal_33406 ;
    wire new_AGEMA_signal_33407 ;
    wire new_AGEMA_signal_33408 ;
    wire new_AGEMA_signal_33409 ;
    wire new_AGEMA_signal_33410 ;
    wire new_AGEMA_signal_33411 ;
    wire new_AGEMA_signal_33412 ;
    wire new_AGEMA_signal_33413 ;
    wire new_AGEMA_signal_33414 ;
    wire new_AGEMA_signal_33415 ;
    wire new_AGEMA_signal_33416 ;
    wire new_AGEMA_signal_33417 ;
    wire new_AGEMA_signal_33418 ;
    wire new_AGEMA_signal_33419 ;
    wire new_AGEMA_signal_33420 ;
    wire new_AGEMA_signal_33421 ;
    wire new_AGEMA_signal_33422 ;
    wire new_AGEMA_signal_33423 ;
    wire new_AGEMA_signal_33424 ;
    wire new_AGEMA_signal_33425 ;
    wire new_AGEMA_signal_33426 ;
    wire new_AGEMA_signal_33427 ;
    wire new_AGEMA_signal_33428 ;
    wire new_AGEMA_signal_33429 ;
    wire new_AGEMA_signal_33430 ;
    wire new_AGEMA_signal_33431 ;
    wire new_AGEMA_signal_33432 ;
    wire new_AGEMA_signal_33433 ;
    wire new_AGEMA_signal_33434 ;
    wire new_AGEMA_signal_33435 ;
    wire new_AGEMA_signal_33436 ;
    wire new_AGEMA_signal_33437 ;
    wire new_AGEMA_signal_33438 ;
    wire new_AGEMA_signal_33439 ;
    wire new_AGEMA_signal_33440 ;
    wire new_AGEMA_signal_33441 ;
    wire new_AGEMA_signal_33442 ;
    wire new_AGEMA_signal_33443 ;
    wire new_AGEMA_signal_33444 ;
    wire new_AGEMA_signal_33445 ;
    wire new_AGEMA_signal_33446 ;
    wire new_AGEMA_signal_33447 ;
    wire new_AGEMA_signal_33448 ;
    wire new_AGEMA_signal_33449 ;
    wire new_AGEMA_signal_33450 ;
    wire new_AGEMA_signal_33451 ;
    wire new_AGEMA_signal_33452 ;
    wire new_AGEMA_signal_33453 ;
    wire new_AGEMA_signal_33454 ;
    wire new_AGEMA_signal_33455 ;
    wire new_AGEMA_signal_33456 ;
    wire new_AGEMA_signal_33457 ;
    wire new_AGEMA_signal_33458 ;
    wire new_AGEMA_signal_33459 ;
    wire new_AGEMA_signal_33460 ;
    wire new_AGEMA_signal_33461 ;
    wire new_AGEMA_signal_33462 ;
    wire new_AGEMA_signal_33463 ;
    wire new_AGEMA_signal_33464 ;
    wire new_AGEMA_signal_33465 ;
    wire new_AGEMA_signal_33466 ;
    wire new_AGEMA_signal_33467 ;
    wire new_AGEMA_signal_33468 ;
    wire new_AGEMA_signal_33469 ;
    wire new_AGEMA_signal_33470 ;
    wire new_AGEMA_signal_33471 ;
    wire new_AGEMA_signal_33472 ;
    wire new_AGEMA_signal_33473 ;
    wire new_AGEMA_signal_33474 ;
    wire new_AGEMA_signal_33475 ;
    wire new_AGEMA_signal_33476 ;
    wire new_AGEMA_signal_33477 ;
    wire new_AGEMA_signal_33478 ;
    wire new_AGEMA_signal_33479 ;
    wire new_AGEMA_signal_33480 ;
    wire new_AGEMA_signal_33481 ;
    wire new_AGEMA_signal_33482 ;
    wire new_AGEMA_signal_33483 ;
    wire new_AGEMA_signal_33484 ;
    wire new_AGEMA_signal_33485 ;
    wire new_AGEMA_signal_33486 ;
    wire new_AGEMA_signal_33487 ;
    wire new_AGEMA_signal_33488 ;
    wire new_AGEMA_signal_33489 ;
    wire new_AGEMA_signal_33490 ;
    wire new_AGEMA_signal_33491 ;
    wire new_AGEMA_signal_33492 ;
    wire new_AGEMA_signal_33493 ;
    wire new_AGEMA_signal_33494 ;
    wire new_AGEMA_signal_33495 ;
    wire new_AGEMA_signal_33496 ;
    wire new_AGEMA_signal_33497 ;
    wire new_AGEMA_signal_33498 ;
    wire new_AGEMA_signal_33499 ;
    wire new_AGEMA_signal_33500 ;
    wire new_AGEMA_signal_33501 ;
    wire new_AGEMA_signal_33502 ;
    wire new_AGEMA_signal_33503 ;
    wire new_AGEMA_signal_33504 ;
    wire new_AGEMA_signal_33505 ;
    wire new_AGEMA_signal_33506 ;
    wire new_AGEMA_signal_33507 ;
    wire new_AGEMA_signal_33508 ;
    wire new_AGEMA_signal_33509 ;
    wire new_AGEMA_signal_33510 ;
    wire new_AGEMA_signal_33511 ;
    wire new_AGEMA_signal_33512 ;
    wire new_AGEMA_signal_33513 ;
    wire new_AGEMA_signal_33514 ;
    wire new_AGEMA_signal_33515 ;
    wire new_AGEMA_signal_33516 ;
    wire new_AGEMA_signal_33517 ;
    wire new_AGEMA_signal_33518 ;
    wire new_AGEMA_signal_33519 ;
    wire new_AGEMA_signal_33520 ;
    wire new_AGEMA_signal_33521 ;
    wire new_AGEMA_signal_33522 ;
    wire new_AGEMA_signal_33523 ;
    wire new_AGEMA_signal_33524 ;
    wire new_AGEMA_signal_33525 ;
    wire new_AGEMA_signal_33526 ;
    wire new_AGEMA_signal_33527 ;
    wire new_AGEMA_signal_33528 ;
    wire new_AGEMA_signal_33529 ;
    wire new_AGEMA_signal_33530 ;
    wire new_AGEMA_signal_33531 ;
    wire new_AGEMA_signal_33532 ;
    wire new_AGEMA_signal_33533 ;
    wire new_AGEMA_signal_33534 ;
    wire new_AGEMA_signal_33535 ;
    wire new_AGEMA_signal_33536 ;
    wire new_AGEMA_signal_33537 ;
    wire new_AGEMA_signal_33538 ;
    wire new_AGEMA_signal_33539 ;
    wire new_AGEMA_signal_33540 ;
    wire new_AGEMA_signal_33541 ;
    wire new_AGEMA_signal_33542 ;
    wire new_AGEMA_signal_33543 ;
    wire new_AGEMA_signal_33544 ;
    wire new_AGEMA_signal_33545 ;
    wire new_AGEMA_signal_33546 ;
    wire new_AGEMA_signal_33547 ;
    wire new_AGEMA_signal_33548 ;
    wire new_AGEMA_signal_33549 ;
    wire new_AGEMA_signal_33550 ;
    wire new_AGEMA_signal_33551 ;
    wire new_AGEMA_signal_33552 ;
    wire new_AGEMA_signal_33553 ;
    wire new_AGEMA_signal_33554 ;
    wire new_AGEMA_signal_33555 ;
    wire new_AGEMA_signal_33556 ;
    wire new_AGEMA_signal_33557 ;
    wire new_AGEMA_signal_33558 ;
    wire new_AGEMA_signal_33559 ;
    wire new_AGEMA_signal_33560 ;
    wire new_AGEMA_signal_33561 ;
    wire new_AGEMA_signal_33562 ;
    wire new_AGEMA_signal_33563 ;
    wire new_AGEMA_signal_33564 ;
    wire new_AGEMA_signal_33565 ;
    wire new_AGEMA_signal_33566 ;
    wire new_AGEMA_signal_33567 ;
    wire new_AGEMA_signal_33568 ;
    wire new_AGEMA_signal_33569 ;
    wire new_AGEMA_signal_33570 ;
    wire new_AGEMA_signal_33571 ;
    wire new_AGEMA_signal_33572 ;
    wire new_AGEMA_signal_33573 ;
    wire new_AGEMA_signal_33574 ;
    wire new_AGEMA_signal_33575 ;
    wire new_AGEMA_signal_33576 ;
    wire new_AGEMA_signal_33577 ;
    wire new_AGEMA_signal_33578 ;
    wire new_AGEMA_signal_33579 ;
    wire new_AGEMA_signal_33580 ;
    wire new_AGEMA_signal_33581 ;
    wire new_AGEMA_signal_33582 ;
    wire new_AGEMA_signal_33583 ;
    wire new_AGEMA_signal_33584 ;
    wire new_AGEMA_signal_33585 ;
    wire new_AGEMA_signal_33586 ;
    wire new_AGEMA_signal_33587 ;
    wire new_AGEMA_signal_33588 ;
    wire new_AGEMA_signal_33589 ;
    wire new_AGEMA_signal_33590 ;
    wire new_AGEMA_signal_33591 ;
    wire new_AGEMA_signal_33592 ;
    wire new_AGEMA_signal_33593 ;
    wire new_AGEMA_signal_33594 ;
    wire new_AGEMA_signal_33595 ;
    wire new_AGEMA_signal_33596 ;
    wire new_AGEMA_signal_33597 ;
    wire new_AGEMA_signal_33598 ;
    wire new_AGEMA_signal_33599 ;
    wire new_AGEMA_signal_33600 ;
    wire new_AGEMA_signal_33601 ;
    wire new_AGEMA_signal_33602 ;
    wire new_AGEMA_signal_33603 ;
    wire new_AGEMA_signal_33604 ;
    wire new_AGEMA_signal_33605 ;
    wire new_AGEMA_signal_33606 ;
    wire new_AGEMA_signal_33607 ;
    wire new_AGEMA_signal_33608 ;
    wire new_AGEMA_signal_33609 ;
    wire new_AGEMA_signal_33610 ;
    wire new_AGEMA_signal_33611 ;
    wire new_AGEMA_signal_33612 ;
    wire new_AGEMA_signal_33613 ;
    wire new_AGEMA_signal_33614 ;
    wire new_AGEMA_signal_33615 ;
    wire new_AGEMA_signal_33616 ;
    wire new_AGEMA_signal_33617 ;
    wire new_AGEMA_signal_33618 ;
    wire new_AGEMA_signal_33619 ;
    wire new_AGEMA_signal_33620 ;
    wire new_AGEMA_signal_33621 ;
    wire new_AGEMA_signal_33622 ;
    wire new_AGEMA_signal_33623 ;
    wire new_AGEMA_signal_33624 ;
    wire new_AGEMA_signal_33625 ;
    wire new_AGEMA_signal_33626 ;
    wire new_AGEMA_signal_33627 ;
    wire new_AGEMA_signal_33628 ;
    wire new_AGEMA_signal_33629 ;
    wire new_AGEMA_signal_33630 ;
    wire new_AGEMA_signal_33631 ;
    wire new_AGEMA_signal_33632 ;
    wire new_AGEMA_signal_33633 ;
    wire new_AGEMA_signal_33634 ;
    wire new_AGEMA_signal_33635 ;
    wire new_AGEMA_signal_33636 ;
    wire new_AGEMA_signal_33637 ;
    wire new_AGEMA_signal_33638 ;
    wire new_AGEMA_signal_33639 ;
    wire new_AGEMA_signal_33640 ;
    wire new_AGEMA_signal_33641 ;
    wire new_AGEMA_signal_33642 ;
    wire new_AGEMA_signal_33643 ;
    wire new_AGEMA_signal_33644 ;
    wire new_AGEMA_signal_33645 ;
    wire new_AGEMA_signal_33646 ;
    wire new_AGEMA_signal_33647 ;
    wire new_AGEMA_signal_33648 ;
    wire new_AGEMA_signal_33649 ;
    wire new_AGEMA_signal_33650 ;
    wire new_AGEMA_signal_33651 ;
    wire new_AGEMA_signal_33652 ;
    wire new_AGEMA_signal_33653 ;
    wire new_AGEMA_signal_33654 ;
    wire new_AGEMA_signal_33655 ;
    wire new_AGEMA_signal_33656 ;
    wire new_AGEMA_signal_33657 ;
    wire new_AGEMA_signal_33658 ;
    wire new_AGEMA_signal_33659 ;
    wire new_AGEMA_signal_33660 ;
    wire new_AGEMA_signal_33661 ;
    wire new_AGEMA_signal_33662 ;
    wire new_AGEMA_signal_33663 ;
    wire new_AGEMA_signal_33664 ;
    wire new_AGEMA_signal_33665 ;
    wire new_AGEMA_signal_33666 ;
    wire new_AGEMA_signal_33667 ;
    wire new_AGEMA_signal_33668 ;
    wire new_AGEMA_signal_33669 ;
    wire new_AGEMA_signal_33670 ;
    wire new_AGEMA_signal_33671 ;
    wire new_AGEMA_signal_33672 ;
    wire new_AGEMA_signal_33673 ;
    wire new_AGEMA_signal_33674 ;
    wire new_AGEMA_signal_33675 ;
    wire new_AGEMA_signal_33676 ;
    wire new_AGEMA_signal_33677 ;
    wire new_AGEMA_signal_33678 ;
    wire new_AGEMA_signal_33679 ;
    wire new_AGEMA_signal_33680 ;
    wire new_AGEMA_signal_33681 ;
    wire new_AGEMA_signal_33682 ;
    wire new_AGEMA_signal_33683 ;
    wire new_AGEMA_signal_33684 ;
    wire new_AGEMA_signal_33685 ;
    wire new_AGEMA_signal_33686 ;
    wire new_AGEMA_signal_33687 ;
    wire new_AGEMA_signal_33688 ;
    wire new_AGEMA_signal_33689 ;
    wire new_AGEMA_signal_33690 ;
    wire new_AGEMA_signal_33691 ;
    wire new_AGEMA_signal_33692 ;
    wire new_AGEMA_signal_33693 ;
    wire new_AGEMA_signal_33694 ;
    wire new_AGEMA_signal_33695 ;
    wire new_AGEMA_signal_33696 ;
    wire new_AGEMA_signal_33697 ;
    wire new_AGEMA_signal_33698 ;
    wire new_AGEMA_signal_33699 ;
    wire new_AGEMA_signal_33700 ;
    wire new_AGEMA_signal_33701 ;
    wire new_AGEMA_signal_33702 ;
    wire new_AGEMA_signal_33703 ;
    wire new_AGEMA_signal_33704 ;
    wire new_AGEMA_signal_33705 ;
    wire new_AGEMA_signal_33706 ;
    wire new_AGEMA_signal_33707 ;
    wire new_AGEMA_signal_33708 ;
    wire new_AGEMA_signal_33709 ;
    wire new_AGEMA_signal_33710 ;
    wire new_AGEMA_signal_33711 ;
    wire new_AGEMA_signal_33712 ;
    wire new_AGEMA_signal_33713 ;
    wire new_AGEMA_signal_33714 ;
    wire new_AGEMA_signal_33715 ;
    wire new_AGEMA_signal_33716 ;
    wire new_AGEMA_signal_33717 ;
    wire new_AGEMA_signal_33718 ;
    wire new_AGEMA_signal_33719 ;
    wire new_AGEMA_signal_33720 ;
    wire new_AGEMA_signal_33721 ;
    wire new_AGEMA_signal_33722 ;
    wire new_AGEMA_signal_33723 ;
    wire new_AGEMA_signal_33724 ;
    wire new_AGEMA_signal_33725 ;
    wire new_AGEMA_signal_33726 ;
    wire new_AGEMA_signal_33727 ;
    wire new_AGEMA_signal_33728 ;
    wire new_AGEMA_signal_33729 ;
    wire new_AGEMA_signal_33730 ;
    wire new_AGEMA_signal_33731 ;
    wire new_AGEMA_signal_33732 ;
    wire new_AGEMA_signal_33733 ;
    wire new_AGEMA_signal_33734 ;
    wire new_AGEMA_signal_33735 ;
    wire new_AGEMA_signal_33736 ;
    wire new_AGEMA_signal_33737 ;
    wire new_AGEMA_signal_33738 ;
    wire new_AGEMA_signal_33739 ;
    wire new_AGEMA_signal_33740 ;
    wire new_AGEMA_signal_33741 ;
    wire new_AGEMA_signal_33742 ;
    wire new_AGEMA_signal_33743 ;
    wire new_AGEMA_signal_33744 ;
    wire new_AGEMA_signal_33745 ;
    wire new_AGEMA_signal_33746 ;
    wire new_AGEMA_signal_33747 ;
    wire new_AGEMA_signal_33748 ;
    wire new_AGEMA_signal_33749 ;
    wire new_AGEMA_signal_33750 ;
    wire new_AGEMA_signal_33751 ;
    wire new_AGEMA_signal_33752 ;
    wire new_AGEMA_signal_33753 ;
    wire new_AGEMA_signal_33754 ;
    wire new_AGEMA_signal_33755 ;
    wire new_AGEMA_signal_33756 ;
    wire new_AGEMA_signal_33757 ;
    wire new_AGEMA_signal_33758 ;
    wire new_AGEMA_signal_33759 ;
    wire new_AGEMA_signal_33760 ;
    wire new_AGEMA_signal_33761 ;
    wire new_AGEMA_signal_33762 ;
    wire new_AGEMA_signal_33763 ;
    wire new_AGEMA_signal_33764 ;
    wire new_AGEMA_signal_33765 ;
    wire new_AGEMA_signal_33766 ;
    wire new_AGEMA_signal_33767 ;
    wire new_AGEMA_signal_33768 ;
    wire new_AGEMA_signal_33769 ;
    wire new_AGEMA_signal_33770 ;
    wire new_AGEMA_signal_33771 ;
    wire new_AGEMA_signal_33772 ;
    wire new_AGEMA_signal_33773 ;
    wire new_AGEMA_signal_33774 ;
    wire new_AGEMA_signal_33775 ;
    wire new_AGEMA_signal_33776 ;
    wire new_AGEMA_signal_33777 ;
    wire new_AGEMA_signal_33778 ;
    wire new_AGEMA_signal_33779 ;
    wire new_AGEMA_signal_33780 ;
    wire new_AGEMA_signal_33781 ;
    wire new_AGEMA_signal_33782 ;
    wire new_AGEMA_signal_33783 ;
    wire new_AGEMA_signal_33784 ;
    wire new_AGEMA_signal_33785 ;
    wire new_AGEMA_signal_33786 ;
    wire new_AGEMA_signal_33787 ;
    wire new_AGEMA_signal_33788 ;
    wire new_AGEMA_signal_33789 ;
    wire new_AGEMA_signal_33790 ;
    wire new_AGEMA_signal_33791 ;
    wire new_AGEMA_signal_33792 ;
    wire new_AGEMA_signal_33793 ;
    wire new_AGEMA_signal_33794 ;
    wire new_AGEMA_signal_33795 ;
    wire new_AGEMA_signal_33796 ;
    wire new_AGEMA_signal_33797 ;
    wire new_AGEMA_signal_33798 ;
    wire new_AGEMA_signal_33799 ;
    wire new_AGEMA_signal_33800 ;
    wire new_AGEMA_signal_33801 ;
    wire new_AGEMA_signal_33802 ;
    wire new_AGEMA_signal_33803 ;
    wire new_AGEMA_signal_33804 ;
    wire new_AGEMA_signal_33805 ;
    wire new_AGEMA_signal_33806 ;
    wire new_AGEMA_signal_33807 ;
    wire new_AGEMA_signal_33808 ;
    wire new_AGEMA_signal_33809 ;
    wire new_AGEMA_signal_33810 ;
    wire new_AGEMA_signal_33811 ;
    wire new_AGEMA_signal_33812 ;
    wire new_AGEMA_signal_33813 ;
    wire new_AGEMA_signal_33814 ;
    wire new_AGEMA_signal_33815 ;
    wire new_AGEMA_signal_33816 ;
    wire new_AGEMA_signal_33817 ;
    wire new_AGEMA_signal_33818 ;
    wire new_AGEMA_signal_33819 ;
    wire new_AGEMA_signal_33820 ;
    wire new_AGEMA_signal_33821 ;
    wire new_AGEMA_signal_33822 ;
    wire new_AGEMA_signal_33823 ;
    wire new_AGEMA_signal_33824 ;
    wire new_AGEMA_signal_33825 ;
    wire new_AGEMA_signal_33826 ;
    wire new_AGEMA_signal_33827 ;
    wire new_AGEMA_signal_33828 ;
    wire new_AGEMA_signal_33829 ;
    wire new_AGEMA_signal_33830 ;
    wire new_AGEMA_signal_33831 ;
    wire new_AGEMA_signal_33832 ;
    wire new_AGEMA_signal_33833 ;
    wire new_AGEMA_signal_33834 ;
    wire new_AGEMA_signal_33835 ;
    wire new_AGEMA_signal_33836 ;
    wire new_AGEMA_signal_33837 ;
    wire new_AGEMA_signal_33838 ;
    wire new_AGEMA_signal_33839 ;
    wire new_AGEMA_signal_33840 ;
    wire new_AGEMA_signal_33841 ;
    wire new_AGEMA_signal_33842 ;
    wire new_AGEMA_signal_33843 ;
    wire new_AGEMA_signal_33844 ;
    wire new_AGEMA_signal_33845 ;
    wire new_AGEMA_signal_33846 ;
    wire new_AGEMA_signal_33847 ;
    wire new_AGEMA_signal_33848 ;
    wire new_AGEMA_signal_33849 ;
    wire new_AGEMA_signal_33850 ;
    wire new_AGEMA_signal_33851 ;
    wire new_AGEMA_signal_33852 ;
    wire new_AGEMA_signal_33853 ;
    wire new_AGEMA_signal_33854 ;
    wire new_AGEMA_signal_33855 ;
    wire new_AGEMA_signal_33856 ;
    wire new_AGEMA_signal_33857 ;
    wire new_AGEMA_signal_33858 ;
    wire new_AGEMA_signal_33859 ;
    wire new_AGEMA_signal_33860 ;
    wire new_AGEMA_signal_33861 ;
    wire new_AGEMA_signal_33862 ;
    wire new_AGEMA_signal_33863 ;
    wire new_AGEMA_signal_33864 ;
    wire new_AGEMA_signal_33865 ;
    wire new_AGEMA_signal_33866 ;
    wire new_AGEMA_signal_33867 ;
    wire new_AGEMA_signal_33868 ;
    wire new_AGEMA_signal_33869 ;
    wire new_AGEMA_signal_33870 ;
    wire new_AGEMA_signal_33871 ;
    wire new_AGEMA_signal_33872 ;
    wire new_AGEMA_signal_33873 ;
    wire new_AGEMA_signal_33874 ;
    wire new_AGEMA_signal_33875 ;
    wire new_AGEMA_signal_33876 ;
    wire new_AGEMA_signal_33877 ;
    wire new_AGEMA_signal_33878 ;
    wire new_AGEMA_signal_33879 ;
    wire new_AGEMA_signal_33880 ;
    wire new_AGEMA_signal_33881 ;
    wire new_AGEMA_signal_33882 ;
    wire new_AGEMA_signal_33883 ;
    wire new_AGEMA_signal_33884 ;
    wire new_AGEMA_signal_33885 ;
    wire new_AGEMA_signal_33886 ;
    wire new_AGEMA_signal_33887 ;
    wire new_AGEMA_signal_33888 ;
    wire new_AGEMA_signal_33889 ;
    wire new_AGEMA_signal_33890 ;
    wire new_AGEMA_signal_33891 ;
    wire new_AGEMA_signal_33892 ;
    wire new_AGEMA_signal_33893 ;
    wire new_AGEMA_signal_33894 ;
    wire new_AGEMA_signal_33895 ;
    wire new_AGEMA_signal_33896 ;
    wire new_AGEMA_signal_33897 ;
    wire new_AGEMA_signal_33898 ;
    wire new_AGEMA_signal_33899 ;
    wire new_AGEMA_signal_33900 ;
    wire new_AGEMA_signal_33901 ;
    wire new_AGEMA_signal_33902 ;
    wire new_AGEMA_signal_33903 ;
    wire new_AGEMA_signal_33904 ;
    wire new_AGEMA_signal_33905 ;
    wire new_AGEMA_signal_33906 ;
    wire new_AGEMA_signal_33907 ;
    wire new_AGEMA_signal_33908 ;
    wire new_AGEMA_signal_33909 ;
    wire new_AGEMA_signal_33910 ;
    wire new_AGEMA_signal_33911 ;
    wire new_AGEMA_signal_33912 ;
    wire new_AGEMA_signal_33913 ;
    wire new_AGEMA_signal_33914 ;
    wire new_AGEMA_signal_33915 ;
    wire new_AGEMA_signal_33916 ;
    wire new_AGEMA_signal_33917 ;
    wire new_AGEMA_signal_33918 ;
    wire new_AGEMA_signal_33919 ;
    wire new_AGEMA_signal_33920 ;
    wire new_AGEMA_signal_33921 ;
    wire new_AGEMA_signal_33922 ;
    wire new_AGEMA_signal_33923 ;
    wire new_AGEMA_signal_33924 ;
    wire new_AGEMA_signal_33925 ;
    wire new_AGEMA_signal_33926 ;
    wire new_AGEMA_signal_33927 ;
    wire new_AGEMA_signal_33928 ;
    wire new_AGEMA_signal_33929 ;
    wire new_AGEMA_signal_33930 ;
    wire new_AGEMA_signal_33931 ;
    wire new_AGEMA_signal_33932 ;
    wire new_AGEMA_signal_33933 ;
    wire new_AGEMA_signal_33934 ;
    wire new_AGEMA_signal_33935 ;
    wire new_AGEMA_signal_33936 ;
    wire new_AGEMA_signal_33937 ;
    wire new_AGEMA_signal_33938 ;
    wire new_AGEMA_signal_33939 ;
    wire new_AGEMA_signal_33940 ;
    wire new_AGEMA_signal_33941 ;
    wire new_AGEMA_signal_33942 ;
    wire new_AGEMA_signal_33943 ;
    wire new_AGEMA_signal_33944 ;
    wire new_AGEMA_signal_33945 ;
    wire new_AGEMA_signal_33946 ;
    wire new_AGEMA_signal_33947 ;
    wire new_AGEMA_signal_33948 ;
    wire new_AGEMA_signal_33949 ;
    wire new_AGEMA_signal_33950 ;
    wire new_AGEMA_signal_33951 ;
    wire new_AGEMA_signal_33952 ;
    wire new_AGEMA_signal_33953 ;
    wire new_AGEMA_signal_33954 ;
    wire new_AGEMA_signal_33955 ;
    wire new_AGEMA_signal_33956 ;
    wire new_AGEMA_signal_33957 ;
    wire new_AGEMA_signal_33958 ;
    wire new_AGEMA_signal_33959 ;
    wire new_AGEMA_signal_33960 ;
    wire new_AGEMA_signal_33961 ;
    wire new_AGEMA_signal_33962 ;
    wire new_AGEMA_signal_33963 ;
    wire new_AGEMA_signal_33964 ;
    wire new_AGEMA_signal_33965 ;
    wire new_AGEMA_signal_33966 ;
    wire new_AGEMA_signal_33967 ;
    wire new_AGEMA_signal_33968 ;
    wire new_AGEMA_signal_33969 ;
    wire new_AGEMA_signal_33970 ;
    wire new_AGEMA_signal_33971 ;
    wire new_AGEMA_signal_33972 ;
    wire new_AGEMA_signal_33973 ;
    wire new_AGEMA_signal_33974 ;
    wire new_AGEMA_signal_33975 ;
    wire new_AGEMA_signal_33976 ;
    wire new_AGEMA_signal_33977 ;
    wire new_AGEMA_signal_33978 ;
    wire new_AGEMA_signal_33979 ;
    wire new_AGEMA_signal_33980 ;
    wire new_AGEMA_signal_33981 ;
    wire new_AGEMA_signal_33982 ;
    wire new_AGEMA_signal_33983 ;
    wire new_AGEMA_signal_33984 ;
    wire new_AGEMA_signal_33985 ;
    wire new_AGEMA_signal_33986 ;
    wire new_AGEMA_signal_33987 ;
    wire new_AGEMA_signal_33988 ;
    wire new_AGEMA_signal_33989 ;
    wire new_AGEMA_signal_33990 ;
    wire new_AGEMA_signal_33991 ;
    wire new_AGEMA_signal_33992 ;
    wire new_AGEMA_signal_33993 ;
    wire new_AGEMA_signal_33994 ;
    wire new_AGEMA_signal_33995 ;
    wire new_AGEMA_signal_33996 ;
    wire new_AGEMA_signal_33997 ;
    wire new_AGEMA_signal_33998 ;
    wire new_AGEMA_signal_33999 ;
    wire new_AGEMA_signal_34000 ;
    wire new_AGEMA_signal_34001 ;
    wire new_AGEMA_signal_34002 ;
    wire new_AGEMA_signal_34003 ;
    wire new_AGEMA_signal_34004 ;
    wire new_AGEMA_signal_34005 ;
    wire new_AGEMA_signal_34006 ;
    wire new_AGEMA_signal_34007 ;
    wire new_AGEMA_signal_34008 ;
    wire new_AGEMA_signal_34009 ;
    wire new_AGEMA_signal_34010 ;
    wire new_AGEMA_signal_34011 ;
    wire new_AGEMA_signal_34012 ;
    wire new_AGEMA_signal_34013 ;
    wire new_AGEMA_signal_34014 ;
    wire new_AGEMA_signal_34015 ;
    wire new_AGEMA_signal_34016 ;
    wire new_AGEMA_signal_34017 ;
    wire new_AGEMA_signal_34018 ;
    wire new_AGEMA_signal_34019 ;
    wire new_AGEMA_signal_34020 ;
    wire new_AGEMA_signal_34021 ;
    wire new_AGEMA_signal_34022 ;
    wire new_AGEMA_signal_34023 ;
    wire new_AGEMA_signal_34024 ;
    wire new_AGEMA_signal_34025 ;
    wire new_AGEMA_signal_34026 ;
    wire new_AGEMA_signal_34027 ;
    wire new_AGEMA_signal_34028 ;
    wire new_AGEMA_signal_34029 ;
    wire new_AGEMA_signal_34030 ;
    wire new_AGEMA_signal_34031 ;
    wire new_AGEMA_signal_34032 ;
    wire new_AGEMA_signal_34033 ;
    wire new_AGEMA_signal_34034 ;
    wire new_AGEMA_signal_34035 ;
    wire new_AGEMA_signal_34036 ;
    wire new_AGEMA_signal_34037 ;
    wire new_AGEMA_signal_34038 ;
    wire new_AGEMA_signal_34039 ;
    wire new_AGEMA_signal_34040 ;
    wire new_AGEMA_signal_34041 ;
    wire new_AGEMA_signal_34042 ;
    wire new_AGEMA_signal_34043 ;
    wire new_AGEMA_signal_34044 ;
    wire new_AGEMA_signal_34045 ;
    wire new_AGEMA_signal_34046 ;
    wire new_AGEMA_signal_34047 ;
    wire new_AGEMA_signal_34048 ;
    wire new_AGEMA_signal_34049 ;
    wire new_AGEMA_signal_34050 ;
    wire new_AGEMA_signal_34051 ;
    wire new_AGEMA_signal_34052 ;
    wire new_AGEMA_signal_34053 ;
    wire new_AGEMA_signal_34054 ;
    wire new_AGEMA_signal_34055 ;
    wire new_AGEMA_signal_34056 ;
    wire new_AGEMA_signal_34057 ;
    wire new_AGEMA_signal_34058 ;
    wire new_AGEMA_signal_34059 ;
    wire new_AGEMA_signal_34060 ;
    wire new_AGEMA_signal_34061 ;
    wire new_AGEMA_signal_34062 ;
    wire new_AGEMA_signal_34063 ;
    wire new_AGEMA_signal_34064 ;
    wire new_AGEMA_signal_34065 ;
    wire new_AGEMA_signal_34066 ;
    wire new_AGEMA_signal_34067 ;
    wire new_AGEMA_signal_34068 ;
    wire new_AGEMA_signal_34069 ;
    wire new_AGEMA_signal_34070 ;
    wire new_AGEMA_signal_34071 ;
    wire new_AGEMA_signal_34072 ;
    wire new_AGEMA_signal_34073 ;
    wire new_AGEMA_signal_34074 ;
    wire new_AGEMA_signal_34075 ;
    wire new_AGEMA_signal_34076 ;
    wire new_AGEMA_signal_34077 ;
    wire new_AGEMA_signal_34078 ;
    wire new_AGEMA_signal_34079 ;
    wire new_AGEMA_signal_34080 ;
    wire new_AGEMA_signal_34081 ;
    wire new_AGEMA_signal_34082 ;
    wire new_AGEMA_signal_34083 ;
    wire new_AGEMA_signal_34084 ;
    wire new_AGEMA_signal_34085 ;
    wire new_AGEMA_signal_34086 ;
    wire new_AGEMA_signal_34087 ;
    wire new_AGEMA_signal_34088 ;
    wire new_AGEMA_signal_34089 ;
    wire new_AGEMA_signal_34090 ;
    wire new_AGEMA_signal_34091 ;
    wire new_AGEMA_signal_34092 ;
    wire new_AGEMA_signal_34093 ;
    wire new_AGEMA_signal_34094 ;
    wire new_AGEMA_signal_34095 ;
    wire new_AGEMA_signal_34096 ;
    wire new_AGEMA_signal_34097 ;
    wire new_AGEMA_signal_34098 ;
    wire new_AGEMA_signal_34099 ;
    wire new_AGEMA_signal_34100 ;
    wire new_AGEMA_signal_34101 ;
    wire new_AGEMA_signal_34102 ;
    wire new_AGEMA_signal_34103 ;
    wire new_AGEMA_signal_34104 ;
    wire new_AGEMA_signal_34105 ;
    wire new_AGEMA_signal_34106 ;
    wire new_AGEMA_signal_34107 ;
    wire new_AGEMA_signal_34108 ;
    wire new_AGEMA_signal_34109 ;
    wire new_AGEMA_signal_34110 ;
    wire new_AGEMA_signal_34111 ;
    wire new_AGEMA_signal_34112 ;
    wire new_AGEMA_signal_34113 ;
    wire new_AGEMA_signal_34114 ;
    wire new_AGEMA_signal_34115 ;
    wire new_AGEMA_signal_34116 ;
    wire new_AGEMA_signal_34117 ;
    wire new_AGEMA_signal_34118 ;
    wire new_AGEMA_signal_34119 ;
    wire new_AGEMA_signal_34120 ;
    wire new_AGEMA_signal_34121 ;
    wire new_AGEMA_signal_34122 ;
    wire new_AGEMA_signal_34123 ;
    wire new_AGEMA_signal_34124 ;
    wire new_AGEMA_signal_34125 ;
    wire new_AGEMA_signal_34126 ;
    wire new_AGEMA_signal_34127 ;
    wire new_AGEMA_signal_34128 ;
    wire new_AGEMA_signal_34129 ;
    wire new_AGEMA_signal_34130 ;
    wire new_AGEMA_signal_34131 ;
    wire new_AGEMA_signal_34132 ;
    wire new_AGEMA_signal_34133 ;
    wire new_AGEMA_signal_34134 ;
    wire new_AGEMA_signal_34135 ;
    wire new_AGEMA_signal_34136 ;
    wire new_AGEMA_signal_34137 ;
    wire new_AGEMA_signal_34138 ;
    wire new_AGEMA_signal_34139 ;
    wire new_AGEMA_signal_34140 ;
    wire new_AGEMA_signal_34141 ;
    wire new_AGEMA_signal_34142 ;
    wire new_AGEMA_signal_34143 ;
    wire new_AGEMA_signal_34144 ;
    wire new_AGEMA_signal_34145 ;
    wire new_AGEMA_signal_34146 ;
    wire new_AGEMA_signal_34147 ;
    wire new_AGEMA_signal_34148 ;
    wire new_AGEMA_signal_34149 ;
    wire new_AGEMA_signal_34150 ;
    wire new_AGEMA_signal_34151 ;
    wire new_AGEMA_signal_34152 ;
    wire new_AGEMA_signal_34153 ;
    wire new_AGEMA_signal_34154 ;
    wire new_AGEMA_signal_34155 ;
    wire new_AGEMA_signal_34156 ;
    wire new_AGEMA_signal_34157 ;
    wire new_AGEMA_signal_34158 ;
    wire new_AGEMA_signal_34159 ;
    wire new_AGEMA_signal_34160 ;
    wire new_AGEMA_signal_34161 ;
    wire new_AGEMA_signal_34162 ;
    wire new_AGEMA_signal_34163 ;
    wire new_AGEMA_signal_34164 ;
    wire new_AGEMA_signal_34165 ;
    wire new_AGEMA_signal_34166 ;
    wire new_AGEMA_signal_34167 ;
    wire new_AGEMA_signal_34168 ;
    wire new_AGEMA_signal_34169 ;
    wire new_AGEMA_signal_34170 ;
    wire new_AGEMA_signal_34171 ;
    wire new_AGEMA_signal_34172 ;
    wire new_AGEMA_signal_34173 ;
    wire new_AGEMA_signal_34174 ;
    wire new_AGEMA_signal_34175 ;
    wire new_AGEMA_signal_34176 ;
    wire new_AGEMA_signal_34177 ;
    wire new_AGEMA_signal_34178 ;
    wire new_AGEMA_signal_34179 ;
    wire new_AGEMA_signal_34180 ;
    wire new_AGEMA_signal_34181 ;
    wire new_AGEMA_signal_34182 ;
    wire new_AGEMA_signal_34183 ;
    wire new_AGEMA_signal_34184 ;
    wire new_AGEMA_signal_34185 ;
    wire new_AGEMA_signal_34186 ;
    wire new_AGEMA_signal_34187 ;
    wire new_AGEMA_signal_34188 ;
    wire new_AGEMA_signal_34189 ;
    wire new_AGEMA_signal_34190 ;
    wire new_AGEMA_signal_34191 ;
    wire new_AGEMA_signal_34192 ;
    wire new_AGEMA_signal_34193 ;
    wire new_AGEMA_signal_34194 ;
    wire new_AGEMA_signal_34195 ;
    wire new_AGEMA_signal_34196 ;
    wire new_AGEMA_signal_34197 ;
    wire new_AGEMA_signal_34198 ;
    wire new_AGEMA_signal_34199 ;
    wire new_AGEMA_signal_34200 ;
    wire new_AGEMA_signal_34201 ;
    wire new_AGEMA_signal_34202 ;
    wire new_AGEMA_signal_34203 ;
    wire new_AGEMA_signal_34204 ;
    wire new_AGEMA_signal_34205 ;
    wire new_AGEMA_signal_34206 ;
    wire new_AGEMA_signal_34207 ;
    wire new_AGEMA_signal_34208 ;
    wire new_AGEMA_signal_34209 ;
    wire new_AGEMA_signal_34210 ;
    wire new_AGEMA_signal_34211 ;
    wire new_AGEMA_signal_34212 ;
    wire new_AGEMA_signal_34213 ;
    wire new_AGEMA_signal_34214 ;
    wire new_AGEMA_signal_34215 ;
    wire new_AGEMA_signal_34216 ;
    wire new_AGEMA_signal_34217 ;
    wire new_AGEMA_signal_34218 ;
    wire new_AGEMA_signal_34219 ;
    wire new_AGEMA_signal_34220 ;
    wire new_AGEMA_signal_34221 ;
    wire new_AGEMA_signal_34222 ;
    wire new_AGEMA_signal_34223 ;
    wire new_AGEMA_signal_34224 ;
    wire new_AGEMA_signal_34225 ;
    wire new_AGEMA_signal_34226 ;
    wire new_AGEMA_signal_34227 ;
    wire new_AGEMA_signal_34228 ;
    wire new_AGEMA_signal_34229 ;
    wire new_AGEMA_signal_34230 ;
    wire new_AGEMA_signal_34231 ;
    wire new_AGEMA_signal_34232 ;
    wire new_AGEMA_signal_34233 ;
    wire new_AGEMA_signal_34234 ;
    wire new_AGEMA_signal_34235 ;
    wire new_AGEMA_signal_34236 ;
    wire new_AGEMA_signal_34237 ;
    wire new_AGEMA_signal_34238 ;
    wire new_AGEMA_signal_34239 ;
    wire new_AGEMA_signal_34240 ;
    wire new_AGEMA_signal_34241 ;
    wire new_AGEMA_signal_34242 ;
    wire new_AGEMA_signal_34243 ;
    wire new_AGEMA_signal_34244 ;
    wire new_AGEMA_signal_34245 ;
    wire new_AGEMA_signal_34246 ;
    wire new_AGEMA_signal_34247 ;
    wire new_AGEMA_signal_34248 ;
    wire new_AGEMA_signal_34249 ;
    wire new_AGEMA_signal_34250 ;
    wire new_AGEMA_signal_34251 ;
    wire new_AGEMA_signal_34252 ;
    wire new_AGEMA_signal_34253 ;
    wire new_AGEMA_signal_34254 ;
    wire new_AGEMA_signal_34255 ;
    wire new_AGEMA_signal_34256 ;
    wire new_AGEMA_signal_34257 ;
    wire new_AGEMA_signal_34258 ;
    wire new_AGEMA_signal_34259 ;
    wire new_AGEMA_signal_34260 ;
    wire new_AGEMA_signal_34261 ;
    wire new_AGEMA_signal_34262 ;
    wire new_AGEMA_signal_34263 ;
    wire new_AGEMA_signal_34264 ;
    wire new_AGEMA_signal_34265 ;
    wire new_AGEMA_signal_34266 ;
    wire new_AGEMA_signal_34267 ;
    wire new_AGEMA_signal_34268 ;
    wire new_AGEMA_signal_34269 ;
    wire new_AGEMA_signal_34270 ;
    wire new_AGEMA_signal_34271 ;
    wire new_AGEMA_signal_34272 ;
    wire new_AGEMA_signal_34273 ;
    wire new_AGEMA_signal_34274 ;
    wire new_AGEMA_signal_34275 ;
    wire new_AGEMA_signal_34276 ;
    wire new_AGEMA_signal_34277 ;
    wire new_AGEMA_signal_34278 ;
    wire new_AGEMA_signal_34279 ;
    wire new_AGEMA_signal_34280 ;
    wire new_AGEMA_signal_34281 ;
    wire new_AGEMA_signal_34282 ;
    wire new_AGEMA_signal_34283 ;
    wire new_AGEMA_signal_34284 ;
    wire new_AGEMA_signal_34285 ;
    wire new_AGEMA_signal_34286 ;
    wire new_AGEMA_signal_34287 ;
    wire new_AGEMA_signal_34288 ;
    wire new_AGEMA_signal_34289 ;
    wire new_AGEMA_signal_34290 ;
    wire new_AGEMA_signal_34291 ;
    wire new_AGEMA_signal_34292 ;
    wire new_AGEMA_signal_34293 ;
    wire new_AGEMA_signal_34294 ;
    wire new_AGEMA_signal_34295 ;
    wire new_AGEMA_signal_34296 ;
    wire new_AGEMA_signal_34297 ;
    wire new_AGEMA_signal_34298 ;
    wire new_AGEMA_signal_34299 ;
    wire new_AGEMA_signal_34300 ;
    wire new_AGEMA_signal_34301 ;
    wire new_AGEMA_signal_34302 ;
    wire new_AGEMA_signal_34303 ;
    wire new_AGEMA_signal_34304 ;
    wire new_AGEMA_signal_34305 ;
    wire new_AGEMA_signal_34306 ;
    wire new_AGEMA_signal_34307 ;
    wire new_AGEMA_signal_34308 ;
    wire new_AGEMA_signal_34309 ;
    wire new_AGEMA_signal_34310 ;
    wire new_AGEMA_signal_34311 ;
    wire new_AGEMA_signal_34312 ;
    wire new_AGEMA_signal_34313 ;
    wire new_AGEMA_signal_34314 ;
    wire new_AGEMA_signal_34315 ;
    wire new_AGEMA_signal_34316 ;
    wire new_AGEMA_signal_34317 ;
    wire new_AGEMA_signal_34318 ;
    wire new_AGEMA_signal_34319 ;
    wire new_AGEMA_signal_34320 ;
    wire new_AGEMA_signal_34321 ;
    wire new_AGEMA_signal_34322 ;
    wire new_AGEMA_signal_34323 ;
    wire new_AGEMA_signal_34324 ;
    wire new_AGEMA_signal_34325 ;
    wire new_AGEMA_signal_34326 ;
    wire new_AGEMA_signal_34327 ;
    wire new_AGEMA_signal_34328 ;
    wire new_AGEMA_signal_34329 ;
    wire new_AGEMA_signal_34330 ;
    wire new_AGEMA_signal_34331 ;
    wire new_AGEMA_signal_34332 ;
    wire new_AGEMA_signal_34333 ;
    wire new_AGEMA_signal_34334 ;
    wire new_AGEMA_signal_34335 ;
    wire new_AGEMA_signal_34336 ;
    wire new_AGEMA_signal_34337 ;
    wire new_AGEMA_signal_34338 ;
    wire new_AGEMA_signal_34339 ;
    wire new_AGEMA_signal_34340 ;
    wire new_AGEMA_signal_34341 ;
    wire new_AGEMA_signal_34342 ;
    wire new_AGEMA_signal_34343 ;
    wire new_AGEMA_signal_34344 ;
    wire new_AGEMA_signal_34345 ;
    wire new_AGEMA_signal_34346 ;
    wire new_AGEMA_signal_34347 ;
    wire new_AGEMA_signal_34348 ;
    wire new_AGEMA_signal_34349 ;
    wire new_AGEMA_signal_34350 ;
    wire new_AGEMA_signal_34351 ;
    wire new_AGEMA_signal_34352 ;
    wire new_AGEMA_signal_34353 ;
    wire new_AGEMA_signal_34354 ;
    wire new_AGEMA_signal_34355 ;
    wire new_AGEMA_signal_34356 ;
    wire new_AGEMA_signal_34357 ;
    wire new_AGEMA_signal_34358 ;
    wire new_AGEMA_signal_34359 ;
    wire new_AGEMA_signal_34360 ;
    wire new_AGEMA_signal_34361 ;
    wire new_AGEMA_signal_34362 ;
    wire new_AGEMA_signal_34363 ;
    wire new_AGEMA_signal_34364 ;
    wire new_AGEMA_signal_34365 ;
    wire new_AGEMA_signal_34366 ;
    wire new_AGEMA_signal_34367 ;
    wire new_AGEMA_signal_34368 ;
    wire new_AGEMA_signal_34369 ;
    wire new_AGEMA_signal_34370 ;
    wire new_AGEMA_signal_34371 ;
    wire new_AGEMA_signal_34372 ;
    wire new_AGEMA_signal_34373 ;
    wire new_AGEMA_signal_34374 ;
    wire new_AGEMA_signal_34375 ;
    wire new_AGEMA_signal_34376 ;
    wire new_AGEMA_signal_34377 ;
    wire new_AGEMA_signal_34378 ;
    wire new_AGEMA_signal_34379 ;
    wire new_AGEMA_signal_34380 ;
    wire new_AGEMA_signal_34381 ;
    wire new_AGEMA_signal_34382 ;
    wire new_AGEMA_signal_34383 ;
    wire new_AGEMA_signal_34384 ;
    wire new_AGEMA_signal_34385 ;
    wire new_AGEMA_signal_34386 ;
    wire new_AGEMA_signal_34387 ;
    wire new_AGEMA_signal_34388 ;
    wire new_AGEMA_signal_34389 ;
    wire new_AGEMA_signal_34390 ;
    wire new_AGEMA_signal_34391 ;
    wire new_AGEMA_signal_34392 ;
    wire new_AGEMA_signal_34393 ;
    wire new_AGEMA_signal_34394 ;
    wire new_AGEMA_signal_34395 ;
    wire new_AGEMA_signal_34396 ;
    wire new_AGEMA_signal_34397 ;
    wire new_AGEMA_signal_34398 ;
    wire new_AGEMA_signal_34399 ;
    wire new_AGEMA_signal_34400 ;
    wire new_AGEMA_signal_34401 ;
    wire new_AGEMA_signal_34402 ;
    wire new_AGEMA_signal_34403 ;
    wire new_AGEMA_signal_34404 ;
    wire new_AGEMA_signal_34405 ;
    wire new_AGEMA_signal_34406 ;
    wire new_AGEMA_signal_34407 ;
    wire new_AGEMA_signal_34408 ;
    wire new_AGEMA_signal_34409 ;
    wire new_AGEMA_signal_34410 ;
    wire new_AGEMA_signal_34411 ;
    wire new_AGEMA_signal_34412 ;
    wire new_AGEMA_signal_34413 ;
    wire new_AGEMA_signal_34414 ;
    wire new_AGEMA_signal_34415 ;
    wire new_AGEMA_signal_34416 ;
    wire new_AGEMA_signal_34417 ;
    wire new_AGEMA_signal_34418 ;
    wire new_AGEMA_signal_34419 ;
    wire new_AGEMA_signal_34420 ;
    wire new_AGEMA_signal_34421 ;
    wire new_AGEMA_signal_34422 ;
    wire new_AGEMA_signal_34423 ;
    wire new_AGEMA_signal_34424 ;
    wire new_AGEMA_signal_34425 ;
    wire new_AGEMA_signal_34426 ;
    wire new_AGEMA_signal_34427 ;
    wire new_AGEMA_signal_34428 ;
    wire new_AGEMA_signal_34429 ;
    wire new_AGEMA_signal_34430 ;
    wire new_AGEMA_signal_34431 ;
    wire new_AGEMA_signal_34432 ;
    wire new_AGEMA_signal_34433 ;
    wire new_AGEMA_signal_34434 ;
    wire new_AGEMA_signal_34435 ;
    wire new_AGEMA_signal_34436 ;
    wire new_AGEMA_signal_34437 ;
    wire new_AGEMA_signal_34438 ;
    wire new_AGEMA_signal_34439 ;
    wire new_AGEMA_signal_34440 ;
    wire new_AGEMA_signal_34441 ;
    wire new_AGEMA_signal_34442 ;
    wire new_AGEMA_signal_34443 ;
    wire new_AGEMA_signal_34444 ;
    wire new_AGEMA_signal_34445 ;
    wire new_AGEMA_signal_34446 ;
    wire new_AGEMA_signal_34447 ;
    wire new_AGEMA_signal_34448 ;
    wire new_AGEMA_signal_34449 ;
    wire new_AGEMA_signal_34450 ;
    wire new_AGEMA_signal_34451 ;
    wire new_AGEMA_signal_34452 ;
    wire new_AGEMA_signal_34453 ;
    wire new_AGEMA_signal_34454 ;
    wire new_AGEMA_signal_34455 ;
    wire new_AGEMA_signal_34456 ;
    wire new_AGEMA_signal_34457 ;
    wire new_AGEMA_signal_34458 ;
    wire new_AGEMA_signal_34459 ;
    wire new_AGEMA_signal_34460 ;
    wire new_AGEMA_signal_34461 ;
    wire new_AGEMA_signal_34462 ;
    wire new_AGEMA_signal_34463 ;
    wire new_AGEMA_signal_34464 ;
    wire new_AGEMA_signal_34465 ;
    wire new_AGEMA_signal_34466 ;
    wire new_AGEMA_signal_34467 ;
    wire new_AGEMA_signal_34468 ;
    wire new_AGEMA_signal_34469 ;
    wire new_AGEMA_signal_34470 ;
    wire new_AGEMA_signal_34471 ;
    wire new_AGEMA_signal_34472 ;
    wire new_AGEMA_signal_34473 ;
    wire new_AGEMA_signal_34474 ;
    wire new_AGEMA_signal_34475 ;
    wire new_AGEMA_signal_34476 ;
    wire new_AGEMA_signal_34477 ;
    wire new_AGEMA_signal_34478 ;
    wire new_AGEMA_signal_34479 ;
    wire new_AGEMA_signal_34480 ;
    wire new_AGEMA_signal_34481 ;
    wire new_AGEMA_signal_34482 ;
    wire new_AGEMA_signal_34483 ;
    wire new_AGEMA_signal_34484 ;
    wire new_AGEMA_signal_34485 ;
    wire new_AGEMA_signal_34486 ;
    wire new_AGEMA_signal_34487 ;
    wire new_AGEMA_signal_34488 ;
    wire new_AGEMA_signal_34489 ;
    wire new_AGEMA_signal_34490 ;
    wire new_AGEMA_signal_34491 ;
    wire new_AGEMA_signal_34492 ;
    wire new_AGEMA_signal_34493 ;
    wire new_AGEMA_signal_34494 ;
    wire new_AGEMA_signal_34495 ;
    wire new_AGEMA_signal_34496 ;
    wire new_AGEMA_signal_34497 ;
    wire new_AGEMA_signal_34498 ;
    wire new_AGEMA_signal_34499 ;
    wire new_AGEMA_signal_34500 ;
    wire new_AGEMA_signal_34501 ;
    wire new_AGEMA_signal_34502 ;
    wire new_AGEMA_signal_34503 ;
    wire new_AGEMA_signal_34504 ;
    wire new_AGEMA_signal_34505 ;
    wire new_AGEMA_signal_34506 ;
    wire new_AGEMA_signal_34507 ;
    wire new_AGEMA_signal_34508 ;
    wire new_AGEMA_signal_34509 ;
    wire new_AGEMA_signal_34510 ;
    wire new_AGEMA_signal_34511 ;
    wire new_AGEMA_signal_34512 ;
    wire new_AGEMA_signal_34513 ;
    wire new_AGEMA_signal_34514 ;
    wire new_AGEMA_signal_34515 ;
    wire new_AGEMA_signal_34516 ;
    wire new_AGEMA_signal_34517 ;
    wire new_AGEMA_signal_34518 ;
    wire new_AGEMA_signal_34519 ;
    wire new_AGEMA_signal_34520 ;
    wire new_AGEMA_signal_34521 ;
    wire new_AGEMA_signal_34522 ;
    wire new_AGEMA_signal_34523 ;
    wire new_AGEMA_signal_34524 ;
    wire new_AGEMA_signal_34525 ;
    wire new_AGEMA_signal_34526 ;
    wire new_AGEMA_signal_34527 ;
    wire new_AGEMA_signal_34528 ;
    wire new_AGEMA_signal_34529 ;
    wire new_AGEMA_signal_34530 ;
    wire new_AGEMA_signal_34531 ;
    wire new_AGEMA_signal_34532 ;
    wire new_AGEMA_signal_34533 ;
    wire new_AGEMA_signal_34534 ;
    wire new_AGEMA_signal_34535 ;
    wire new_AGEMA_signal_34536 ;
    wire new_AGEMA_signal_34537 ;
    wire new_AGEMA_signal_34538 ;
    wire new_AGEMA_signal_34539 ;
    wire new_AGEMA_signal_34540 ;
    wire new_AGEMA_signal_34541 ;
    wire new_AGEMA_signal_34542 ;
    wire new_AGEMA_signal_34543 ;
    wire new_AGEMA_signal_34544 ;
    wire new_AGEMA_signal_34545 ;
    wire new_AGEMA_signal_34546 ;
    wire new_AGEMA_signal_34547 ;
    wire new_AGEMA_signal_34548 ;
    wire new_AGEMA_signal_34549 ;
    wire new_AGEMA_signal_34550 ;
    wire new_AGEMA_signal_34551 ;
    wire new_AGEMA_signal_34552 ;
    wire new_AGEMA_signal_34553 ;
    wire new_AGEMA_signal_34554 ;
    wire new_AGEMA_signal_34555 ;
    wire new_AGEMA_signal_34556 ;
    wire new_AGEMA_signal_34557 ;
    wire new_AGEMA_signal_34558 ;
    wire new_AGEMA_signal_34559 ;
    wire new_AGEMA_signal_34560 ;
    wire new_AGEMA_signal_34561 ;
    wire new_AGEMA_signal_34562 ;
    wire new_AGEMA_signal_34563 ;
    wire new_AGEMA_signal_34564 ;
    wire new_AGEMA_signal_34565 ;
    wire new_AGEMA_signal_34566 ;
    wire new_AGEMA_signal_34567 ;
    wire new_AGEMA_signal_34568 ;
    wire new_AGEMA_signal_34569 ;
    wire new_AGEMA_signal_34570 ;
    wire new_AGEMA_signal_34571 ;
    wire new_AGEMA_signal_34572 ;
    wire new_AGEMA_signal_34573 ;
    wire new_AGEMA_signal_34574 ;
    wire new_AGEMA_signal_34575 ;
    wire new_AGEMA_signal_34576 ;
    wire new_AGEMA_signal_34577 ;
    wire new_AGEMA_signal_34578 ;
    wire new_AGEMA_signal_34579 ;
    wire new_AGEMA_signal_34580 ;
    wire new_AGEMA_signal_34581 ;
    wire new_AGEMA_signal_34582 ;
    wire new_AGEMA_signal_34583 ;
    wire new_AGEMA_signal_34584 ;
    wire new_AGEMA_signal_34585 ;
    wire new_AGEMA_signal_34586 ;
    wire new_AGEMA_signal_34587 ;
    wire new_AGEMA_signal_34588 ;
    wire new_AGEMA_signal_34589 ;
    wire new_AGEMA_signal_34590 ;
    wire new_AGEMA_signal_34591 ;
    wire new_AGEMA_signal_34592 ;
    wire new_AGEMA_signal_34593 ;
    wire new_AGEMA_signal_34594 ;
    wire new_AGEMA_signal_34595 ;
    wire new_AGEMA_signal_34596 ;
    wire new_AGEMA_signal_34597 ;
    wire new_AGEMA_signal_34598 ;
    wire new_AGEMA_signal_34599 ;
    wire new_AGEMA_signal_34600 ;
    wire new_AGEMA_signal_34601 ;
    wire new_AGEMA_signal_34602 ;
    wire new_AGEMA_signal_34603 ;
    wire new_AGEMA_signal_34604 ;
    wire new_AGEMA_signal_34605 ;
    wire new_AGEMA_signal_34606 ;
    wire new_AGEMA_signal_34607 ;
    wire new_AGEMA_signal_34608 ;
    wire new_AGEMA_signal_34609 ;
    wire new_AGEMA_signal_34610 ;
    wire new_AGEMA_signal_34611 ;
    wire new_AGEMA_signal_34612 ;
    wire new_AGEMA_signal_34613 ;
    wire new_AGEMA_signal_34614 ;
    wire new_AGEMA_signal_34615 ;
    wire new_AGEMA_signal_34616 ;
    wire new_AGEMA_signal_34617 ;
    wire new_AGEMA_signal_34618 ;
    wire new_AGEMA_signal_34619 ;
    wire new_AGEMA_signal_34620 ;
    wire new_AGEMA_signal_34621 ;
    wire new_AGEMA_signal_34622 ;
    wire new_AGEMA_signal_34623 ;
    wire new_AGEMA_signal_34624 ;
    wire new_AGEMA_signal_34625 ;
    wire new_AGEMA_signal_34626 ;
    wire new_AGEMA_signal_34627 ;
    wire new_AGEMA_signal_34628 ;
    wire new_AGEMA_signal_34629 ;
    wire new_AGEMA_signal_34630 ;
    wire new_AGEMA_signal_34631 ;
    wire new_AGEMA_signal_34632 ;
    wire new_AGEMA_signal_34633 ;
    wire new_AGEMA_signal_34634 ;
    wire new_AGEMA_signal_34635 ;
    wire new_AGEMA_signal_34636 ;
    wire new_AGEMA_signal_34637 ;
    wire new_AGEMA_signal_34638 ;
    wire new_AGEMA_signal_34639 ;
    wire new_AGEMA_signal_34640 ;
    wire new_AGEMA_signal_34641 ;
    wire new_AGEMA_signal_34642 ;
    wire new_AGEMA_signal_34643 ;
    wire new_AGEMA_signal_34644 ;
    wire new_AGEMA_signal_34645 ;
    wire new_AGEMA_signal_34646 ;
    wire new_AGEMA_signal_34647 ;
    wire new_AGEMA_signal_34648 ;
    wire new_AGEMA_signal_34649 ;
    wire new_AGEMA_signal_34650 ;
    wire new_AGEMA_signal_34651 ;
    wire new_AGEMA_signal_34652 ;
    wire new_AGEMA_signal_34653 ;
    wire new_AGEMA_signal_34654 ;
    wire new_AGEMA_signal_34655 ;
    wire new_AGEMA_signal_34656 ;
    wire new_AGEMA_signal_34657 ;
    wire new_AGEMA_signal_34658 ;
    wire new_AGEMA_signal_34659 ;
    wire new_AGEMA_signal_34660 ;
    wire new_AGEMA_signal_34661 ;
    wire new_AGEMA_signal_34662 ;
    wire new_AGEMA_signal_34663 ;
    wire new_AGEMA_signal_34664 ;
    wire new_AGEMA_signal_34665 ;
    wire new_AGEMA_signal_34666 ;
    wire new_AGEMA_signal_34667 ;
    wire new_AGEMA_signal_34668 ;
    wire new_AGEMA_signal_34669 ;
    wire new_AGEMA_signal_34670 ;
    wire new_AGEMA_signal_34671 ;
    wire new_AGEMA_signal_34672 ;
    wire new_AGEMA_signal_34673 ;
    wire new_AGEMA_signal_34674 ;
    wire new_AGEMA_signal_34675 ;
    wire new_AGEMA_signal_34676 ;
    wire new_AGEMA_signal_34677 ;
    wire new_AGEMA_signal_34678 ;
    wire new_AGEMA_signal_34679 ;
    wire new_AGEMA_signal_34680 ;
    wire new_AGEMA_signal_34681 ;
    wire new_AGEMA_signal_34682 ;
    wire new_AGEMA_signal_34683 ;
    wire new_AGEMA_signal_34684 ;
    wire new_AGEMA_signal_34685 ;
    wire new_AGEMA_signal_34686 ;
    wire new_AGEMA_signal_34687 ;
    wire new_AGEMA_signal_34688 ;
    wire new_AGEMA_signal_34689 ;
    wire new_AGEMA_signal_34690 ;
    wire new_AGEMA_signal_34691 ;
    wire new_AGEMA_signal_34692 ;
    wire new_AGEMA_signal_34693 ;
    wire new_AGEMA_signal_34694 ;
    wire new_AGEMA_signal_34695 ;
    wire new_AGEMA_signal_34696 ;
    wire new_AGEMA_signal_34697 ;
    wire new_AGEMA_signal_34698 ;
    wire new_AGEMA_signal_34699 ;
    wire new_AGEMA_signal_34700 ;
    wire new_AGEMA_signal_34701 ;
    wire new_AGEMA_signal_34702 ;
    wire new_AGEMA_signal_34703 ;
    wire new_AGEMA_signal_34704 ;
    wire new_AGEMA_signal_34705 ;
    wire new_AGEMA_signal_34706 ;
    wire new_AGEMA_signal_34707 ;
    wire new_AGEMA_signal_34708 ;
    wire new_AGEMA_signal_34709 ;
    wire new_AGEMA_signal_34710 ;
    wire new_AGEMA_signal_34711 ;
    wire new_AGEMA_signal_34712 ;
    wire new_AGEMA_signal_34713 ;
    wire new_AGEMA_signal_34714 ;
    wire new_AGEMA_signal_34715 ;
    wire new_AGEMA_signal_34716 ;
    wire new_AGEMA_signal_34717 ;
    wire new_AGEMA_signal_34718 ;
    wire new_AGEMA_signal_34719 ;
    wire new_AGEMA_signal_34720 ;
    wire new_AGEMA_signal_34721 ;
    wire new_AGEMA_signal_34722 ;
    wire new_AGEMA_signal_34723 ;
    wire new_AGEMA_signal_34724 ;
    wire new_AGEMA_signal_34725 ;
    wire new_AGEMA_signal_34726 ;
    wire new_AGEMA_signal_34727 ;
    wire new_AGEMA_signal_34728 ;
    wire new_AGEMA_signal_34729 ;
    wire new_AGEMA_signal_34730 ;
    wire new_AGEMA_signal_34731 ;
    wire new_AGEMA_signal_34732 ;
    wire new_AGEMA_signal_34733 ;
    wire new_AGEMA_signal_34734 ;
    wire new_AGEMA_signal_34735 ;
    wire new_AGEMA_signal_34736 ;
    wire new_AGEMA_signal_34737 ;
    wire new_AGEMA_signal_34738 ;
    wire new_AGEMA_signal_34739 ;
    wire new_AGEMA_signal_34740 ;
    wire new_AGEMA_signal_34741 ;
    wire new_AGEMA_signal_34742 ;
    wire new_AGEMA_signal_34743 ;
    wire new_AGEMA_signal_34744 ;
    wire new_AGEMA_signal_34745 ;
    wire new_AGEMA_signal_34746 ;
    wire new_AGEMA_signal_34747 ;
    wire new_AGEMA_signal_34748 ;
    wire new_AGEMA_signal_34749 ;
    wire new_AGEMA_signal_34750 ;
    wire new_AGEMA_signal_34751 ;
    wire new_AGEMA_signal_34752 ;
    wire new_AGEMA_signal_34753 ;
    wire new_AGEMA_signal_34754 ;
    wire new_AGEMA_signal_34755 ;
    wire new_AGEMA_signal_34756 ;
    wire new_AGEMA_signal_34757 ;
    wire new_AGEMA_signal_34758 ;
    wire new_AGEMA_signal_34759 ;
    wire new_AGEMA_signal_34760 ;
    wire new_AGEMA_signal_34761 ;
    wire new_AGEMA_signal_34762 ;
    wire new_AGEMA_signal_34763 ;
    wire new_AGEMA_signal_34764 ;
    wire new_AGEMA_signal_34765 ;
    wire new_AGEMA_signal_34766 ;
    wire new_AGEMA_signal_34767 ;
    wire new_AGEMA_signal_34768 ;
    wire new_AGEMA_signal_34769 ;
    wire new_AGEMA_signal_34770 ;
    wire new_AGEMA_signal_34771 ;
    wire new_AGEMA_signal_34772 ;
    wire new_AGEMA_signal_34773 ;
    wire new_AGEMA_signal_34774 ;
    wire new_AGEMA_signal_34775 ;
    wire new_AGEMA_signal_34776 ;
    wire new_AGEMA_signal_34777 ;
    wire new_AGEMA_signal_34778 ;
    wire new_AGEMA_signal_34779 ;
    wire new_AGEMA_signal_34780 ;
    wire new_AGEMA_signal_34781 ;
    wire new_AGEMA_signal_34782 ;
    wire new_AGEMA_signal_34783 ;
    wire new_AGEMA_signal_34784 ;
    wire new_AGEMA_signal_34785 ;
    wire new_AGEMA_signal_34786 ;
    wire new_AGEMA_signal_34787 ;
    wire new_AGEMA_signal_34788 ;
    wire new_AGEMA_signal_34789 ;
    wire new_AGEMA_signal_34790 ;
    wire new_AGEMA_signal_34791 ;
    wire new_AGEMA_signal_34792 ;
    wire new_AGEMA_signal_34793 ;
    wire new_AGEMA_signal_34794 ;
    wire new_AGEMA_signal_34795 ;
    wire new_AGEMA_signal_34796 ;
    wire new_AGEMA_signal_34797 ;
    wire new_AGEMA_signal_34798 ;
    wire new_AGEMA_signal_34799 ;
    wire new_AGEMA_signal_34800 ;
    wire new_AGEMA_signal_34801 ;
    wire new_AGEMA_signal_34802 ;
    wire new_AGEMA_signal_34803 ;
    wire new_AGEMA_signal_34804 ;
    wire new_AGEMA_signal_34805 ;
    wire new_AGEMA_signal_34806 ;
    wire new_AGEMA_signal_34807 ;
    wire new_AGEMA_signal_34808 ;
    wire new_AGEMA_signal_34809 ;
    wire new_AGEMA_signal_34810 ;
    wire new_AGEMA_signal_34811 ;
    wire new_AGEMA_signal_34812 ;
    wire new_AGEMA_signal_34813 ;
    wire new_AGEMA_signal_34814 ;
    wire new_AGEMA_signal_34815 ;
    wire new_AGEMA_signal_34816 ;
    wire new_AGEMA_signal_34817 ;
    wire new_AGEMA_signal_34818 ;
    wire new_AGEMA_signal_34819 ;
    wire new_AGEMA_signal_34820 ;
    wire new_AGEMA_signal_34821 ;
    wire new_AGEMA_signal_34822 ;
    wire new_AGEMA_signal_34823 ;
    wire new_AGEMA_signal_34824 ;
    wire new_AGEMA_signal_34825 ;
    wire new_AGEMA_signal_34826 ;
    wire new_AGEMA_signal_34827 ;
    wire new_AGEMA_signal_34828 ;
    wire new_AGEMA_signal_34829 ;
    wire new_AGEMA_signal_34830 ;
    wire new_AGEMA_signal_34831 ;
    wire new_AGEMA_signal_34832 ;
    wire new_AGEMA_signal_34833 ;
    wire new_AGEMA_signal_34834 ;
    wire new_AGEMA_signal_34835 ;
    wire new_AGEMA_signal_34836 ;
    wire new_AGEMA_signal_34837 ;
    wire new_AGEMA_signal_34838 ;
    wire new_AGEMA_signal_34839 ;
    wire new_AGEMA_signal_34840 ;
    wire new_AGEMA_signal_34841 ;
    wire new_AGEMA_signal_34842 ;
    wire new_AGEMA_signal_34843 ;
    wire new_AGEMA_signal_34844 ;
    wire new_AGEMA_signal_34845 ;
    wire new_AGEMA_signal_34846 ;
    wire new_AGEMA_signal_34847 ;
    wire new_AGEMA_signal_34848 ;
    wire new_AGEMA_signal_34849 ;
    wire new_AGEMA_signal_34850 ;
    wire new_AGEMA_signal_34851 ;
    wire new_AGEMA_signal_34852 ;
    wire new_AGEMA_signal_34853 ;
    wire new_AGEMA_signal_34854 ;
    wire new_AGEMA_signal_34855 ;
    wire new_AGEMA_signal_34856 ;
    wire new_AGEMA_signal_34857 ;
    wire new_AGEMA_signal_34858 ;
    wire new_AGEMA_signal_34859 ;
    wire new_AGEMA_signal_34860 ;
    wire new_AGEMA_signal_34861 ;
    wire new_AGEMA_signal_34862 ;
    wire new_AGEMA_signal_34863 ;
    wire new_AGEMA_signal_34864 ;
    wire new_AGEMA_signal_34865 ;
    wire new_AGEMA_signal_34866 ;
    wire new_AGEMA_signal_34867 ;
    wire new_AGEMA_signal_34868 ;
    wire new_AGEMA_signal_34869 ;
    wire new_AGEMA_signal_34870 ;
    wire new_AGEMA_signal_34871 ;
    wire new_AGEMA_signal_34872 ;
    wire new_AGEMA_signal_34873 ;
    wire new_AGEMA_signal_34874 ;
    wire new_AGEMA_signal_34875 ;
    wire new_AGEMA_signal_34876 ;
    wire new_AGEMA_signal_34877 ;
    wire new_AGEMA_signal_34878 ;
    wire new_AGEMA_signal_34879 ;
    wire new_AGEMA_signal_34880 ;
    wire new_AGEMA_signal_34881 ;
    wire new_AGEMA_signal_34882 ;
    wire new_AGEMA_signal_34883 ;
    wire new_AGEMA_signal_34884 ;
    wire new_AGEMA_signal_34885 ;
    wire new_AGEMA_signal_34886 ;
    wire new_AGEMA_signal_34887 ;
    wire new_AGEMA_signal_34888 ;
    wire new_AGEMA_signal_34889 ;
    wire new_AGEMA_signal_34890 ;
    wire new_AGEMA_signal_34891 ;
    wire new_AGEMA_signal_34892 ;
    wire new_AGEMA_signal_34893 ;
    wire new_AGEMA_signal_34894 ;
    wire new_AGEMA_signal_34895 ;
    wire new_AGEMA_signal_34896 ;
    wire new_AGEMA_signal_34897 ;
    wire new_AGEMA_signal_34898 ;
    wire new_AGEMA_signal_34899 ;
    wire new_AGEMA_signal_34900 ;
    wire new_AGEMA_signal_34901 ;
    wire new_AGEMA_signal_34902 ;
    wire new_AGEMA_signal_34903 ;
    wire new_AGEMA_signal_34904 ;
    wire new_AGEMA_signal_34905 ;
    wire new_AGEMA_signal_34906 ;
    wire new_AGEMA_signal_34907 ;
    wire new_AGEMA_signal_34908 ;
    wire new_AGEMA_signal_34909 ;
    wire new_AGEMA_signal_34910 ;
    wire new_AGEMA_signal_34911 ;
    wire new_AGEMA_signal_34912 ;
    wire new_AGEMA_signal_34913 ;
    wire new_AGEMA_signal_34914 ;
    wire new_AGEMA_signal_34915 ;
    wire new_AGEMA_signal_34916 ;
    wire new_AGEMA_signal_34917 ;
    wire new_AGEMA_signal_34918 ;
    wire new_AGEMA_signal_34919 ;
    wire new_AGEMA_signal_34920 ;
    wire new_AGEMA_signal_34921 ;
    wire new_AGEMA_signal_34922 ;
    wire new_AGEMA_signal_34923 ;
    wire new_AGEMA_signal_34924 ;
    wire new_AGEMA_signal_34925 ;
    wire new_AGEMA_signal_34926 ;
    wire new_AGEMA_signal_34927 ;
    wire new_AGEMA_signal_34928 ;
    wire new_AGEMA_signal_34929 ;
    wire new_AGEMA_signal_34930 ;
    wire new_AGEMA_signal_34931 ;
    wire new_AGEMA_signal_34932 ;
    wire new_AGEMA_signal_34933 ;
    wire new_AGEMA_signal_34934 ;
    wire new_AGEMA_signal_34935 ;
    wire new_AGEMA_signal_34936 ;
    wire new_AGEMA_signal_34937 ;
    wire new_AGEMA_signal_34938 ;
    wire new_AGEMA_signal_34939 ;
    wire new_AGEMA_signal_34940 ;
    wire new_AGEMA_signal_34941 ;
    wire new_AGEMA_signal_34942 ;
    wire new_AGEMA_signal_34943 ;
    wire new_AGEMA_signal_34944 ;
    wire new_AGEMA_signal_34945 ;
    wire new_AGEMA_signal_34946 ;
    wire new_AGEMA_signal_34947 ;
    wire new_AGEMA_signal_34948 ;
    wire new_AGEMA_signal_34949 ;
    wire new_AGEMA_signal_34950 ;
    wire new_AGEMA_signal_34951 ;
    wire new_AGEMA_signal_34952 ;
    wire new_AGEMA_signal_34953 ;
    wire new_AGEMA_signal_34954 ;
    wire new_AGEMA_signal_34955 ;
    wire new_AGEMA_signal_34956 ;
    wire new_AGEMA_signal_34957 ;
    wire new_AGEMA_signal_34958 ;
    wire new_AGEMA_signal_34959 ;
    wire new_AGEMA_signal_34960 ;
    wire new_AGEMA_signal_34961 ;
    wire new_AGEMA_signal_34962 ;
    wire new_AGEMA_signal_34963 ;
    wire new_AGEMA_signal_34964 ;
    wire new_AGEMA_signal_34965 ;
    wire new_AGEMA_signal_34966 ;
    wire new_AGEMA_signal_34967 ;
    wire new_AGEMA_signal_34968 ;
    wire new_AGEMA_signal_34969 ;
    wire new_AGEMA_signal_34970 ;
    wire new_AGEMA_signal_34971 ;
    wire new_AGEMA_signal_34972 ;
    wire new_AGEMA_signal_34973 ;
    wire new_AGEMA_signal_34974 ;
    wire new_AGEMA_signal_34975 ;
    wire new_AGEMA_signal_34976 ;
    wire new_AGEMA_signal_34977 ;
    wire new_AGEMA_signal_34978 ;
    wire new_AGEMA_signal_34979 ;
    wire new_AGEMA_signal_34980 ;
    wire new_AGEMA_signal_34981 ;
    wire new_AGEMA_signal_34982 ;
    wire new_AGEMA_signal_34983 ;
    wire new_AGEMA_signal_34984 ;
    wire new_AGEMA_signal_34985 ;
    wire new_AGEMA_signal_34986 ;
    wire new_AGEMA_signal_34987 ;
    wire new_AGEMA_signal_34988 ;
    wire new_AGEMA_signal_34989 ;
    wire new_AGEMA_signal_34990 ;
    wire new_AGEMA_signal_34991 ;
    wire new_AGEMA_signal_34992 ;
    wire new_AGEMA_signal_34993 ;
    wire new_AGEMA_signal_34994 ;
    wire new_AGEMA_signal_34995 ;
    wire new_AGEMA_signal_34996 ;
    wire new_AGEMA_signal_34997 ;
    wire new_AGEMA_signal_34998 ;
    wire new_AGEMA_signal_34999 ;
    wire new_AGEMA_signal_35000 ;
    wire new_AGEMA_signal_35001 ;
    wire new_AGEMA_signal_35002 ;
    wire new_AGEMA_signal_35003 ;
    wire new_AGEMA_signal_35004 ;
    wire new_AGEMA_signal_35005 ;
    wire new_AGEMA_signal_35006 ;
    wire new_AGEMA_signal_35007 ;
    wire new_AGEMA_signal_35008 ;
    wire new_AGEMA_signal_35009 ;
    wire new_AGEMA_signal_35010 ;
    wire new_AGEMA_signal_35011 ;
    wire new_AGEMA_signal_35012 ;
    wire new_AGEMA_signal_35013 ;
    wire new_AGEMA_signal_35014 ;
    wire new_AGEMA_signal_35015 ;
    wire new_AGEMA_signal_35016 ;
    wire new_AGEMA_signal_35017 ;
    wire new_AGEMA_signal_35018 ;
    wire new_AGEMA_signal_35019 ;
    wire new_AGEMA_signal_35020 ;
    wire new_AGEMA_signal_35021 ;
    wire new_AGEMA_signal_35022 ;
    wire new_AGEMA_signal_35023 ;
    wire new_AGEMA_signal_35024 ;
    wire new_AGEMA_signal_35025 ;
    wire new_AGEMA_signal_35026 ;
    wire new_AGEMA_signal_35027 ;
    wire new_AGEMA_signal_35028 ;
    wire new_AGEMA_signal_35029 ;
    wire new_AGEMA_signal_35030 ;
    wire new_AGEMA_signal_35031 ;
    wire new_AGEMA_signal_35032 ;
    wire new_AGEMA_signal_35033 ;
    wire new_AGEMA_signal_35034 ;
    wire new_AGEMA_signal_35035 ;
    wire new_AGEMA_signal_35036 ;
    wire new_AGEMA_signal_35037 ;
    wire new_AGEMA_signal_35038 ;
    wire new_AGEMA_signal_35039 ;
    wire new_AGEMA_signal_35040 ;
    wire new_AGEMA_signal_35041 ;
    wire new_AGEMA_signal_35042 ;
    wire new_AGEMA_signal_35043 ;
    wire new_AGEMA_signal_35044 ;
    wire new_AGEMA_signal_35045 ;
    wire new_AGEMA_signal_35046 ;
    wire new_AGEMA_signal_35047 ;
    wire new_AGEMA_signal_35048 ;
    wire new_AGEMA_signal_35049 ;
    wire new_AGEMA_signal_35050 ;
    wire new_AGEMA_signal_35051 ;
    wire new_AGEMA_signal_35052 ;
    wire new_AGEMA_signal_35053 ;
    wire new_AGEMA_signal_35054 ;
    wire new_AGEMA_signal_35055 ;
    wire new_AGEMA_signal_35056 ;
    wire new_AGEMA_signal_35057 ;
    wire new_AGEMA_signal_35058 ;
    wire new_AGEMA_signal_35059 ;
    wire new_AGEMA_signal_35060 ;
    wire new_AGEMA_signal_35061 ;
    wire new_AGEMA_signal_35062 ;
    wire new_AGEMA_signal_35063 ;
    wire new_AGEMA_signal_35064 ;
    wire new_AGEMA_signal_35065 ;
    wire new_AGEMA_signal_35066 ;
    wire new_AGEMA_signal_35067 ;
    wire new_AGEMA_signal_35068 ;
    wire new_AGEMA_signal_35069 ;
    wire new_AGEMA_signal_35070 ;
    wire new_AGEMA_signal_35071 ;
    wire new_AGEMA_signal_35072 ;
    wire new_AGEMA_signal_35073 ;
    wire new_AGEMA_signal_35074 ;
    wire new_AGEMA_signal_35075 ;
    wire new_AGEMA_signal_35076 ;
    wire new_AGEMA_signal_35077 ;
    wire new_AGEMA_signal_35078 ;
    wire new_AGEMA_signal_35079 ;
    wire new_AGEMA_signal_35080 ;
    wire new_AGEMA_signal_35081 ;
    wire new_AGEMA_signal_35082 ;
    wire new_AGEMA_signal_35083 ;
    wire new_AGEMA_signal_35084 ;
    wire new_AGEMA_signal_35085 ;
    wire new_AGEMA_signal_35086 ;
    wire new_AGEMA_signal_35087 ;
    wire new_AGEMA_signal_35088 ;
    wire new_AGEMA_signal_35089 ;
    wire new_AGEMA_signal_35090 ;
    wire new_AGEMA_signal_35091 ;
    wire new_AGEMA_signal_35092 ;
    wire new_AGEMA_signal_35093 ;
    wire new_AGEMA_signal_35094 ;
    wire new_AGEMA_signal_35095 ;
    wire new_AGEMA_signal_35096 ;
    wire new_AGEMA_signal_35097 ;
    wire new_AGEMA_signal_35098 ;
    wire new_AGEMA_signal_35099 ;
    wire new_AGEMA_signal_35100 ;
    wire new_AGEMA_signal_35101 ;
    wire new_AGEMA_signal_35102 ;
    wire new_AGEMA_signal_35103 ;
    wire new_AGEMA_signal_35104 ;
    wire new_AGEMA_signal_35105 ;
    wire new_AGEMA_signal_35106 ;
    wire new_AGEMA_signal_35107 ;
    wire new_AGEMA_signal_35108 ;
    wire new_AGEMA_signal_35109 ;
    wire new_AGEMA_signal_35110 ;
    wire new_AGEMA_signal_35111 ;
    wire new_AGEMA_signal_35112 ;
    wire new_AGEMA_signal_35113 ;
    wire new_AGEMA_signal_35114 ;
    wire new_AGEMA_signal_35115 ;
    wire new_AGEMA_signal_35116 ;
    wire new_AGEMA_signal_35117 ;
    wire new_AGEMA_signal_35118 ;
    wire new_AGEMA_signal_35119 ;
    wire new_AGEMA_signal_35120 ;
    wire new_AGEMA_signal_35121 ;
    wire new_AGEMA_signal_35122 ;
    wire new_AGEMA_signal_35123 ;
    wire new_AGEMA_signal_35124 ;
    wire new_AGEMA_signal_35125 ;
    wire new_AGEMA_signal_35126 ;
    wire new_AGEMA_signal_35127 ;
    wire new_AGEMA_signal_35128 ;
    wire new_AGEMA_signal_35129 ;
    wire new_AGEMA_signal_35130 ;
    wire new_AGEMA_signal_35131 ;
    wire new_AGEMA_signal_35132 ;
    wire new_AGEMA_signal_35133 ;
    wire new_AGEMA_signal_35134 ;
    wire new_AGEMA_signal_35135 ;
    wire new_AGEMA_signal_35136 ;
    wire new_AGEMA_signal_35137 ;
    wire new_AGEMA_signal_35138 ;
    wire new_AGEMA_signal_35139 ;
    wire new_AGEMA_signal_35140 ;
    wire new_AGEMA_signal_35141 ;
    wire new_AGEMA_signal_35142 ;
    wire new_AGEMA_signal_35143 ;
    wire new_AGEMA_signal_35144 ;
    wire new_AGEMA_signal_35145 ;
    wire new_AGEMA_signal_35146 ;
    wire new_AGEMA_signal_35147 ;
    wire new_AGEMA_signal_35148 ;
    wire new_AGEMA_signal_35149 ;
    wire new_AGEMA_signal_35150 ;
    wire new_AGEMA_signal_35151 ;
    wire new_AGEMA_signal_35152 ;
    wire new_AGEMA_signal_35153 ;
    wire new_AGEMA_signal_35154 ;
    wire new_AGEMA_signal_35155 ;
    wire new_AGEMA_signal_35156 ;
    wire new_AGEMA_signal_35157 ;
    wire new_AGEMA_signal_35158 ;
    wire new_AGEMA_signal_35159 ;
    wire new_AGEMA_signal_35160 ;
    wire new_AGEMA_signal_35161 ;
    wire new_AGEMA_signal_35162 ;
    wire new_AGEMA_signal_35163 ;
    wire new_AGEMA_signal_35164 ;
    wire new_AGEMA_signal_35165 ;
    wire new_AGEMA_signal_35166 ;
    wire new_AGEMA_signal_35167 ;
    wire new_AGEMA_signal_35168 ;
    wire new_AGEMA_signal_35169 ;
    wire new_AGEMA_signal_35170 ;
    wire new_AGEMA_signal_35171 ;
    wire new_AGEMA_signal_35172 ;
    wire new_AGEMA_signal_35173 ;
    wire new_AGEMA_signal_35174 ;
    wire new_AGEMA_signal_35175 ;
    wire new_AGEMA_signal_35176 ;
    wire new_AGEMA_signal_35177 ;
    wire new_AGEMA_signal_35178 ;
    wire new_AGEMA_signal_35179 ;
    wire new_AGEMA_signal_35180 ;
    wire new_AGEMA_signal_35181 ;
    wire new_AGEMA_signal_35182 ;
    wire new_AGEMA_signal_35183 ;
    wire new_AGEMA_signal_35184 ;
    wire new_AGEMA_signal_35185 ;
    wire new_AGEMA_signal_35186 ;
    wire new_AGEMA_signal_35187 ;
    wire new_AGEMA_signal_35188 ;
    wire new_AGEMA_signal_35189 ;
    wire new_AGEMA_signal_35190 ;
    wire new_AGEMA_signal_35191 ;
    wire new_AGEMA_signal_35192 ;
    wire new_AGEMA_signal_35193 ;
    wire new_AGEMA_signal_35194 ;
    wire new_AGEMA_signal_35195 ;
    wire new_AGEMA_signal_35196 ;
    wire new_AGEMA_signal_35197 ;
    wire new_AGEMA_signal_35198 ;
    wire new_AGEMA_signal_35199 ;
    wire new_AGEMA_signal_35200 ;
    wire new_AGEMA_signal_35201 ;
    wire new_AGEMA_signal_35202 ;
    wire new_AGEMA_signal_35203 ;
    wire new_AGEMA_signal_35204 ;
    wire new_AGEMA_signal_35205 ;
    wire new_AGEMA_signal_35206 ;
    wire new_AGEMA_signal_35207 ;
    wire new_AGEMA_signal_35208 ;
    wire new_AGEMA_signal_35209 ;
    wire new_AGEMA_signal_35210 ;
    wire new_AGEMA_signal_35211 ;
    wire new_AGEMA_signal_35212 ;
    wire new_AGEMA_signal_35213 ;
    wire new_AGEMA_signal_35214 ;
    wire new_AGEMA_signal_35215 ;
    wire new_AGEMA_signal_35216 ;
    wire new_AGEMA_signal_35217 ;
    wire new_AGEMA_signal_35218 ;
    wire new_AGEMA_signal_35219 ;
    wire new_AGEMA_signal_35220 ;
    wire new_AGEMA_signal_35221 ;
    wire new_AGEMA_signal_35222 ;
    wire new_AGEMA_signal_35223 ;
    wire new_AGEMA_signal_35224 ;
    wire new_AGEMA_signal_35225 ;
    wire new_AGEMA_signal_35226 ;
    wire new_AGEMA_signal_35227 ;
    wire new_AGEMA_signal_35228 ;
    wire new_AGEMA_signal_35229 ;
    wire new_AGEMA_signal_35230 ;
    wire new_AGEMA_signal_35231 ;
    wire new_AGEMA_signal_35232 ;
    wire new_AGEMA_signal_35233 ;
    wire new_AGEMA_signal_35234 ;
    wire new_AGEMA_signal_35235 ;
    wire new_AGEMA_signal_35236 ;
    wire new_AGEMA_signal_35237 ;
    wire new_AGEMA_signal_35238 ;
    wire new_AGEMA_signal_35239 ;
    wire new_AGEMA_signal_35240 ;
    wire new_AGEMA_signal_35241 ;
    wire new_AGEMA_signal_35242 ;
    wire new_AGEMA_signal_35243 ;
    wire new_AGEMA_signal_35244 ;
    wire new_AGEMA_signal_35245 ;
    wire new_AGEMA_signal_35246 ;
    wire new_AGEMA_signal_35247 ;
    wire new_AGEMA_signal_35248 ;
    wire new_AGEMA_signal_35249 ;
    wire new_AGEMA_signal_35250 ;
    wire new_AGEMA_signal_35251 ;
    wire new_AGEMA_signal_35252 ;
    wire new_AGEMA_signal_35253 ;
    wire new_AGEMA_signal_35254 ;
    wire new_AGEMA_signal_35255 ;
    wire new_AGEMA_signal_35256 ;
    wire new_AGEMA_signal_35257 ;
    wire new_AGEMA_signal_35258 ;
    wire new_AGEMA_signal_35259 ;
    wire new_AGEMA_signal_35260 ;
    wire new_AGEMA_signal_35261 ;
    wire new_AGEMA_signal_35262 ;
    wire new_AGEMA_signal_35263 ;
    wire new_AGEMA_signal_35264 ;
    wire new_AGEMA_signal_35265 ;
    wire new_AGEMA_signal_35266 ;
    wire new_AGEMA_signal_35267 ;
    wire new_AGEMA_signal_35268 ;
    wire new_AGEMA_signal_35269 ;
    wire new_AGEMA_signal_35270 ;
    wire new_AGEMA_signal_35271 ;
    wire new_AGEMA_signal_35272 ;
    wire new_AGEMA_signal_35273 ;
    wire new_AGEMA_signal_35274 ;
    wire new_AGEMA_signal_35275 ;
    wire new_AGEMA_signal_35276 ;
    wire new_AGEMA_signal_35277 ;
    wire new_AGEMA_signal_35278 ;
    wire new_AGEMA_signal_35279 ;
    wire new_AGEMA_signal_35280 ;
    wire new_AGEMA_signal_35281 ;
    wire new_AGEMA_signal_35282 ;
    wire new_AGEMA_signal_35283 ;
    wire new_AGEMA_signal_35284 ;
    wire new_AGEMA_signal_35285 ;
    wire new_AGEMA_signal_35286 ;
    wire new_AGEMA_signal_35287 ;
    wire new_AGEMA_signal_35288 ;
    wire new_AGEMA_signal_35289 ;
    wire new_AGEMA_signal_35290 ;
    wire new_AGEMA_signal_35291 ;
    wire new_AGEMA_signal_35292 ;
    wire new_AGEMA_signal_35293 ;
    wire new_AGEMA_signal_35294 ;
    wire new_AGEMA_signal_35295 ;
    wire new_AGEMA_signal_35296 ;
    wire new_AGEMA_signal_35297 ;
    wire new_AGEMA_signal_35298 ;
    wire new_AGEMA_signal_35299 ;
    wire new_AGEMA_signal_35300 ;
    wire new_AGEMA_signal_35301 ;
    wire new_AGEMA_signal_35302 ;
    wire new_AGEMA_signal_35303 ;
    wire new_AGEMA_signal_35304 ;
    wire new_AGEMA_signal_35305 ;
    wire new_AGEMA_signal_35306 ;
    wire new_AGEMA_signal_35307 ;
    wire new_AGEMA_signal_35308 ;
    wire new_AGEMA_signal_35309 ;
    wire new_AGEMA_signal_35310 ;
    wire new_AGEMA_signal_35311 ;
    wire new_AGEMA_signal_35312 ;
    wire new_AGEMA_signal_35313 ;
    wire new_AGEMA_signal_35314 ;
    wire new_AGEMA_signal_35315 ;
    wire new_AGEMA_signal_35316 ;
    wire new_AGEMA_signal_35317 ;
    wire new_AGEMA_signal_35318 ;
    wire new_AGEMA_signal_35319 ;
    wire new_AGEMA_signal_35320 ;
    wire new_AGEMA_signal_35321 ;
    wire new_AGEMA_signal_35322 ;
    wire new_AGEMA_signal_35323 ;
    wire new_AGEMA_signal_35324 ;
    wire new_AGEMA_signal_35325 ;
    wire new_AGEMA_signal_35326 ;
    wire new_AGEMA_signal_35327 ;
    wire new_AGEMA_signal_35328 ;
    wire new_AGEMA_signal_35329 ;
    wire new_AGEMA_signal_35330 ;
    wire new_AGEMA_signal_35331 ;
    wire new_AGEMA_signal_35332 ;
    wire new_AGEMA_signal_35333 ;
    wire new_AGEMA_signal_35334 ;
    wire new_AGEMA_signal_35335 ;
    wire new_AGEMA_signal_35336 ;
    wire new_AGEMA_signal_35337 ;
    wire new_AGEMA_signal_35338 ;
    wire new_AGEMA_signal_35339 ;
    wire new_AGEMA_signal_35340 ;
    wire new_AGEMA_signal_35341 ;
    wire new_AGEMA_signal_35342 ;
    wire new_AGEMA_signal_35343 ;
    wire new_AGEMA_signal_35344 ;
    wire new_AGEMA_signal_35345 ;
    wire new_AGEMA_signal_35346 ;
    wire new_AGEMA_signal_35347 ;
    wire new_AGEMA_signal_35348 ;
    wire new_AGEMA_signal_35349 ;
    wire new_AGEMA_signal_35350 ;
    wire new_AGEMA_signal_35351 ;
    wire new_AGEMA_signal_35352 ;
    wire new_AGEMA_signal_35353 ;
    wire new_AGEMA_signal_35354 ;
    wire new_AGEMA_signal_35355 ;
    wire new_AGEMA_signal_35356 ;
    wire new_AGEMA_signal_35357 ;
    wire new_AGEMA_signal_35358 ;
    wire new_AGEMA_signal_35359 ;
    wire new_AGEMA_signal_35360 ;
    wire new_AGEMA_signal_35361 ;
    wire new_AGEMA_signal_35362 ;
    wire new_AGEMA_signal_35363 ;
    wire new_AGEMA_signal_35364 ;
    wire new_AGEMA_signal_35365 ;
    wire new_AGEMA_signal_35366 ;
    wire new_AGEMA_signal_35367 ;
    wire new_AGEMA_signal_35368 ;
    wire new_AGEMA_signal_35369 ;
    wire new_AGEMA_signal_35370 ;
    wire new_AGEMA_signal_35371 ;
    wire new_AGEMA_signal_35372 ;
    wire new_AGEMA_signal_35373 ;
    wire new_AGEMA_signal_35374 ;
    wire new_AGEMA_signal_35375 ;
    wire new_AGEMA_signal_35376 ;
    wire new_AGEMA_signal_35377 ;
    wire new_AGEMA_signal_35378 ;
    wire new_AGEMA_signal_35379 ;
    wire new_AGEMA_signal_35380 ;
    wire new_AGEMA_signal_35381 ;
    wire new_AGEMA_signal_35382 ;
    wire new_AGEMA_signal_35383 ;
    wire new_AGEMA_signal_35384 ;
    wire new_AGEMA_signal_35385 ;
    wire new_AGEMA_signal_35386 ;
    wire new_AGEMA_signal_35387 ;
    wire new_AGEMA_signal_35388 ;
    wire new_AGEMA_signal_35389 ;
    wire new_AGEMA_signal_35390 ;
    wire new_AGEMA_signal_35391 ;
    wire new_AGEMA_signal_35392 ;
    wire new_AGEMA_signal_35393 ;
    wire new_AGEMA_signal_35394 ;
    wire new_AGEMA_signal_35395 ;
    wire new_AGEMA_signal_35396 ;
    wire new_AGEMA_signal_35397 ;
    wire new_AGEMA_signal_35398 ;
    wire new_AGEMA_signal_35399 ;
    wire new_AGEMA_signal_35400 ;
    wire new_AGEMA_signal_35401 ;
    wire new_AGEMA_signal_35402 ;
    wire new_AGEMA_signal_35403 ;
    wire new_AGEMA_signal_35404 ;
    wire new_AGEMA_signal_35405 ;
    wire new_AGEMA_signal_35406 ;
    wire new_AGEMA_signal_35407 ;
    wire new_AGEMA_signal_35408 ;
    wire new_AGEMA_signal_35409 ;
    wire new_AGEMA_signal_35410 ;
    wire new_AGEMA_signal_35411 ;
    wire new_AGEMA_signal_35412 ;
    wire new_AGEMA_signal_35413 ;
    wire new_AGEMA_signal_35414 ;
    wire new_AGEMA_signal_35415 ;
    wire new_AGEMA_signal_35416 ;
    wire new_AGEMA_signal_35417 ;
    wire new_AGEMA_signal_35418 ;
    wire new_AGEMA_signal_35419 ;
    wire new_AGEMA_signal_35420 ;
    wire new_AGEMA_signal_35421 ;
    wire new_AGEMA_signal_35422 ;
    wire new_AGEMA_signal_35423 ;
    wire new_AGEMA_signal_35424 ;
    wire new_AGEMA_signal_35425 ;
    wire new_AGEMA_signal_35426 ;
    wire new_AGEMA_signal_35427 ;
    wire new_AGEMA_signal_35428 ;
    wire new_AGEMA_signal_35429 ;
    wire new_AGEMA_signal_35430 ;
    wire new_AGEMA_signal_35431 ;
    wire new_AGEMA_signal_35432 ;
    wire new_AGEMA_signal_35433 ;
    wire new_AGEMA_signal_35434 ;
    wire new_AGEMA_signal_35435 ;
    wire new_AGEMA_signal_35436 ;
    wire new_AGEMA_signal_35437 ;
    wire new_AGEMA_signal_35438 ;
    wire new_AGEMA_signal_35439 ;
    wire new_AGEMA_signal_35440 ;
    wire new_AGEMA_signal_35441 ;
    wire new_AGEMA_signal_35442 ;
    wire new_AGEMA_signal_35443 ;
    wire new_AGEMA_signal_35444 ;
    wire new_AGEMA_signal_35445 ;
    wire new_AGEMA_signal_35446 ;
    wire new_AGEMA_signal_35447 ;
    wire new_AGEMA_signal_35448 ;
    wire new_AGEMA_signal_35449 ;
    wire new_AGEMA_signal_35450 ;
    wire new_AGEMA_signal_35451 ;
    wire new_AGEMA_signal_35452 ;
    wire new_AGEMA_signal_35453 ;
    wire new_AGEMA_signal_35454 ;
    wire new_AGEMA_signal_35455 ;
    wire new_AGEMA_signal_35456 ;
    wire new_AGEMA_signal_35457 ;
    wire new_AGEMA_signal_35458 ;
    wire new_AGEMA_signal_35459 ;
    wire new_AGEMA_signal_35460 ;
    wire new_AGEMA_signal_35461 ;
    wire new_AGEMA_signal_35462 ;
    wire new_AGEMA_signal_35463 ;
    wire new_AGEMA_signal_35464 ;
    wire new_AGEMA_signal_35465 ;
    wire new_AGEMA_signal_35466 ;
    wire new_AGEMA_signal_35467 ;
    wire new_AGEMA_signal_35468 ;
    wire new_AGEMA_signal_35469 ;
    wire new_AGEMA_signal_35470 ;
    wire new_AGEMA_signal_35471 ;
    wire new_AGEMA_signal_35472 ;
    wire new_AGEMA_signal_35473 ;
    wire new_AGEMA_signal_35474 ;
    wire new_AGEMA_signal_35475 ;
    wire new_AGEMA_signal_35476 ;
    wire new_AGEMA_signal_35477 ;
    wire new_AGEMA_signal_35478 ;
    wire new_AGEMA_signal_35479 ;
    wire new_AGEMA_signal_35480 ;
    wire new_AGEMA_signal_35481 ;
    wire new_AGEMA_signal_35482 ;
    wire new_AGEMA_signal_35483 ;
    wire new_AGEMA_signal_35484 ;
    wire new_AGEMA_signal_35485 ;
    wire new_AGEMA_signal_35486 ;
    wire new_AGEMA_signal_35487 ;
    wire new_AGEMA_signal_35488 ;
    wire new_AGEMA_signal_35489 ;
    wire new_AGEMA_signal_35490 ;
    wire new_AGEMA_signal_35491 ;
    wire new_AGEMA_signal_35492 ;
    wire new_AGEMA_signal_35493 ;
    wire new_AGEMA_signal_35494 ;
    wire new_AGEMA_signal_35495 ;
    wire new_AGEMA_signal_35496 ;
    wire new_AGEMA_signal_35497 ;
    wire new_AGEMA_signal_35498 ;
    wire new_AGEMA_signal_35499 ;
    wire new_AGEMA_signal_35500 ;
    wire new_AGEMA_signal_35501 ;
    wire new_AGEMA_signal_35502 ;
    wire new_AGEMA_signal_35503 ;
    wire new_AGEMA_signal_35504 ;
    wire new_AGEMA_signal_35505 ;
    wire new_AGEMA_signal_35506 ;
    wire new_AGEMA_signal_35507 ;
    wire new_AGEMA_signal_35508 ;
    wire new_AGEMA_signal_35509 ;
    wire new_AGEMA_signal_35510 ;
    wire new_AGEMA_signal_35511 ;
    wire new_AGEMA_signal_35512 ;
    wire new_AGEMA_signal_35513 ;
    wire new_AGEMA_signal_35514 ;
    wire new_AGEMA_signal_35515 ;
    wire new_AGEMA_signal_35516 ;
    wire new_AGEMA_signal_35517 ;
    wire new_AGEMA_signal_35518 ;
    wire new_AGEMA_signal_35519 ;
    wire new_AGEMA_signal_35520 ;
    wire new_AGEMA_signal_35521 ;
    wire new_AGEMA_signal_35522 ;
    wire new_AGEMA_signal_35523 ;
    wire new_AGEMA_signal_35524 ;
    wire new_AGEMA_signal_35525 ;
    wire new_AGEMA_signal_35526 ;
    wire new_AGEMA_signal_35527 ;
    wire new_AGEMA_signal_35528 ;
    wire new_AGEMA_signal_35529 ;
    wire new_AGEMA_signal_35530 ;
    wire new_AGEMA_signal_35531 ;
    wire new_AGEMA_signal_35532 ;
    wire new_AGEMA_signal_35533 ;
    wire new_AGEMA_signal_35534 ;
    wire new_AGEMA_signal_35535 ;
    wire new_AGEMA_signal_35536 ;
    wire new_AGEMA_signal_35537 ;
    wire new_AGEMA_signal_35538 ;
    wire new_AGEMA_signal_35539 ;
    wire new_AGEMA_signal_35540 ;
    wire new_AGEMA_signal_35541 ;
    wire new_AGEMA_signal_35542 ;
    wire new_AGEMA_signal_35543 ;
    wire new_AGEMA_signal_35544 ;
    wire new_AGEMA_signal_35545 ;
    wire new_AGEMA_signal_35546 ;
    wire new_AGEMA_signal_35547 ;
    wire new_AGEMA_signal_35548 ;
    wire new_AGEMA_signal_35549 ;
    wire new_AGEMA_signal_35550 ;
    wire new_AGEMA_signal_35551 ;
    wire new_AGEMA_signal_35552 ;
    wire new_AGEMA_signal_35553 ;
    wire new_AGEMA_signal_35554 ;
    wire new_AGEMA_signal_35555 ;
    wire new_AGEMA_signal_35556 ;
    wire new_AGEMA_signal_35557 ;
    wire new_AGEMA_signal_35558 ;
    wire new_AGEMA_signal_35559 ;
    wire new_AGEMA_signal_35560 ;
    wire new_AGEMA_signal_35561 ;
    wire new_AGEMA_signal_35562 ;
    wire new_AGEMA_signal_35563 ;
    wire new_AGEMA_signal_35564 ;
    wire new_AGEMA_signal_35565 ;
    wire new_AGEMA_signal_35566 ;
    wire new_AGEMA_signal_35567 ;
    wire new_AGEMA_signal_35568 ;
    wire new_AGEMA_signal_35569 ;
    wire new_AGEMA_signal_35570 ;
    wire new_AGEMA_signal_35571 ;
    wire new_AGEMA_signal_35572 ;
    wire new_AGEMA_signal_35573 ;
    wire new_AGEMA_signal_35574 ;
    wire new_AGEMA_signal_35575 ;
    wire new_AGEMA_signal_35576 ;
    wire new_AGEMA_signal_35577 ;
    wire new_AGEMA_signal_35578 ;
    wire new_AGEMA_signal_35579 ;
    wire new_AGEMA_signal_35580 ;
    wire new_AGEMA_signal_35581 ;
    wire new_AGEMA_signal_35582 ;
    wire new_AGEMA_signal_35583 ;
    wire new_AGEMA_signal_35584 ;
    wire new_AGEMA_signal_35585 ;
    wire new_AGEMA_signal_35586 ;
    wire new_AGEMA_signal_35587 ;
    wire new_AGEMA_signal_35588 ;
    wire new_AGEMA_signal_35589 ;
    wire new_AGEMA_signal_35590 ;
    wire new_AGEMA_signal_35591 ;
    wire new_AGEMA_signal_35592 ;
    wire new_AGEMA_signal_35593 ;
    wire new_AGEMA_signal_35594 ;
    wire new_AGEMA_signal_35595 ;
    wire new_AGEMA_signal_35596 ;
    wire new_AGEMA_signal_35597 ;
    wire new_AGEMA_signal_35598 ;
    wire new_AGEMA_signal_35599 ;
    wire new_AGEMA_signal_35600 ;
    wire new_AGEMA_signal_35601 ;
    wire new_AGEMA_signal_35602 ;
    wire new_AGEMA_signal_35603 ;
    wire new_AGEMA_signal_35604 ;
    wire new_AGEMA_signal_35605 ;
    wire new_AGEMA_signal_35606 ;
    wire new_AGEMA_signal_35607 ;
    wire new_AGEMA_signal_35608 ;
    wire new_AGEMA_signal_35609 ;
    wire new_AGEMA_signal_35610 ;
    wire new_AGEMA_signal_35611 ;
    wire new_AGEMA_signal_35612 ;
    wire new_AGEMA_signal_35613 ;
    wire new_AGEMA_signal_35614 ;
    wire new_AGEMA_signal_35615 ;
    wire new_AGEMA_signal_35616 ;
    wire new_AGEMA_signal_35617 ;
    wire new_AGEMA_signal_35618 ;
    wire new_AGEMA_signal_35619 ;
    wire new_AGEMA_signal_35620 ;
    wire new_AGEMA_signal_35621 ;
    wire new_AGEMA_signal_35622 ;
    wire new_AGEMA_signal_35623 ;
    wire new_AGEMA_signal_35624 ;
    wire new_AGEMA_signal_35625 ;
    wire new_AGEMA_signal_35626 ;
    wire new_AGEMA_signal_35627 ;
    wire new_AGEMA_signal_35628 ;
    wire new_AGEMA_signal_35629 ;
    wire new_AGEMA_signal_35630 ;
    wire new_AGEMA_signal_35631 ;
    wire new_AGEMA_signal_35632 ;
    wire new_AGEMA_signal_35633 ;
    wire new_AGEMA_signal_35634 ;
    wire new_AGEMA_signal_35635 ;
    wire new_AGEMA_signal_35636 ;
    wire new_AGEMA_signal_35637 ;
    wire new_AGEMA_signal_35638 ;
    wire new_AGEMA_signal_35639 ;
    wire new_AGEMA_signal_35640 ;
    wire new_AGEMA_signal_35641 ;
    wire new_AGEMA_signal_35642 ;
    wire new_AGEMA_signal_35643 ;
    wire new_AGEMA_signal_35644 ;
    wire new_AGEMA_signal_35645 ;
    wire new_AGEMA_signal_35646 ;
    wire new_AGEMA_signal_35647 ;
    wire new_AGEMA_signal_35648 ;
    wire new_AGEMA_signal_35649 ;
    wire new_AGEMA_signal_35650 ;
    wire new_AGEMA_signal_35651 ;
    wire new_AGEMA_signal_35652 ;
    wire new_AGEMA_signal_35653 ;
    wire new_AGEMA_signal_35654 ;
    wire new_AGEMA_signal_35655 ;
    wire new_AGEMA_signal_35656 ;
    wire new_AGEMA_signal_35657 ;
    wire new_AGEMA_signal_35658 ;
    wire new_AGEMA_signal_35659 ;
    wire new_AGEMA_signal_35660 ;
    wire new_AGEMA_signal_35661 ;
    wire new_AGEMA_signal_35662 ;
    wire new_AGEMA_signal_35663 ;
    wire new_AGEMA_signal_35664 ;
    wire new_AGEMA_signal_35665 ;
    wire new_AGEMA_signal_35666 ;
    wire new_AGEMA_signal_35667 ;
    wire new_AGEMA_signal_35668 ;
    wire new_AGEMA_signal_35669 ;
    wire new_AGEMA_signal_35670 ;
    wire new_AGEMA_signal_35671 ;
    wire new_AGEMA_signal_35672 ;
    wire new_AGEMA_signal_35673 ;
    wire new_AGEMA_signal_35674 ;
    wire new_AGEMA_signal_35675 ;
    wire new_AGEMA_signal_35676 ;
    wire new_AGEMA_signal_35677 ;
    wire new_AGEMA_signal_35678 ;
    wire new_AGEMA_signal_35679 ;
    wire new_AGEMA_signal_35680 ;
    wire new_AGEMA_signal_35681 ;
    wire new_AGEMA_signal_35682 ;
    wire new_AGEMA_signal_35683 ;
    wire new_AGEMA_signal_35684 ;
    wire new_AGEMA_signal_35685 ;
    wire new_AGEMA_signal_35686 ;
    wire new_AGEMA_signal_35687 ;
    wire new_AGEMA_signal_35688 ;
    wire new_AGEMA_signal_35689 ;
    wire new_AGEMA_signal_35690 ;
    wire new_AGEMA_signal_35691 ;
    wire new_AGEMA_signal_35692 ;
    wire new_AGEMA_signal_35693 ;
    wire new_AGEMA_signal_35694 ;
    wire new_AGEMA_signal_35695 ;
    wire new_AGEMA_signal_35696 ;
    wire new_AGEMA_signal_35697 ;
    wire new_AGEMA_signal_35698 ;
    wire new_AGEMA_signal_35699 ;
    wire new_AGEMA_signal_35700 ;
    wire new_AGEMA_signal_35701 ;
    wire new_AGEMA_signal_35702 ;
    wire new_AGEMA_signal_35703 ;
    wire new_AGEMA_signal_35704 ;
    wire new_AGEMA_signal_35705 ;
    wire new_AGEMA_signal_35706 ;
    wire new_AGEMA_signal_35707 ;
    wire new_AGEMA_signal_35708 ;
    wire new_AGEMA_signal_35709 ;
    wire new_AGEMA_signal_35710 ;
    wire new_AGEMA_signal_35711 ;
    wire new_AGEMA_signal_35712 ;
    wire new_AGEMA_signal_35713 ;
    wire new_AGEMA_signal_35714 ;
    wire new_AGEMA_signal_35715 ;
    wire new_AGEMA_signal_35716 ;
    wire new_AGEMA_signal_35717 ;
    wire new_AGEMA_signal_35718 ;
    wire new_AGEMA_signal_35719 ;
    wire new_AGEMA_signal_35720 ;
    wire new_AGEMA_signal_35721 ;
    wire new_AGEMA_signal_35722 ;
    wire new_AGEMA_signal_35723 ;
    wire new_AGEMA_signal_35724 ;
    wire new_AGEMA_signal_35725 ;
    wire new_AGEMA_signal_35726 ;
    wire new_AGEMA_signal_35727 ;
    wire new_AGEMA_signal_35728 ;
    wire new_AGEMA_signal_35729 ;
    wire new_AGEMA_signal_35730 ;
    wire new_AGEMA_signal_35731 ;
    wire new_AGEMA_signal_35732 ;
    wire new_AGEMA_signal_35733 ;
    wire new_AGEMA_signal_35734 ;
    wire new_AGEMA_signal_35735 ;
    wire new_AGEMA_signal_35736 ;
    wire new_AGEMA_signal_35737 ;
    wire new_AGEMA_signal_35738 ;
    wire new_AGEMA_signal_35739 ;
    wire new_AGEMA_signal_35740 ;
    wire new_AGEMA_signal_35741 ;
    wire new_AGEMA_signal_35742 ;
    wire new_AGEMA_signal_35743 ;
    wire new_AGEMA_signal_35744 ;
    wire new_AGEMA_signal_35745 ;
    wire new_AGEMA_signal_35746 ;
    wire new_AGEMA_signal_35747 ;
    wire new_AGEMA_signal_35748 ;
    wire new_AGEMA_signal_35749 ;
    wire new_AGEMA_signal_35750 ;
    wire new_AGEMA_signal_35751 ;
    wire new_AGEMA_signal_35752 ;
    wire new_AGEMA_signal_35753 ;
    wire new_AGEMA_signal_35754 ;
    wire new_AGEMA_signal_35755 ;
    wire new_AGEMA_signal_35756 ;
    wire new_AGEMA_signal_35757 ;
    wire new_AGEMA_signal_35758 ;
    wire new_AGEMA_signal_35759 ;
    wire new_AGEMA_signal_35760 ;
    wire new_AGEMA_signal_35761 ;
    wire new_AGEMA_signal_35762 ;
    wire new_AGEMA_signal_35763 ;
    wire new_AGEMA_signal_35764 ;
    wire new_AGEMA_signal_35765 ;
    wire new_AGEMA_signal_35766 ;
    wire new_AGEMA_signal_35767 ;
    wire new_AGEMA_signal_35768 ;
    wire new_AGEMA_signal_35769 ;
    wire new_AGEMA_signal_35770 ;
    wire new_AGEMA_signal_35771 ;
    wire new_AGEMA_signal_35772 ;
    wire new_AGEMA_signal_35773 ;
    wire new_AGEMA_signal_35774 ;
    wire new_AGEMA_signal_35775 ;
    wire new_AGEMA_signal_35776 ;
    wire new_AGEMA_signal_35777 ;
    wire new_AGEMA_signal_35778 ;
    wire new_AGEMA_signal_35779 ;
    wire new_AGEMA_signal_35780 ;
    wire new_AGEMA_signal_35781 ;
    wire new_AGEMA_signal_35782 ;
    wire new_AGEMA_signal_35783 ;
    wire new_AGEMA_signal_35784 ;
    wire new_AGEMA_signal_35785 ;
    wire new_AGEMA_signal_35786 ;
    wire new_AGEMA_signal_35787 ;
    wire new_AGEMA_signal_35788 ;
    wire new_AGEMA_signal_35789 ;
    wire new_AGEMA_signal_35790 ;
    wire new_AGEMA_signal_35791 ;
    wire new_AGEMA_signal_35792 ;
    wire new_AGEMA_signal_35793 ;
    wire new_AGEMA_signal_35794 ;
    wire new_AGEMA_signal_35795 ;
    wire new_AGEMA_signal_35796 ;
    wire new_AGEMA_signal_35797 ;
    wire new_AGEMA_signal_35798 ;
    wire new_AGEMA_signal_35799 ;
    wire new_AGEMA_signal_35800 ;
    wire new_AGEMA_signal_35801 ;
    wire new_AGEMA_signal_35802 ;
    wire new_AGEMA_signal_35803 ;
    wire new_AGEMA_signal_35804 ;
    wire new_AGEMA_signal_35805 ;
    wire new_AGEMA_signal_35806 ;
    wire new_AGEMA_signal_35807 ;
    wire new_AGEMA_signal_35808 ;
    wire new_AGEMA_signal_35809 ;
    wire new_AGEMA_signal_35810 ;
    wire new_AGEMA_signal_35811 ;
    wire new_AGEMA_signal_35812 ;
    wire new_AGEMA_signal_35813 ;
    wire new_AGEMA_signal_35814 ;
    wire new_AGEMA_signal_35815 ;
    wire new_AGEMA_signal_35816 ;
    wire new_AGEMA_signal_35817 ;
    wire new_AGEMA_signal_35818 ;
    wire new_AGEMA_signal_35819 ;
    wire new_AGEMA_signal_35820 ;
    wire new_AGEMA_signal_35821 ;
    wire new_AGEMA_signal_35822 ;
    wire new_AGEMA_signal_35823 ;
    wire new_AGEMA_signal_35824 ;
    wire new_AGEMA_signal_35825 ;
    wire new_AGEMA_signal_35826 ;
    wire new_AGEMA_signal_35827 ;
    wire new_AGEMA_signal_35828 ;
    wire new_AGEMA_signal_35829 ;
    wire new_AGEMA_signal_35830 ;
    wire new_AGEMA_signal_35831 ;
    wire new_AGEMA_signal_35832 ;
    wire new_AGEMA_signal_35833 ;
    wire new_AGEMA_signal_35834 ;
    wire new_AGEMA_signal_35835 ;
    wire new_AGEMA_signal_35836 ;
    wire new_AGEMA_signal_35837 ;
    wire new_AGEMA_signal_35838 ;
    wire new_AGEMA_signal_35839 ;
    wire new_AGEMA_signal_35840 ;
    wire new_AGEMA_signal_35841 ;
    wire new_AGEMA_signal_35842 ;
    wire new_AGEMA_signal_35843 ;
    wire new_AGEMA_signal_35844 ;
    wire new_AGEMA_signal_35845 ;
    wire new_AGEMA_signal_35846 ;
    wire new_AGEMA_signal_35847 ;
    wire new_AGEMA_signal_35848 ;
    wire new_AGEMA_signal_35849 ;
    wire new_AGEMA_signal_35850 ;
    wire new_AGEMA_signal_35851 ;
    wire new_AGEMA_signal_35852 ;
    wire new_AGEMA_signal_35853 ;
    wire new_AGEMA_signal_35854 ;
    wire new_AGEMA_signal_35855 ;
    wire new_AGEMA_signal_35856 ;
    wire new_AGEMA_signal_35857 ;
    wire new_AGEMA_signal_35858 ;
    wire new_AGEMA_signal_35859 ;
    wire new_AGEMA_signal_35860 ;
    wire new_AGEMA_signal_35861 ;
    wire new_AGEMA_signal_35862 ;
    wire new_AGEMA_signal_35863 ;
    wire new_AGEMA_signal_35864 ;
    wire new_AGEMA_signal_35865 ;
    wire new_AGEMA_signal_35866 ;
    wire new_AGEMA_signal_35867 ;
    wire new_AGEMA_signal_35868 ;
    wire new_AGEMA_signal_35869 ;
    wire new_AGEMA_signal_35870 ;
    wire new_AGEMA_signal_35871 ;
    wire new_AGEMA_signal_35872 ;
    wire new_AGEMA_signal_35873 ;
    wire new_AGEMA_signal_35874 ;
    wire new_AGEMA_signal_35875 ;
    wire new_AGEMA_signal_35876 ;
    wire new_AGEMA_signal_35877 ;
    wire new_AGEMA_signal_35878 ;
    wire new_AGEMA_signal_35879 ;
    wire new_AGEMA_signal_35880 ;
    wire new_AGEMA_signal_35881 ;
    wire new_AGEMA_signal_35882 ;
    wire new_AGEMA_signal_35883 ;
    wire new_AGEMA_signal_35884 ;
    wire new_AGEMA_signal_35885 ;
    wire new_AGEMA_signal_35886 ;
    wire new_AGEMA_signal_35887 ;
    wire new_AGEMA_signal_35888 ;
    wire new_AGEMA_signal_35889 ;
    wire new_AGEMA_signal_35890 ;
    wire new_AGEMA_signal_35891 ;
    wire new_AGEMA_signal_35892 ;
    wire new_AGEMA_signal_35893 ;
    wire new_AGEMA_signal_35894 ;
    wire new_AGEMA_signal_35895 ;
    wire new_AGEMA_signal_35896 ;
    wire new_AGEMA_signal_35897 ;
    wire new_AGEMA_signal_35898 ;
    wire new_AGEMA_signal_35899 ;
    wire new_AGEMA_signal_35900 ;
    wire new_AGEMA_signal_35901 ;
    wire new_AGEMA_signal_35902 ;
    wire new_AGEMA_signal_35903 ;
    wire new_AGEMA_signal_35904 ;
    wire new_AGEMA_signal_35905 ;
    wire new_AGEMA_signal_35906 ;
    wire new_AGEMA_signal_35907 ;
    wire new_AGEMA_signal_35908 ;
    wire new_AGEMA_signal_35909 ;
    wire new_AGEMA_signal_35910 ;
    wire new_AGEMA_signal_35911 ;
    wire new_AGEMA_signal_35912 ;
    wire new_AGEMA_signal_35913 ;
    wire new_AGEMA_signal_35914 ;
    wire new_AGEMA_signal_35915 ;
    wire new_AGEMA_signal_35916 ;
    wire new_AGEMA_signal_35917 ;
    wire new_AGEMA_signal_35918 ;
    wire new_AGEMA_signal_35919 ;
    wire new_AGEMA_signal_35920 ;
    wire new_AGEMA_signal_35921 ;
    wire new_AGEMA_signal_35922 ;
    wire new_AGEMA_signal_35923 ;
    wire new_AGEMA_signal_35924 ;
    wire new_AGEMA_signal_35925 ;
    wire new_AGEMA_signal_35926 ;
    wire new_AGEMA_signal_35927 ;
    wire new_AGEMA_signal_35928 ;
    wire new_AGEMA_signal_35929 ;
    wire new_AGEMA_signal_35930 ;
    wire new_AGEMA_signal_35931 ;
    wire new_AGEMA_signal_35932 ;
    wire new_AGEMA_signal_35933 ;
    wire new_AGEMA_signal_35934 ;
    wire new_AGEMA_signal_35935 ;
    wire new_AGEMA_signal_35936 ;
    wire new_AGEMA_signal_35937 ;
    wire new_AGEMA_signal_35938 ;
    wire new_AGEMA_signal_35939 ;
    wire new_AGEMA_signal_35940 ;
    wire new_AGEMA_signal_35941 ;
    wire new_AGEMA_signal_35942 ;
    wire new_AGEMA_signal_35943 ;
    wire new_AGEMA_signal_35944 ;
    wire new_AGEMA_signal_35945 ;
    wire new_AGEMA_signal_35946 ;
    wire new_AGEMA_signal_35947 ;
    wire new_AGEMA_signal_35948 ;
    wire new_AGEMA_signal_35949 ;
    wire new_AGEMA_signal_35950 ;
    wire new_AGEMA_signal_35951 ;
    wire new_AGEMA_signal_35952 ;
    wire new_AGEMA_signal_35953 ;
    wire new_AGEMA_signal_35954 ;
    wire new_AGEMA_signal_35955 ;
    wire new_AGEMA_signal_35956 ;
    wire new_AGEMA_signal_35957 ;
    wire new_AGEMA_signal_35958 ;
    wire new_AGEMA_signal_35959 ;
    wire new_AGEMA_signal_35960 ;
    wire new_AGEMA_signal_35961 ;
    wire new_AGEMA_signal_35962 ;
    wire new_AGEMA_signal_35963 ;
    wire new_AGEMA_signal_35964 ;
    wire new_AGEMA_signal_35965 ;
    wire new_AGEMA_signal_35966 ;
    wire new_AGEMA_signal_35967 ;
    wire new_AGEMA_signal_35968 ;
    wire new_AGEMA_signal_35969 ;
    wire new_AGEMA_signal_35970 ;
    wire new_AGEMA_signal_35971 ;
    wire new_AGEMA_signal_35972 ;
    wire new_AGEMA_signal_35973 ;
    wire new_AGEMA_signal_35974 ;
    wire new_AGEMA_signal_35975 ;
    wire new_AGEMA_signal_35976 ;
    wire new_AGEMA_signal_35977 ;
    wire new_AGEMA_signal_35978 ;
    wire new_AGEMA_signal_35979 ;
    wire new_AGEMA_signal_35980 ;
    wire new_AGEMA_signal_35981 ;
    wire new_AGEMA_signal_35982 ;
    wire new_AGEMA_signal_35983 ;
    wire new_AGEMA_signal_35984 ;
    wire new_AGEMA_signal_35985 ;
    wire new_AGEMA_signal_35986 ;
    wire new_AGEMA_signal_35987 ;
    wire new_AGEMA_signal_35988 ;
    wire new_AGEMA_signal_35989 ;
    wire new_AGEMA_signal_35990 ;
    wire new_AGEMA_signal_35991 ;
    wire new_AGEMA_signal_35992 ;
    wire new_AGEMA_signal_35993 ;
    wire new_AGEMA_signal_35994 ;
    wire new_AGEMA_signal_35995 ;
    wire new_AGEMA_signal_35996 ;
    wire new_AGEMA_signal_35997 ;
    wire new_AGEMA_signal_35998 ;
    wire new_AGEMA_signal_35999 ;
    wire new_AGEMA_signal_36000 ;
    wire new_AGEMA_signal_36001 ;
    wire new_AGEMA_signal_36002 ;
    wire new_AGEMA_signal_36003 ;
    wire new_AGEMA_signal_36004 ;
    wire new_AGEMA_signal_36005 ;
    wire new_AGEMA_signal_36006 ;
    wire new_AGEMA_signal_36007 ;
    wire new_AGEMA_signal_36008 ;
    wire new_AGEMA_signal_36009 ;
    wire new_AGEMA_signal_36010 ;
    wire new_AGEMA_signal_36011 ;
    wire new_AGEMA_signal_36012 ;
    wire new_AGEMA_signal_36013 ;
    wire new_AGEMA_signal_36014 ;
    wire new_AGEMA_signal_36015 ;
    wire new_AGEMA_signal_36016 ;
    wire new_AGEMA_signal_36017 ;
    wire new_AGEMA_signal_36018 ;
    wire new_AGEMA_signal_36019 ;
    wire new_AGEMA_signal_36020 ;
    wire new_AGEMA_signal_36021 ;
    wire new_AGEMA_signal_36022 ;
    wire new_AGEMA_signal_36023 ;
    wire new_AGEMA_signal_36024 ;
    wire new_AGEMA_signal_36025 ;
    wire new_AGEMA_signal_36026 ;
    wire new_AGEMA_signal_36027 ;
    wire new_AGEMA_signal_36028 ;
    wire new_AGEMA_signal_36029 ;
    wire new_AGEMA_signal_36030 ;
    wire new_AGEMA_signal_36031 ;
    wire new_AGEMA_signal_36032 ;
    wire new_AGEMA_signal_36033 ;
    wire new_AGEMA_signal_36034 ;
    wire new_AGEMA_signal_36035 ;
    wire new_AGEMA_signal_36036 ;
    wire new_AGEMA_signal_36037 ;
    wire new_AGEMA_signal_36038 ;
    wire new_AGEMA_signal_36039 ;
    wire new_AGEMA_signal_36040 ;
    wire new_AGEMA_signal_36041 ;
    wire new_AGEMA_signal_36042 ;
    wire new_AGEMA_signal_36043 ;
    wire new_AGEMA_signal_36044 ;
    wire new_AGEMA_signal_36045 ;
    wire new_AGEMA_signal_36046 ;
    wire new_AGEMA_signal_36047 ;
    wire new_AGEMA_signal_36048 ;
    wire new_AGEMA_signal_36049 ;
    wire new_AGEMA_signal_36050 ;
    wire new_AGEMA_signal_36051 ;
    wire new_AGEMA_signal_36052 ;
    wire new_AGEMA_signal_36053 ;
    wire new_AGEMA_signal_36054 ;
    wire new_AGEMA_signal_36055 ;
    wire new_AGEMA_signal_36056 ;
    wire new_AGEMA_signal_36057 ;
    wire new_AGEMA_signal_36058 ;
    wire new_AGEMA_signal_36059 ;
    wire new_AGEMA_signal_36060 ;
    wire new_AGEMA_signal_36061 ;
    wire new_AGEMA_signal_36062 ;
    wire new_AGEMA_signal_36063 ;
    wire new_AGEMA_signal_36064 ;
    wire new_AGEMA_signal_36065 ;
    wire new_AGEMA_signal_36066 ;
    wire new_AGEMA_signal_36067 ;
    wire new_AGEMA_signal_36068 ;
    wire new_AGEMA_signal_36069 ;
    wire new_AGEMA_signal_36070 ;
    wire new_AGEMA_signal_36071 ;
    wire new_AGEMA_signal_36072 ;
    wire new_AGEMA_signal_36073 ;
    wire new_AGEMA_signal_36074 ;
    wire new_AGEMA_signal_36075 ;
    wire new_AGEMA_signal_36076 ;
    wire new_AGEMA_signal_36077 ;
    wire new_AGEMA_signal_36078 ;
    wire new_AGEMA_signal_36079 ;
    wire new_AGEMA_signal_36080 ;
    wire new_AGEMA_signal_36081 ;
    wire new_AGEMA_signal_36082 ;
    wire new_AGEMA_signal_36083 ;
    wire new_AGEMA_signal_36084 ;
    wire new_AGEMA_signal_36085 ;
    wire new_AGEMA_signal_36086 ;
    wire new_AGEMA_signal_36087 ;
    wire new_AGEMA_signal_36088 ;
    wire new_AGEMA_signal_36089 ;
    wire new_AGEMA_signal_36090 ;
    wire new_AGEMA_signal_36091 ;
    wire new_AGEMA_signal_36092 ;
    wire new_AGEMA_signal_36093 ;
    wire new_AGEMA_signal_36094 ;
    wire new_AGEMA_signal_36095 ;
    wire new_AGEMA_signal_36096 ;
    wire new_AGEMA_signal_36097 ;
    wire new_AGEMA_signal_36098 ;
    wire new_AGEMA_signal_36099 ;
    wire new_AGEMA_signal_36100 ;
    wire new_AGEMA_signal_36101 ;
    wire new_AGEMA_signal_36102 ;
    wire new_AGEMA_signal_36103 ;
    wire new_AGEMA_signal_36104 ;
    wire new_AGEMA_signal_36105 ;
    wire new_AGEMA_signal_36106 ;
    wire new_AGEMA_signal_36107 ;
    wire new_AGEMA_signal_36108 ;
    wire new_AGEMA_signal_36109 ;
    wire new_AGEMA_signal_36110 ;
    wire new_AGEMA_signal_36111 ;
    wire new_AGEMA_signal_36112 ;
    wire new_AGEMA_signal_36113 ;
    wire new_AGEMA_signal_36114 ;
    wire new_AGEMA_signal_36115 ;
    wire new_AGEMA_signal_36116 ;
    wire new_AGEMA_signal_36117 ;
    wire new_AGEMA_signal_36118 ;
    wire new_AGEMA_signal_36119 ;
    wire new_AGEMA_signal_36120 ;
    wire new_AGEMA_signal_36121 ;
    wire new_AGEMA_signal_36122 ;
    wire new_AGEMA_signal_36123 ;
    wire new_AGEMA_signal_36124 ;
    wire new_AGEMA_signal_36125 ;
    wire new_AGEMA_signal_36126 ;
    wire new_AGEMA_signal_36127 ;
    wire new_AGEMA_signal_36128 ;
    wire new_AGEMA_signal_36129 ;
    wire new_AGEMA_signal_36130 ;
    wire new_AGEMA_signal_36131 ;
    wire new_AGEMA_signal_36132 ;
    wire new_AGEMA_signal_36133 ;
    wire new_AGEMA_signal_36134 ;
    wire new_AGEMA_signal_36135 ;
    wire new_AGEMA_signal_36136 ;
    wire new_AGEMA_signal_36137 ;
    wire new_AGEMA_signal_36138 ;
    wire new_AGEMA_signal_36139 ;
    wire new_AGEMA_signal_36140 ;
    wire new_AGEMA_signal_36141 ;
    wire new_AGEMA_signal_36142 ;
    wire new_AGEMA_signal_36143 ;
    wire new_AGEMA_signal_36144 ;
    wire new_AGEMA_signal_36145 ;
    wire new_AGEMA_signal_36146 ;
    wire new_AGEMA_signal_36147 ;
    wire new_AGEMA_signal_36148 ;
    wire new_AGEMA_signal_36149 ;
    wire new_AGEMA_signal_36150 ;
    wire new_AGEMA_signal_36151 ;
    wire new_AGEMA_signal_36152 ;
    wire new_AGEMA_signal_36153 ;
    wire new_AGEMA_signal_36154 ;
    wire new_AGEMA_signal_36155 ;
    wire new_AGEMA_signal_36156 ;
    wire new_AGEMA_signal_36157 ;
    wire new_AGEMA_signal_36158 ;
    wire new_AGEMA_signal_36159 ;
    wire new_AGEMA_signal_36160 ;
    wire new_AGEMA_signal_36161 ;
    wire new_AGEMA_signal_36162 ;
    wire new_AGEMA_signal_36163 ;
    wire new_AGEMA_signal_36164 ;
    wire new_AGEMA_signal_36165 ;
    wire new_AGEMA_signal_36166 ;
    wire new_AGEMA_signal_36167 ;
    wire new_AGEMA_signal_36168 ;
    wire new_AGEMA_signal_36169 ;
    wire new_AGEMA_signal_36170 ;
    wire new_AGEMA_signal_36171 ;
    wire new_AGEMA_signal_36172 ;
    wire new_AGEMA_signal_36173 ;
    wire new_AGEMA_signal_36174 ;
    wire new_AGEMA_signal_36175 ;
    wire new_AGEMA_signal_36176 ;
    wire new_AGEMA_signal_36177 ;
    wire new_AGEMA_signal_36178 ;
    wire new_AGEMA_signal_36179 ;
    wire new_AGEMA_signal_36180 ;
    wire new_AGEMA_signal_36181 ;
    wire new_AGEMA_signal_36182 ;
    wire new_AGEMA_signal_36183 ;
    wire new_AGEMA_signal_36184 ;
    wire new_AGEMA_signal_36185 ;
    wire new_AGEMA_signal_36186 ;
    wire new_AGEMA_signal_36187 ;
    wire new_AGEMA_signal_36188 ;
    wire new_AGEMA_signal_36189 ;
    wire new_AGEMA_signal_36190 ;
    wire new_AGEMA_signal_36191 ;
    wire new_AGEMA_signal_36192 ;
    wire new_AGEMA_signal_36193 ;
    wire new_AGEMA_signal_36194 ;
    wire new_AGEMA_signal_36195 ;
    wire new_AGEMA_signal_36196 ;
    wire new_AGEMA_signal_36197 ;
    wire new_AGEMA_signal_36198 ;
    wire new_AGEMA_signal_36199 ;
    wire new_AGEMA_signal_36200 ;
    wire new_AGEMA_signal_36201 ;
    wire new_AGEMA_signal_36202 ;
    wire new_AGEMA_signal_36203 ;
    wire new_AGEMA_signal_36204 ;
    wire new_AGEMA_signal_36205 ;
    wire new_AGEMA_signal_36206 ;
    wire new_AGEMA_signal_36207 ;
    wire new_AGEMA_signal_36208 ;
    wire new_AGEMA_signal_36209 ;
    wire new_AGEMA_signal_36210 ;
    wire new_AGEMA_signal_36211 ;
    wire new_AGEMA_signal_36212 ;
    wire new_AGEMA_signal_36213 ;
    wire new_AGEMA_signal_36214 ;
    wire new_AGEMA_signal_36215 ;
    wire new_AGEMA_signal_36216 ;
    wire new_AGEMA_signal_36217 ;
    wire new_AGEMA_signal_36218 ;
    wire new_AGEMA_signal_36219 ;
    wire new_AGEMA_signal_36220 ;
    wire new_AGEMA_signal_36221 ;
    wire new_AGEMA_signal_36222 ;
    wire new_AGEMA_signal_36223 ;
    wire new_AGEMA_signal_36224 ;
    wire new_AGEMA_signal_36225 ;
    wire new_AGEMA_signal_36226 ;
    wire new_AGEMA_signal_36227 ;
    wire new_AGEMA_signal_36228 ;
    wire new_AGEMA_signal_36229 ;
    wire new_AGEMA_signal_36230 ;
    wire new_AGEMA_signal_36231 ;
    wire new_AGEMA_signal_36232 ;
    wire new_AGEMA_signal_36233 ;
    wire new_AGEMA_signal_36234 ;
    wire new_AGEMA_signal_36235 ;
    wire new_AGEMA_signal_36236 ;
    wire new_AGEMA_signal_36237 ;
    wire new_AGEMA_signal_36238 ;
    wire new_AGEMA_signal_36239 ;
    wire new_AGEMA_signal_36240 ;
    wire new_AGEMA_signal_36241 ;
    wire new_AGEMA_signal_36242 ;
    wire new_AGEMA_signal_36243 ;
    wire new_AGEMA_signal_36244 ;
    wire new_AGEMA_signal_36245 ;
    wire new_AGEMA_signal_36246 ;
    wire new_AGEMA_signal_36247 ;
    wire new_AGEMA_signal_36248 ;
    wire new_AGEMA_signal_36249 ;
    wire new_AGEMA_signal_36250 ;
    wire new_AGEMA_signal_36251 ;
    wire new_AGEMA_signal_36252 ;
    wire new_AGEMA_signal_36253 ;
    wire new_AGEMA_signal_36254 ;
    wire new_AGEMA_signal_36255 ;
    wire new_AGEMA_signal_36256 ;
    wire new_AGEMA_signal_36257 ;
    wire new_AGEMA_signal_36258 ;
    wire new_AGEMA_signal_36259 ;
    wire new_AGEMA_signal_36260 ;
    wire new_AGEMA_signal_36261 ;
    wire new_AGEMA_signal_36262 ;
    wire new_AGEMA_signal_36263 ;
    wire new_AGEMA_signal_36264 ;
    wire new_AGEMA_signal_36265 ;
    wire new_AGEMA_signal_36266 ;
    wire new_AGEMA_signal_36267 ;
    wire new_AGEMA_signal_36268 ;
    wire new_AGEMA_signal_36269 ;
    wire new_AGEMA_signal_36270 ;
    wire new_AGEMA_signal_36271 ;
    wire new_AGEMA_signal_36272 ;
    wire new_AGEMA_signal_36273 ;
    wire new_AGEMA_signal_36274 ;
    wire new_AGEMA_signal_36275 ;
    wire new_AGEMA_signal_36276 ;
    wire new_AGEMA_signal_36277 ;
    wire new_AGEMA_signal_36278 ;
    wire new_AGEMA_signal_36279 ;
    wire new_AGEMA_signal_36280 ;
    wire new_AGEMA_signal_36281 ;
    wire new_AGEMA_signal_36282 ;
    wire new_AGEMA_signal_36283 ;
    wire new_AGEMA_signal_36284 ;
    wire new_AGEMA_signal_36285 ;
    wire new_AGEMA_signal_36286 ;
    wire new_AGEMA_signal_36287 ;
    wire new_AGEMA_signal_36288 ;
    wire new_AGEMA_signal_36289 ;
    wire new_AGEMA_signal_36290 ;
    wire new_AGEMA_signal_36291 ;
    wire new_AGEMA_signal_36292 ;
    wire new_AGEMA_signal_36293 ;
    wire new_AGEMA_signal_36294 ;
    wire new_AGEMA_signal_36295 ;
    wire new_AGEMA_signal_36296 ;
    wire new_AGEMA_signal_36297 ;
    wire new_AGEMA_signal_36298 ;
    wire new_AGEMA_signal_36299 ;
    wire new_AGEMA_signal_36300 ;
    wire new_AGEMA_signal_36301 ;
    wire new_AGEMA_signal_36302 ;
    wire new_AGEMA_signal_36303 ;
    wire new_AGEMA_signal_36304 ;
    wire new_AGEMA_signal_36305 ;
    wire new_AGEMA_signal_36306 ;
    wire new_AGEMA_signal_36307 ;
    wire new_AGEMA_signal_36308 ;
    wire new_AGEMA_signal_36309 ;
    wire new_AGEMA_signal_36310 ;
    wire new_AGEMA_signal_36311 ;
    wire new_AGEMA_signal_36312 ;
    wire new_AGEMA_signal_36313 ;
    wire new_AGEMA_signal_36314 ;
    wire new_AGEMA_signal_36315 ;
    wire new_AGEMA_signal_36316 ;
    wire new_AGEMA_signal_36317 ;
    wire new_AGEMA_signal_36318 ;
    wire new_AGEMA_signal_36319 ;
    wire new_AGEMA_signal_36320 ;
    wire new_AGEMA_signal_36321 ;
    wire new_AGEMA_signal_36322 ;
    wire new_AGEMA_signal_36323 ;
    wire new_AGEMA_signal_36324 ;
    wire new_AGEMA_signal_36325 ;
    wire new_AGEMA_signal_36326 ;
    wire new_AGEMA_signal_36327 ;
    wire new_AGEMA_signal_36328 ;
    wire new_AGEMA_signal_36329 ;
    wire new_AGEMA_signal_36330 ;
    wire new_AGEMA_signal_36331 ;
    wire new_AGEMA_signal_36332 ;
    wire new_AGEMA_signal_36333 ;
    wire new_AGEMA_signal_36334 ;
    wire new_AGEMA_signal_36335 ;
    wire new_AGEMA_signal_36336 ;
    wire new_AGEMA_signal_36337 ;
    wire new_AGEMA_signal_36338 ;
    wire new_AGEMA_signal_36339 ;
    wire new_AGEMA_signal_36340 ;
    wire new_AGEMA_signal_36341 ;
    wire new_AGEMA_signal_36342 ;
    wire new_AGEMA_signal_36343 ;
    wire new_AGEMA_signal_36344 ;
    wire new_AGEMA_signal_36345 ;
    wire new_AGEMA_signal_36346 ;
    wire new_AGEMA_signal_36347 ;
    wire new_AGEMA_signal_36348 ;
    wire new_AGEMA_signal_36349 ;
    wire new_AGEMA_signal_36350 ;
    wire new_AGEMA_signal_36351 ;
    wire new_AGEMA_signal_36352 ;
    wire new_AGEMA_signal_36353 ;
    wire new_AGEMA_signal_36354 ;
    wire new_AGEMA_signal_36355 ;
    wire new_AGEMA_signal_36356 ;
    wire new_AGEMA_signal_36357 ;
    wire new_AGEMA_signal_36358 ;
    wire new_AGEMA_signal_36359 ;
    wire new_AGEMA_signal_36360 ;
    wire new_AGEMA_signal_36361 ;
    wire new_AGEMA_signal_36362 ;
    wire new_AGEMA_signal_36363 ;
    wire new_AGEMA_signal_36364 ;
    wire new_AGEMA_signal_36365 ;
    wire new_AGEMA_signal_36366 ;
    wire new_AGEMA_signal_36367 ;
    wire new_AGEMA_signal_36368 ;
    wire new_AGEMA_signal_36369 ;
    wire new_AGEMA_signal_36370 ;
    wire new_AGEMA_signal_36371 ;
    wire new_AGEMA_signal_36372 ;
    wire new_AGEMA_signal_36373 ;
    wire new_AGEMA_signal_36374 ;
    wire new_AGEMA_signal_36375 ;
    wire new_AGEMA_signal_36376 ;
    wire new_AGEMA_signal_36377 ;
    wire new_AGEMA_signal_36378 ;
    wire new_AGEMA_signal_36379 ;
    wire new_AGEMA_signal_36380 ;
    wire new_AGEMA_signal_36381 ;
    wire new_AGEMA_signal_36382 ;
    wire new_AGEMA_signal_36383 ;
    wire new_AGEMA_signal_36384 ;
    wire new_AGEMA_signal_36385 ;
    wire new_AGEMA_signal_36386 ;
    wire new_AGEMA_signal_36387 ;
    wire new_AGEMA_signal_36388 ;
    wire new_AGEMA_signal_36389 ;
    wire new_AGEMA_signal_36390 ;
    wire new_AGEMA_signal_36391 ;
    wire new_AGEMA_signal_36392 ;
    wire new_AGEMA_signal_36393 ;
    wire new_AGEMA_signal_36394 ;
    wire new_AGEMA_signal_36395 ;
    wire new_AGEMA_signal_36396 ;
    wire new_AGEMA_signal_36397 ;
    wire new_AGEMA_signal_36398 ;
    wire new_AGEMA_signal_36399 ;
    wire new_AGEMA_signal_36400 ;
    wire new_AGEMA_signal_36401 ;
    wire new_AGEMA_signal_36402 ;
    wire new_AGEMA_signal_36403 ;
    wire new_AGEMA_signal_36404 ;
    wire new_AGEMA_signal_36405 ;
    wire new_AGEMA_signal_36406 ;
    wire new_AGEMA_signal_36407 ;
    wire new_AGEMA_signal_36408 ;
    wire new_AGEMA_signal_36409 ;
    wire new_AGEMA_signal_36410 ;
    wire new_AGEMA_signal_36411 ;
    wire new_AGEMA_signal_36412 ;
    wire new_AGEMA_signal_36413 ;
    wire new_AGEMA_signal_36414 ;
    wire new_AGEMA_signal_36415 ;
    wire new_AGEMA_signal_36416 ;
    wire new_AGEMA_signal_36417 ;
    wire new_AGEMA_signal_36418 ;
    wire new_AGEMA_signal_36419 ;
    wire new_AGEMA_signal_36420 ;
    wire new_AGEMA_signal_36421 ;
    wire new_AGEMA_signal_36422 ;
    wire new_AGEMA_signal_36423 ;
    wire new_AGEMA_signal_36424 ;
    wire new_AGEMA_signal_36425 ;
    wire new_AGEMA_signal_36426 ;
    wire new_AGEMA_signal_36427 ;
    wire new_AGEMA_signal_36428 ;
    wire new_AGEMA_signal_36429 ;
    wire new_AGEMA_signal_36430 ;
    wire new_AGEMA_signal_36431 ;
    wire new_AGEMA_signal_36432 ;
    wire new_AGEMA_signal_36433 ;
    wire new_AGEMA_signal_36434 ;
    wire new_AGEMA_signal_36435 ;
    wire new_AGEMA_signal_36436 ;
    wire new_AGEMA_signal_36437 ;
    wire new_AGEMA_signal_36438 ;
    wire new_AGEMA_signal_36439 ;
    wire new_AGEMA_signal_36440 ;
    wire new_AGEMA_signal_36441 ;
    wire new_AGEMA_signal_36442 ;
    wire new_AGEMA_signal_36443 ;
    wire new_AGEMA_signal_36444 ;
    wire new_AGEMA_signal_36445 ;
    wire new_AGEMA_signal_36446 ;
    wire new_AGEMA_signal_36447 ;
    wire new_AGEMA_signal_36448 ;
    wire new_AGEMA_signal_36449 ;
    wire new_AGEMA_signal_36450 ;
    wire new_AGEMA_signal_36451 ;
    wire new_AGEMA_signal_36452 ;
    wire new_AGEMA_signal_36453 ;
    wire new_AGEMA_signal_36454 ;
    wire new_AGEMA_signal_36455 ;
    wire new_AGEMA_signal_36456 ;
    wire new_AGEMA_signal_36457 ;
    wire new_AGEMA_signal_36458 ;
    wire new_AGEMA_signal_36459 ;
    wire new_AGEMA_signal_36460 ;
    wire new_AGEMA_signal_36461 ;
    wire new_AGEMA_signal_36462 ;
    wire new_AGEMA_signal_36463 ;
    wire new_AGEMA_signal_36464 ;
    wire new_AGEMA_signal_36465 ;
    wire new_AGEMA_signal_36466 ;
    wire new_AGEMA_signal_36467 ;
    wire new_AGEMA_signal_36468 ;
    wire new_AGEMA_signal_36469 ;
    wire new_AGEMA_signal_36470 ;
    wire new_AGEMA_signal_36471 ;
    wire new_AGEMA_signal_36472 ;
    wire new_AGEMA_signal_36473 ;
    wire new_AGEMA_signal_36474 ;
    wire new_AGEMA_signal_36475 ;
    wire new_AGEMA_signal_36476 ;
    wire new_AGEMA_signal_36477 ;
    wire new_AGEMA_signal_36478 ;
    wire new_AGEMA_signal_36479 ;
    wire new_AGEMA_signal_36480 ;
    wire new_AGEMA_signal_36481 ;
    wire new_AGEMA_signal_36482 ;
    wire new_AGEMA_signal_36483 ;
    wire new_AGEMA_signal_36484 ;
    wire new_AGEMA_signal_36485 ;
    wire new_AGEMA_signal_36486 ;
    wire new_AGEMA_signal_36487 ;
    wire new_AGEMA_signal_36488 ;
    wire new_AGEMA_signal_36489 ;
    wire new_AGEMA_signal_36490 ;
    wire new_AGEMA_signal_36491 ;
    wire new_AGEMA_signal_36492 ;
    wire new_AGEMA_signal_36493 ;
    wire new_AGEMA_signal_36494 ;
    wire new_AGEMA_signal_36495 ;
    wire new_AGEMA_signal_36496 ;
    wire new_AGEMA_signal_36497 ;
    wire new_AGEMA_signal_36498 ;
    wire new_AGEMA_signal_36499 ;
    wire new_AGEMA_signal_36500 ;
    wire new_AGEMA_signal_36501 ;
    wire new_AGEMA_signal_36502 ;
    wire new_AGEMA_signal_36503 ;
    wire new_AGEMA_signal_36504 ;
    wire new_AGEMA_signal_36505 ;
    wire new_AGEMA_signal_36506 ;
    wire new_AGEMA_signal_36507 ;
    wire new_AGEMA_signal_36508 ;
    wire new_AGEMA_signal_36509 ;
    wire new_AGEMA_signal_36510 ;
    wire new_AGEMA_signal_36511 ;
    wire new_AGEMA_signal_36512 ;
    wire new_AGEMA_signal_36513 ;
    wire new_AGEMA_signal_36514 ;
    wire new_AGEMA_signal_36515 ;
    wire new_AGEMA_signal_36516 ;
    wire new_AGEMA_signal_36517 ;
    wire new_AGEMA_signal_36518 ;
    wire new_AGEMA_signal_36519 ;
    wire new_AGEMA_signal_36520 ;
    wire new_AGEMA_signal_36521 ;
    wire new_AGEMA_signal_36522 ;
    wire new_AGEMA_signal_36523 ;
    wire new_AGEMA_signal_36524 ;
    wire new_AGEMA_signal_36525 ;
    wire new_AGEMA_signal_36526 ;
    wire new_AGEMA_signal_36527 ;
    wire new_AGEMA_signal_36528 ;
    wire new_AGEMA_signal_36529 ;
    wire new_AGEMA_signal_36530 ;
    wire new_AGEMA_signal_36531 ;
    wire new_AGEMA_signal_36532 ;
    wire new_AGEMA_signal_36533 ;
    wire new_AGEMA_signal_36534 ;
    wire new_AGEMA_signal_36535 ;
    wire new_AGEMA_signal_36536 ;
    wire new_AGEMA_signal_36537 ;
    wire new_AGEMA_signal_36538 ;
    wire new_AGEMA_signal_36539 ;
    wire new_AGEMA_signal_36540 ;
    wire new_AGEMA_signal_36541 ;
    wire new_AGEMA_signal_36542 ;
    wire new_AGEMA_signal_36543 ;
    wire new_AGEMA_signal_36544 ;
    wire new_AGEMA_signal_36545 ;
    wire new_AGEMA_signal_36546 ;
    wire new_AGEMA_signal_36547 ;
    wire new_AGEMA_signal_36548 ;
    wire new_AGEMA_signal_36549 ;
    wire new_AGEMA_signal_36550 ;
    wire new_AGEMA_signal_36551 ;
    wire new_AGEMA_signal_36552 ;
    wire new_AGEMA_signal_36553 ;
    wire new_AGEMA_signal_36554 ;
    wire new_AGEMA_signal_36555 ;
    wire new_AGEMA_signal_36556 ;
    wire new_AGEMA_signal_36557 ;
    wire new_AGEMA_signal_36558 ;
    wire new_AGEMA_signal_36559 ;
    wire new_AGEMA_signal_36560 ;
    wire new_AGEMA_signal_36561 ;
    wire new_AGEMA_signal_36562 ;
    wire new_AGEMA_signal_36563 ;
    wire new_AGEMA_signal_36564 ;
    wire new_AGEMA_signal_36565 ;
    wire new_AGEMA_signal_36566 ;
    wire new_AGEMA_signal_36567 ;
    wire new_AGEMA_signal_36568 ;
    wire new_AGEMA_signal_36569 ;
    wire new_AGEMA_signal_36570 ;
    wire new_AGEMA_signal_36571 ;
    wire new_AGEMA_signal_36572 ;
    wire new_AGEMA_signal_36573 ;
    wire new_AGEMA_signal_36574 ;
    wire new_AGEMA_signal_36575 ;
    wire new_AGEMA_signal_36576 ;
    wire new_AGEMA_signal_36577 ;
    wire new_AGEMA_signal_36578 ;
    wire new_AGEMA_signal_36579 ;
    wire new_AGEMA_signal_36580 ;
    wire new_AGEMA_signal_36581 ;
    wire new_AGEMA_signal_36582 ;
    wire new_AGEMA_signal_36583 ;
    wire new_AGEMA_signal_36584 ;
    wire new_AGEMA_signal_36585 ;
    wire new_AGEMA_signal_36586 ;
    wire new_AGEMA_signal_36587 ;
    wire new_AGEMA_signal_36588 ;
    wire new_AGEMA_signal_36589 ;
    wire new_AGEMA_signal_36590 ;
    wire new_AGEMA_signal_36591 ;
    wire new_AGEMA_signal_36592 ;
    wire new_AGEMA_signal_36593 ;
    wire new_AGEMA_signal_36594 ;
    wire new_AGEMA_signal_36595 ;
    wire new_AGEMA_signal_36596 ;
    wire new_AGEMA_signal_36597 ;
    wire new_AGEMA_signal_36598 ;
    wire new_AGEMA_signal_36599 ;
    wire new_AGEMA_signal_36600 ;
    wire new_AGEMA_signal_36601 ;
    wire new_AGEMA_signal_36602 ;
    wire new_AGEMA_signal_36603 ;
    wire new_AGEMA_signal_36604 ;
    wire new_AGEMA_signal_36605 ;
    wire new_AGEMA_signal_36606 ;
    wire new_AGEMA_signal_36607 ;
    wire new_AGEMA_signal_36608 ;
    wire new_AGEMA_signal_36609 ;
    wire new_AGEMA_signal_36610 ;
    wire new_AGEMA_signal_36611 ;
    wire new_AGEMA_signal_36612 ;
    wire new_AGEMA_signal_36613 ;
    wire new_AGEMA_signal_36614 ;
    wire new_AGEMA_signal_36615 ;
    wire new_AGEMA_signal_36616 ;
    wire new_AGEMA_signal_36617 ;
    wire new_AGEMA_signal_36618 ;
    wire new_AGEMA_signal_36619 ;
    wire new_AGEMA_signal_36620 ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U986 ( .a ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U987 ( .a ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, RoundInput[100]}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundKey[100]}), .c ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U988 ( .a ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[101]}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, RoundKey[101]}), .c ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U989 ( .a ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, RoundInput[102]}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundKey[102]}), .c ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U990 ( .a ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[103]}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, RoundKey[103]}), .c ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U991 ( .a ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, RoundInput[104]}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundKey[104]}), .c ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U992 ( .a ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[105]}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, RoundKey[105]}), .c ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U993 ( .a ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, RoundInput[106]}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundKey[106]}), .c ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U994 ( .a ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[107]}), .b ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, RoundKey[107]}), .c ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U995 ( .a ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, RoundInput[108]}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundKey[108]}), .c ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U996 ( .a ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[109]}), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, RoundKey[109]}), .c ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U997 ( .a ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, RoundInput[10]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U998 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[110]}), .b ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, RoundKey[110]}), .c ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U999 ( .a ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, RoundInput[111]}), .b ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundKey[111]}), .c ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1000 ( .a ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[112]}), .b ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, RoundKey[112]}), .c ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1001 ( .a ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, RoundInput[113]}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundKey[113]}), .c ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1002 ( .a ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[114]}), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, RoundKey[114]}), .c ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1003 ( .a ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, RoundInput[115]}), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundKey[115]}), .c ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1004 ( .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[116]}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, RoundKey[116]}), .c ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1005 ( .a ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, RoundInput[117]}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundKey[117]}), .c ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1006 ( .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[118]}), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, RoundKey[118]}), .c ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1007 ( .a ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, RoundInput[119]}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundKey[119]}), .c ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1008 ( .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[11]}), .b ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}), .c ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1009 ( .a ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, RoundInput[120]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundKey[120]}), .c ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1010 ( .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[121]}), .b ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, RoundKey[121]}), .c ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1011 ( .a ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, RoundInput[122]}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundKey[122]}), .c ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1012 ( .a ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[123]}), .b ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, RoundKey[123]}), .c ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1013 ( .a ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, RoundInput[124]}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundKey[124]}), .c ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1014 ( .a ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[125]}), .b ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, RoundKey[125]}), .c ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1015 ( .a ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, RoundInput[126]}), .b ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundKey[126]}), .c ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1016 ( .a ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[127]}), .b ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, RoundKey[127]}), .c ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1017 ( .a ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, RoundInput[12]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .c ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1018 ( .a ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[13]}), .b ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .c ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1019 ( .a ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, RoundInput[14]}), .b ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .c ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1020 ( .a ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[15]}), .b ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .c ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1021 ( .a ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, RoundInput[16]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1022 ( .a ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[17]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1023 ( .a ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, RoundInput[18]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1024 ( .a ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[19]}), .b ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}), .c ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1025 ( .a ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, RoundInput[1]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1026 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[20]}), .b ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .c ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1027 ( .a ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, RoundInput[21]}), .b ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .c ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1028 ( .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[22]}), .b ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .c ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1029 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, RoundInput[23]}), .b ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .c ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1030 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[24]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1031 ( .a ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, RoundInput[25]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1032 ( .a ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[26]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1033 ( .a ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, RoundInput[27]}), .b ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}), .c ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1034 ( .a ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[28]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .c ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1035 ( .a ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, RoundInput[29]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .c ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1036 ( .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[2]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1037 ( .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, RoundInput[30]}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .c ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1038 ( .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[31]}), .b ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .c ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1039 ( .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, RoundInput[32]}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundKey[32]}), .c ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1040 ( .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[33]}), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, RoundKey[33]}), .c ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1041 ( .a ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, RoundInput[34]}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundKey[34]}), .c ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1042 ( .a ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[35]}), .b ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKey[35]}), .c ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1043 ( .a ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundInput[36]}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundKey[36]}), .c ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1044 ( .a ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[37]}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKey[37]}), .c ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1045 ( .a ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundInput[38]}), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundKey[38]}), .c ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1046 ( .a ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[39]}), .b ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKey[39]}), .c ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1047 ( .a ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundInput[3]}), .b ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}), .c ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1048 ( .a ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[40]}), .b ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, RoundKey[40]}), .c ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1049 ( .a ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, RoundInput[41]}), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundKey[41]}), .c ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1050 ( .a ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[42]}), .b ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, RoundKey[42]}), .c ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1051 ( .a ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, RoundInput[43]}), .b ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundKey[43]}), .c ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1052 ( .a ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[44]}), .b ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, RoundKey[44]}), .c ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1053 ( .a ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, RoundInput[45]}), .b ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundKey[45]}), .c ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1054 ( .a ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[46]}), .b ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, RoundKey[46]}), .c ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1055 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, RoundInput[47]}), .b ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundKey[47]}), .c ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1056 ( .a ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[48]}), .b ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, RoundKey[48]}), .c ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1057 ( .a ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, RoundInput[49]}), .b ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundKey[49]}), .c ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1058 ( .a ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[4]}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .c ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1059 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, RoundInput[50]}), .b ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundKey[50]}), .c ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1060 ( .a ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[51]}), .b ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, RoundKey[51]}), .c ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1061 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, RoundInput[52]}), .b ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundKey[52]}), .c ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1062 ( .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[53]}), .b ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, RoundKey[53]}), .c ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1063 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, RoundInput[54]}), .b ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundKey[54]}), .c ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1064 ( .a ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[55]}), .b ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, RoundKey[55]}), .c ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1065 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, RoundInput[56]}), .b ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundKey[56]}), .c ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1066 ( .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[57]}), .b ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, RoundKey[57]}), .c ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1067 ( .a ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, RoundInput[58]}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundKey[58]}), .c ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1068 ( .a ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[59]}), .b ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, RoundKey[59]}), .c ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1069 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, RoundInput[5]}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .c ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1070 ( .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[60]}), .b ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, RoundKey[60]}), .c ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1071 ( .a ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, RoundInput[61]}), .b ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, RoundKey[61]}), .c ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1072 ( .a ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, RoundInput[62]}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, RoundKey[62]}), .c ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1073 ( .a ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundInput[63]}), .b ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, RoundKey[63]}), .c ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1074 ( .a ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, RoundInput[64]}), .b ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKey[64]}), .c ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1075 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundInput[65]}), .b ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, RoundKey[65]}), .c ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1076 ( .a ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, RoundInput[66]}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKey[66]}), .c ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1077 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundInput[67]}), .b ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, RoundKey[67]}), .c ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1078 ( .a ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, RoundInput[68]}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKey[68]}), .c ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1079 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundInput[69]}), .b ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, RoundKey[69]}), .c ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1080 ( .a ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, RoundInput[6]}), .b ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .c ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1081 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, RoundInput[70]}), .b ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, RoundKey[70]}), .c ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1082 ( .a ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, RoundInput[71]}), .b ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, RoundKey[71]}), .c ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1083 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, RoundInput[72]}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, RoundKey[72]}), .c ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1084 ( .a ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, RoundInput[73]}), .b ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, RoundKey[73]}), .c ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1085 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, RoundInput[74]}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, RoundKey[74]}), .c ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1086 ( .a ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, RoundInput[75]}), .b ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, RoundKey[75]}), .c ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1087 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, RoundInput[76]}), .b ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, RoundKey[76]}), .c ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1088 ( .a ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, RoundInput[77]}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, RoundKey[77]}), .c ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1089 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, RoundInput[78]}), .b ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, RoundKey[78]}), .c ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1090 ( .a ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, RoundInput[79]}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, RoundKey[79]}), .c ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1091 ( .a ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, RoundInput[7]}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .c ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1092 ( .a ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, RoundInput[80]}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, RoundKey[80]}), .c ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1093 ( .a ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, RoundInput[81]}), .b ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, RoundKey[81]}), .c ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1094 ( .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, RoundInput[82]}), .b ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, RoundKey[82]}), .c ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1095 ( .a ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, RoundInput[83]}), .b ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, RoundKey[83]}), .c ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1096 ( .a ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, RoundInput[84]}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, RoundKey[84]}), .c ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1097 ( .a ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, RoundInput[85]}), .b ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, RoundKey[85]}), .c ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1098 ( .a ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, RoundInput[86]}), .b ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, RoundKey[86]}), .c ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1099 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, RoundInput[87]}), .b ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, RoundKey[87]}), .c ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1100 ( .a ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, RoundInput[88]}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, RoundKey[88]}), .c ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1101 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, RoundInput[89]}), .b ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, RoundKey[89]}), .c ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1102 ( .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, RoundInput[8]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1103 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, RoundInput[90]}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, RoundKey[90]}), .c ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1104 ( .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, RoundInput[91]}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, RoundKey[91]}), .c ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1105 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, RoundInput[92]}), .b ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, RoundKey[92]}), .c ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1106 ( .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, RoundInput[93]}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, RoundKey[93]}), .c ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1107 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, RoundInput[94]}), .b ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, RoundKey[94]}), .c ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1108 ( .a ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, RoundInput[95]}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKey[95]}), .c ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1109 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundInput[96]}), .b ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, RoundKey[96]}), .c ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1110 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, RoundInput[97]}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKey[97]}), .c ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1111 ( .a ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundInput[98]}), .b ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, RoundKey[98]}), .c ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1112 ( .a ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, RoundInput[99]}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKey[99]}), .c ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U1113 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundInput[9]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, new_AGEMA_signal_7669, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, new_AGEMA_signal_7672, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, new_AGEMA_signal_6955, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, new_AGEMA_signal_6982, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, new_AGEMA_signal_7696, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, new_AGEMA_signal_7726, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, new_AGEMA_signal_7750, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, new_AGEMA_signal_7780, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, new_AGEMA_signal_7138, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, new_AGEMA_signal_7804, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, new_AGEMA_signal_7150, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, new_AGEMA_signal_7834, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, new_AGEMA_signal_7858, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, new_AGEMA_signal_7861, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, new_AGEMA_signal_7888, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, new_AGEMA_signal_7912, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, new_AGEMA_signal_7942, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, new_AGEMA_signal_7372, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, new_AGEMA_signal_7966, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, new_AGEMA_signal_7384, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_7995, new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, new_AGEMA_signal_7996, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, new_AGEMA_signal_7450, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, new_AGEMA_signal_8020, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_8025, new_AGEMA_signal_8024, new_AGEMA_signal_8023, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, new_AGEMA_signal_7462, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_8049, new_AGEMA_signal_8048, new_AGEMA_signal_8047, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, new_AGEMA_signal_8050, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, new_AGEMA_signal_7528, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_6297, new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_6297, new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, new_AGEMA_signal_8074, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_8079, new_AGEMA_signal_8078, new_AGEMA_signal_8077, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, new_AGEMA_signal_7540, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .c ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .b ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .c ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_6309, new_AGEMA_signal_6308, new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, new_AGEMA_signal_7561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, new_AGEMA_signal_7564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .c ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .b ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .c ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, new_AGEMA_signal_6826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, new_AGEMA_signal_7588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, new_AGEMA_signal_7591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, new_AGEMA_signal_6838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .c ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .c ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, new_AGEMA_signal_6865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, new_AGEMA_signal_7615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, new_AGEMA_signal_7618, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, new_AGEMA_signal_6877, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .c ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .c ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, new_AGEMA_signal_6904, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, new_AGEMA_signal_7642, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, new_AGEMA_signal_6916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, new_AGEMA_signal_7675, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_25168, new_AGEMA_signal_25167, new_AGEMA_signal_25166, new_AGEMA_signal_25165}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_25172, new_AGEMA_signal_25171, new_AGEMA_signal_25170, new_AGEMA_signal_25169}), .b ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, new_AGEMA_signal_7675, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_25176, new_AGEMA_signal_25175, new_AGEMA_signal_25174, new_AGEMA_signal_25173}), .c ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, new_AGEMA_signal_8170, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, new_AGEMA_signal_8170, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_25180, new_AGEMA_signal_25179, new_AGEMA_signal_25178, new_AGEMA_signal_25177}), .c ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_25184, new_AGEMA_signal_25183, new_AGEMA_signal_25182, new_AGEMA_signal_25181}), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_25188, new_AGEMA_signal_25187, new_AGEMA_signal_25186, new_AGEMA_signal_25185}), .b ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, new_AGEMA_signal_8176, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, new_AGEMA_signal_8182, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_25192, new_AGEMA_signal_25191, new_AGEMA_signal_25190, new_AGEMA_signal_25189}), .c ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, new_AGEMA_signal_8188, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, new_AGEMA_signal_8176, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, new_AGEMA_signal_8182, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, new_AGEMA_signal_8188, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_25196, new_AGEMA_signal_25195, new_AGEMA_signal_25194, new_AGEMA_signal_25193}), .c ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, new_AGEMA_signal_8956, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_25200, new_AGEMA_signal_25199, new_AGEMA_signal_25198, new_AGEMA_signal_25197}), .b ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_25204, new_AGEMA_signal_25203, new_AGEMA_signal_25202, new_AGEMA_signal_25201}), .b ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_25208, new_AGEMA_signal_25207, new_AGEMA_signal_25206, new_AGEMA_signal_25205}), .c ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, new_AGEMA_signal_8200, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, new_AGEMA_signal_8200, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_25212, new_AGEMA_signal_25211, new_AGEMA_signal_25210, new_AGEMA_signal_25209}), .c ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, new_AGEMA_signal_8971, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_25216, new_AGEMA_signal_25215, new_AGEMA_signal_25214, new_AGEMA_signal_25213}), .b ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_25220, new_AGEMA_signal_25219, new_AGEMA_signal_25218, new_AGEMA_signal_25217}), .b ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, new_AGEMA_signal_8206, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, new_AGEMA_signal_8212, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_25224, new_AGEMA_signal_25223, new_AGEMA_signal_25222, new_AGEMA_signal_25221}), .c ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, new_AGEMA_signal_8218, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, new_AGEMA_signal_8206, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, new_AGEMA_signal_8485, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, new_AGEMA_signal_8212, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, new_AGEMA_signal_8218, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, new_AGEMA_signal_8485, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_25228, new_AGEMA_signal_25227, new_AGEMA_signal_25226, new_AGEMA_signal_25225}), .c ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, new_AGEMA_signal_8986, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_25232, new_AGEMA_signal_25231, new_AGEMA_signal_25230, new_AGEMA_signal_25229}), .b ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_25236, new_AGEMA_signal_25235, new_AGEMA_signal_25234, new_AGEMA_signal_25233}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_25240, new_AGEMA_signal_25239, new_AGEMA_signal_25238, new_AGEMA_signal_25237}), .c ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, new_AGEMA_signal_8230, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, new_AGEMA_signal_8497, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, new_AGEMA_signal_8230, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, new_AGEMA_signal_8497, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_25244, new_AGEMA_signal_25243, new_AGEMA_signal_25242, new_AGEMA_signal_25241}), .c ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, new_AGEMA_signal_9001, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_25248, new_AGEMA_signal_25247, new_AGEMA_signal_25246, new_AGEMA_signal_25245}), .b ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, new_AGEMA_signal_7156, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, new_AGEMA_signal_7156, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, new_AGEMA_signal_7162, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_25252, new_AGEMA_signal_25251, new_AGEMA_signal_25250, new_AGEMA_signal_25249}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, new_AGEMA_signal_8236, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, new_AGEMA_signal_7168, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, new_AGEMA_signal_7168, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, new_AGEMA_signal_8242, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_25256, new_AGEMA_signal_25255, new_AGEMA_signal_25254, new_AGEMA_signal_25253}), .c ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, new_AGEMA_signal_7162, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, new_AGEMA_signal_8248, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, new_AGEMA_signal_8236, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, new_AGEMA_signal_8509, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, new_AGEMA_signal_8242, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, new_AGEMA_signal_8248, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, new_AGEMA_signal_8509, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_25260, new_AGEMA_signal_25259, new_AGEMA_signal_25258, new_AGEMA_signal_25257}), .c ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, new_AGEMA_signal_9016, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, new_AGEMA_signal_7837, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_25264, new_AGEMA_signal_25263, new_AGEMA_signal_25262, new_AGEMA_signal_25261}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, new_AGEMA_signal_7843, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_25268, new_AGEMA_signal_25267, new_AGEMA_signal_25266, new_AGEMA_signal_25265}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, new_AGEMA_signal_7849, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, new_AGEMA_signal_7849, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, new_AGEMA_signal_7855, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, new_AGEMA_signal_7855, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, new_AGEMA_signal_7837, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, new_AGEMA_signal_7843, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_25272, new_AGEMA_signal_25271, new_AGEMA_signal_25270, new_AGEMA_signal_25269}), .c ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, new_AGEMA_signal_8260, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, new_AGEMA_signal_8521, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, new_AGEMA_signal_8260, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, new_AGEMA_signal_8521, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_25276, new_AGEMA_signal_25275, new_AGEMA_signal_25274, new_AGEMA_signal_25273}), .c ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, new_AGEMA_signal_9031, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_25280, new_AGEMA_signal_25279, new_AGEMA_signal_25278, new_AGEMA_signal_25277}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, new_AGEMA_signal_7867, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_25284, new_AGEMA_signal_25283, new_AGEMA_signal_25282, new_AGEMA_signal_25281}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, new_AGEMA_signal_8266, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, new_AGEMA_signal_7867, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, new_AGEMA_signal_8272, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_25288, new_AGEMA_signal_25287, new_AGEMA_signal_25286, new_AGEMA_signal_25285}), .c ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, new_AGEMA_signal_8278, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, new_AGEMA_signal_8266, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, new_AGEMA_signal_8533, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, new_AGEMA_signal_8272, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, new_AGEMA_signal_8278, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, new_AGEMA_signal_8533, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_25292, new_AGEMA_signal_25291, new_AGEMA_signal_25290, new_AGEMA_signal_25289}), .c ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, new_AGEMA_signal_9046, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_25296, new_AGEMA_signal_25295, new_AGEMA_signal_25294, new_AGEMA_signal_25293}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_25300, new_AGEMA_signal_25299, new_AGEMA_signal_25298, new_AGEMA_signal_25297}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_25304, new_AGEMA_signal_25303, new_AGEMA_signal_25302, new_AGEMA_signal_25301}), .c ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, new_AGEMA_signal_8290, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, new_AGEMA_signal_8545, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, new_AGEMA_signal_8290, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, new_AGEMA_signal_8545, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_25308, new_AGEMA_signal_25307, new_AGEMA_signal_25306, new_AGEMA_signal_25305}), .c ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_25312, new_AGEMA_signal_25311, new_AGEMA_signal_25310, new_AGEMA_signal_25309}), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_25316, new_AGEMA_signal_25315, new_AGEMA_signal_25314, new_AGEMA_signal_25313}), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, new_AGEMA_signal_8296, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, new_AGEMA_signal_8302, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_25320, new_AGEMA_signal_25319, new_AGEMA_signal_25318, new_AGEMA_signal_25317}), .c ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, new_AGEMA_signal_8308, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, new_AGEMA_signal_8296, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, new_AGEMA_signal_8557, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, new_AGEMA_signal_8302, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, new_AGEMA_signal_8308, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, new_AGEMA_signal_8557, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_25324, new_AGEMA_signal_25323, new_AGEMA_signal_25322, new_AGEMA_signal_25321}), .c ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, new_AGEMA_signal_9076, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_25328, new_AGEMA_signal_25327, new_AGEMA_signal_25326, new_AGEMA_signal_25325}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_25332, new_AGEMA_signal_25331, new_AGEMA_signal_25330, new_AGEMA_signal_25329}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_25336, new_AGEMA_signal_25335, new_AGEMA_signal_25334, new_AGEMA_signal_25333}), .c ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, new_AGEMA_signal_8320, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, new_AGEMA_signal_8569, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, new_AGEMA_signal_8320, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, new_AGEMA_signal_8569, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_25340, new_AGEMA_signal_25339, new_AGEMA_signal_25338, new_AGEMA_signal_25337}), .c ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_25344, new_AGEMA_signal_25343, new_AGEMA_signal_25342, new_AGEMA_signal_25341}), .b ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_25348, new_AGEMA_signal_25347, new_AGEMA_signal_25346, new_AGEMA_signal_25345}), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, new_AGEMA_signal_8326, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, new_AGEMA_signal_8332, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_25352, new_AGEMA_signal_25351, new_AGEMA_signal_25350, new_AGEMA_signal_25349}), .c ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, new_AGEMA_signal_8338, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, new_AGEMA_signal_8326, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, new_AGEMA_signal_8332, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, new_AGEMA_signal_8338, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_25356, new_AGEMA_signal_25355, new_AGEMA_signal_25354, new_AGEMA_signal_25353}), .c ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, new_AGEMA_signal_9106, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, new_AGEMA_signal_7999, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_25360, new_AGEMA_signal_25359, new_AGEMA_signal_25358, new_AGEMA_signal_25357}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, new_AGEMA_signal_8005, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_25364, new_AGEMA_signal_25363, new_AGEMA_signal_25362, new_AGEMA_signal_25361}), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, new_AGEMA_signal_8011, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, new_AGEMA_signal_8011, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, new_AGEMA_signal_8017, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, new_AGEMA_signal_8017, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, new_AGEMA_signal_7999, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, new_AGEMA_signal_8005, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_25368, new_AGEMA_signal_25367, new_AGEMA_signal_25366, new_AGEMA_signal_25365}), .c ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, new_AGEMA_signal_8350, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, new_AGEMA_signal_8350, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_25372, new_AGEMA_signal_25371, new_AGEMA_signal_25370, new_AGEMA_signal_25369}), .c ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_25376, new_AGEMA_signal_25375, new_AGEMA_signal_25374, new_AGEMA_signal_25373}), .b ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, new_AGEMA_signal_8029, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_25380, new_AGEMA_signal_25379, new_AGEMA_signal_25378, new_AGEMA_signal_25377}), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, new_AGEMA_signal_8035, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, new_AGEMA_signal_8356, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, new_AGEMA_signal_8029, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, new_AGEMA_signal_8362, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_25384, new_AGEMA_signal_25383, new_AGEMA_signal_25382, new_AGEMA_signal_25381}), .c ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, new_AGEMA_signal_8035, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, new_AGEMA_signal_8368, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, new_AGEMA_signal_8356, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, new_AGEMA_signal_8362, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, new_AGEMA_signal_8368, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_25388, new_AGEMA_signal_25387, new_AGEMA_signal_25386, new_AGEMA_signal_25385}), .c ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, new_AGEMA_signal_9136, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, new_AGEMA_signal_8053, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_25392, new_AGEMA_signal_25391, new_AGEMA_signal_25390, new_AGEMA_signal_25389}), .b ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, new_AGEMA_signal_8059, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_25396, new_AGEMA_signal_25395, new_AGEMA_signal_25394, new_AGEMA_signal_25393}), .b ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, new_AGEMA_signal_8065, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, new_AGEMA_signal_8065, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, new_AGEMA_signal_8071, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, new_AGEMA_signal_8071, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, new_AGEMA_signal_8053, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, new_AGEMA_signal_8059, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_25400, new_AGEMA_signal_25399, new_AGEMA_signal_25398, new_AGEMA_signal_25397}), .c ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, new_AGEMA_signal_8380, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, new_AGEMA_signal_8380, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_25404, new_AGEMA_signal_25403, new_AGEMA_signal_25402, new_AGEMA_signal_25401}), .c ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_25408, new_AGEMA_signal_25407, new_AGEMA_signal_25406, new_AGEMA_signal_25405}), .b ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, new_AGEMA_signal_8083, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650], Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_25412, new_AGEMA_signal_25411, new_AGEMA_signal_25410, new_AGEMA_signal_25409}), .b ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, new_AGEMA_signal_8089, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, new_AGEMA_signal_8386, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710], Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, new_AGEMA_signal_8083, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, new_AGEMA_signal_8392, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_25416, new_AGEMA_signal_25415, new_AGEMA_signal_25414, new_AGEMA_signal_25413}), .c ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, new_AGEMA_signal_8089, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, new_AGEMA_signal_8398, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, new_AGEMA_signal_8386, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, new_AGEMA_signal_8392, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, new_AGEMA_signal_8398, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_25420, new_AGEMA_signal_25419, new_AGEMA_signal_25418, new_AGEMA_signal_25417}), .c ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, new_AGEMA_signal_9166, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6308, new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, new_AGEMA_signal_7567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_25424, new_AGEMA_signal_25423, new_AGEMA_signal_25422, new_AGEMA_signal_25421}), .b ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, new_AGEMA_signal_7573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770], Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_25428, new_AGEMA_signal_25427, new_AGEMA_signal_25426, new_AGEMA_signal_25425}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, new_AGEMA_signal_7579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, new_AGEMA_signal_7579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, new_AGEMA_signal_8101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830], Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, new_AGEMA_signal_7585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, new_AGEMA_signal_7585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, new_AGEMA_signal_7567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, new_AGEMA_signal_8107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, new_AGEMA_signal_7573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_25432, new_AGEMA_signal_25431, new_AGEMA_signal_25430, new_AGEMA_signal_25429}), .c ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, new_AGEMA_signal_8113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, new_AGEMA_signal_8101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, new_AGEMA_signal_8401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, new_AGEMA_signal_8107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, new_AGEMA_signal_8113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, new_AGEMA_signal_8401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_25436, new_AGEMA_signal_25435, new_AGEMA_signal_25434, new_AGEMA_signal_25433}), .c ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, new_AGEMA_signal_8881, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, new_AGEMA_signal_8647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_25440, new_AGEMA_signal_25439, new_AGEMA_signal_25438, new_AGEMA_signal_25437}), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, new_AGEMA_signal_7597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890], Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_25444, new_AGEMA_signal_25443, new_AGEMA_signal_25442, new_AGEMA_signal_25441}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, new_AGEMA_signal_7603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, new_AGEMA_signal_7597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_25448, new_AGEMA_signal_25447, new_AGEMA_signal_25446, new_AGEMA_signal_25445}), .c ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, new_AGEMA_signal_7603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, new_AGEMA_signal_8413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, new_AGEMA_signal_8413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_25452, new_AGEMA_signal_25451, new_AGEMA_signal_25450, new_AGEMA_signal_25449}), .c ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, new_AGEMA_signal_8896, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, new_AGEMA_signal_8659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950], Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, new_AGEMA_signal_7621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_25456, new_AGEMA_signal_25455, new_AGEMA_signal_25454, new_AGEMA_signal_25453}), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, new_AGEMA_signal_7627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_25460, new_AGEMA_signal_25459, new_AGEMA_signal_25458, new_AGEMA_signal_25457}), .b ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010], Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, new_AGEMA_signal_7633, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, new_AGEMA_signal_7633, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, new_AGEMA_signal_7621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, new_AGEMA_signal_7627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_25464, new_AGEMA_signal_25463, new_AGEMA_signal_25462, new_AGEMA_signal_25461}), .c ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, new_AGEMA_signal_8140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, new_AGEMA_signal_8425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, new_AGEMA_signal_8140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, new_AGEMA_signal_8425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_25468, new_AGEMA_signal_25467, new_AGEMA_signal_25466, new_AGEMA_signal_25465}), .c ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, new_AGEMA_signal_8911, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, new_AGEMA_signal_8671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070], Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_25472, new_AGEMA_signal_25471, new_AGEMA_signal_25470, new_AGEMA_signal_25469}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_25476, new_AGEMA_signal_25475, new_AGEMA_signal_25474, new_AGEMA_signal_25473}), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, new_AGEMA_signal_8146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130], Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, new_AGEMA_signal_8152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_25480, new_AGEMA_signal_25479, new_AGEMA_signal_25478, new_AGEMA_signal_25477}), .c ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, new_AGEMA_signal_8158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, new_AGEMA_signal_8146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, new_AGEMA_signal_8437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, new_AGEMA_signal_8152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, new_AGEMA_signal_8158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, new_AGEMA_signal_8437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_25484, new_AGEMA_signal_25483, new_AGEMA_signal_25482, new_AGEMA_signal_25481}), .c ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, new_AGEMA_signal_8926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, new_AGEMA_signal_8683, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_25165) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_25166) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_6944), .Q (new_AGEMA_signal_25167) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_6945), .Q (new_AGEMA_signal_25168) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_25169) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_25170) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_6956), .Q (new_AGEMA_signal_25171) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_6957), .Q (new_AGEMA_signal_25172) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_25173) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_7669), .Q (new_AGEMA_signal_25174) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_7670), .Q (new_AGEMA_signal_25175) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_7671), .Q (new_AGEMA_signal_25176) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_25177) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_25178) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_7673), .Q (new_AGEMA_signal_25179) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_7674), .Q (new_AGEMA_signal_25180) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_25181) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_6982), .Q (new_AGEMA_signal_25182) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_6983), .Q (new_AGEMA_signal_25183) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_6984), .Q (new_AGEMA_signal_25184) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_25185) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_6994), .Q (new_AGEMA_signal_25186) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_6995), .Q (new_AGEMA_signal_25187) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_6996), .Q (new_AGEMA_signal_25188) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_25189) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_25190) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_7697), .Q (new_AGEMA_signal_25191) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_7698), .Q (new_AGEMA_signal_25192) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_25193) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_7699), .Q (new_AGEMA_signal_25194) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_25195) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_7701), .Q (new_AGEMA_signal_25196) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_25197) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_7021), .Q (new_AGEMA_signal_25198) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_7022), .Q (new_AGEMA_signal_25199) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_25200) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_25201) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_7033), .Q (new_AGEMA_signal_25202) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_7034), .Q (new_AGEMA_signal_25203) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_25204) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_25205) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_7723), .Q (new_AGEMA_signal_25206) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_25207) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_7725), .Q (new_AGEMA_signal_25208) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_25209) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_7726), .Q (new_AGEMA_signal_25210) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_25211) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_7728), .Q (new_AGEMA_signal_25212) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_25213) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_7060), .Q (new_AGEMA_signal_25214) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_7061), .Q (new_AGEMA_signal_25215) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_7062), .Q (new_AGEMA_signal_25216) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_25217) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_7072), .Q (new_AGEMA_signal_25218) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_7073), .Q (new_AGEMA_signal_25219) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_7074), .Q (new_AGEMA_signal_25220) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_25221) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_7750), .Q (new_AGEMA_signal_25222) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_25223) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_7752), .Q (new_AGEMA_signal_25224) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_25225) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_7753), .Q (new_AGEMA_signal_25226) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_7754), .Q (new_AGEMA_signal_25227) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_7755), .Q (new_AGEMA_signal_25228) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T14), .Q (new_AGEMA_signal_25229) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_7099), .Q (new_AGEMA_signal_25230) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_7100), .Q (new_AGEMA_signal_25231) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_7101), .Q (new_AGEMA_signal_25232) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T26), .Q (new_AGEMA_signal_25233) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_25234) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_7112), .Q (new_AGEMA_signal_25235) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_7113), .Q (new_AGEMA_signal_25236) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T24), .Q (new_AGEMA_signal_25237) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_7777), .Q (new_AGEMA_signal_25238) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_7778), .Q (new_AGEMA_signal_25239) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_7779), .Q (new_AGEMA_signal_25240) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T25), .Q (new_AGEMA_signal_25241) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_25242) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_7781), .Q (new_AGEMA_signal_25243) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_7782), .Q (new_AGEMA_signal_25244) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T14), .Q (new_AGEMA_signal_25245) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_7138), .Q (new_AGEMA_signal_25246) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_7139), .Q (new_AGEMA_signal_25247) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_7140), .Q (new_AGEMA_signal_25248) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T26), .Q (new_AGEMA_signal_25249) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_25250) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_25251) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_7152), .Q (new_AGEMA_signal_25252) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T24), .Q (new_AGEMA_signal_25253) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_25254) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_25255) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_7806), .Q (new_AGEMA_signal_25256) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T25), .Q (new_AGEMA_signal_25257) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_25258) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_25259) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_7809), .Q (new_AGEMA_signal_25260) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T14), .Q (new_AGEMA_signal_25261) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_7177), .Q (new_AGEMA_signal_25262) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_7178), .Q (new_AGEMA_signal_25263) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_7179), .Q (new_AGEMA_signal_25264) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T26), .Q (new_AGEMA_signal_25265) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_7189), .Q (new_AGEMA_signal_25266) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_7190), .Q (new_AGEMA_signal_25267) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_7191), .Q (new_AGEMA_signal_25268) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T24), .Q (new_AGEMA_signal_25269) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_25270) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_25271) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_7833), .Q (new_AGEMA_signal_25272) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T25), .Q (new_AGEMA_signal_25273) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_7834), .Q (new_AGEMA_signal_25274) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_25275) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_25276) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T14), .Q (new_AGEMA_signal_25277) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_7216), .Q (new_AGEMA_signal_25278) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_7217), .Q (new_AGEMA_signal_25279) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_7218), .Q (new_AGEMA_signal_25280) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T26), .Q (new_AGEMA_signal_25281) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_7228), .Q (new_AGEMA_signal_25282) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_7229), .Q (new_AGEMA_signal_25283) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_7230), .Q (new_AGEMA_signal_25284) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T24), .Q (new_AGEMA_signal_25285) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_7858), .Q (new_AGEMA_signal_25286) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_7859), .Q (new_AGEMA_signal_25287) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_7860), .Q (new_AGEMA_signal_25288) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T25), .Q (new_AGEMA_signal_25289) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_7861), .Q (new_AGEMA_signal_25290) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_7862), .Q (new_AGEMA_signal_25291) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_7863), .Q (new_AGEMA_signal_25292) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T14), .Q (new_AGEMA_signal_25293) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_25294) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_25295) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_7257), .Q (new_AGEMA_signal_25296) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T26), .Q (new_AGEMA_signal_25297) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_25298) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_25299) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_7269), .Q (new_AGEMA_signal_25300) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T24), .Q (new_AGEMA_signal_25301) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_7885), .Q (new_AGEMA_signal_25302) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_7886), .Q (new_AGEMA_signal_25303) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_7887), .Q (new_AGEMA_signal_25304) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T25), .Q (new_AGEMA_signal_25305) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_25306) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_7889), .Q (new_AGEMA_signal_25307) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_7890), .Q (new_AGEMA_signal_25308) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T14), .Q (new_AGEMA_signal_25309) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_25310) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_25311) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_25312) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T26), .Q (new_AGEMA_signal_25313) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_25314) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_25315) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_25316) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T24), .Q (new_AGEMA_signal_25317) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_25318) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_7913), .Q (new_AGEMA_signal_25319) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_7914), .Q (new_AGEMA_signal_25320) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T25), .Q (new_AGEMA_signal_25321) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_7915), .Q (new_AGEMA_signal_25322) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_25323) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_7917), .Q (new_AGEMA_signal_25324) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T14), .Q (new_AGEMA_signal_25325) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_7333), .Q (new_AGEMA_signal_25326) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_25327) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_25328) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T26), .Q (new_AGEMA_signal_25329) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_7345), .Q (new_AGEMA_signal_25330) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_25331) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_25332) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T24), .Q (new_AGEMA_signal_25333) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_7939), .Q (new_AGEMA_signal_25334) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_25335) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_7941), .Q (new_AGEMA_signal_25336) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T25), .Q (new_AGEMA_signal_25337) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_7942), .Q (new_AGEMA_signal_25338) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_25339) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_7944), .Q (new_AGEMA_signal_25340) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T14), .Q (new_AGEMA_signal_25341) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_25342) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_7373), .Q (new_AGEMA_signal_25343) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_25344) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T26), .Q (new_AGEMA_signal_25345) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_25346) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_7385), .Q (new_AGEMA_signal_25347) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_25348) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T24), .Q (new_AGEMA_signal_25349) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_7966), .Q (new_AGEMA_signal_25350) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_7967), .Q (new_AGEMA_signal_25351) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_7968), .Q (new_AGEMA_signal_25352) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T25), .Q (new_AGEMA_signal_25353) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_7969), .Q (new_AGEMA_signal_25354) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_7970), .Q (new_AGEMA_signal_25355) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_7971), .Q (new_AGEMA_signal_25356) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T14), .Q (new_AGEMA_signal_25357) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_25358) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_25359) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_7413), .Q (new_AGEMA_signal_25360) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T26), .Q (new_AGEMA_signal_25361) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_25362) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_25363) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_7425), .Q (new_AGEMA_signal_25364) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T24), .Q (new_AGEMA_signal_25365) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_7993), .Q (new_AGEMA_signal_25366) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_7994), .Q (new_AGEMA_signal_25367) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_7995), .Q (new_AGEMA_signal_25368) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T25), .Q (new_AGEMA_signal_25369) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_7996), .Q (new_AGEMA_signal_25370) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_7997), .Q (new_AGEMA_signal_25371) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_7998), .Q (new_AGEMA_signal_25372) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T14), .Q (new_AGEMA_signal_25373) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_7450), .Q (new_AGEMA_signal_25374) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_25375) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_25376) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T26), .Q (new_AGEMA_signal_25377) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_25378) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_25379) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_25380) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T24), .Q (new_AGEMA_signal_25381) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_8020), .Q (new_AGEMA_signal_25382) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_8021), .Q (new_AGEMA_signal_25383) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_8022), .Q (new_AGEMA_signal_25384) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T25), .Q (new_AGEMA_signal_25385) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_8023), .Q (new_AGEMA_signal_25386) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_25387) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_8025), .Q (new_AGEMA_signal_25388) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T14), .Q (new_AGEMA_signal_25389) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_7489), .Q (new_AGEMA_signal_25390) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_7490), .Q (new_AGEMA_signal_25391) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_25392) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T26), .Q (new_AGEMA_signal_25393) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_7501), .Q (new_AGEMA_signal_25394) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_25395) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_25396) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T24), .Q (new_AGEMA_signal_25397) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_8047), .Q (new_AGEMA_signal_25398) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_8048), .Q (new_AGEMA_signal_25399) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_8049), .Q (new_AGEMA_signal_25400) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T25), .Q (new_AGEMA_signal_25401) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_8050), .Q (new_AGEMA_signal_25402) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_8051), .Q (new_AGEMA_signal_25403) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_8052), .Q (new_AGEMA_signal_25404) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T14), .Q (new_AGEMA_signal_25405) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_25406) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_7529), .Q (new_AGEMA_signal_25407) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_7530), .Q (new_AGEMA_signal_25408) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T26), .Q (new_AGEMA_signal_25409) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_25410) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_7541), .Q (new_AGEMA_signal_25411) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_7542), .Q (new_AGEMA_signal_25412) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T24), .Q (new_AGEMA_signal_25413) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_8074), .Q (new_AGEMA_signal_25414) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_8075), .Q (new_AGEMA_signal_25415) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_8076), .Q (new_AGEMA_signal_25416) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T25), .Q (new_AGEMA_signal_25417) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_8077), .Q (new_AGEMA_signal_25418) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_8078), .Q (new_AGEMA_signal_25419) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_8079), .Q (new_AGEMA_signal_25420) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_25421) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_6787), .Q (new_AGEMA_signal_25422) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_6788), .Q (new_AGEMA_signal_25423) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_6789), .Q (new_AGEMA_signal_25424) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_25425) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_25426) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_25427) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_6801), .Q (new_AGEMA_signal_25428) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_25429) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_7561), .Q (new_AGEMA_signal_25430) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_7562), .Q (new_AGEMA_signal_25431) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_7563), .Q (new_AGEMA_signal_25432) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_25433) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_25434) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_7565), .Q (new_AGEMA_signal_25435) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_7566), .Q (new_AGEMA_signal_25436) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_25437) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_6826), .Q (new_AGEMA_signal_25438) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_25439) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_25440) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_25441) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_6838), .Q (new_AGEMA_signal_25442) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_6839), .Q (new_AGEMA_signal_25443) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_25444) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_25445) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_25446) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_7589), .Q (new_AGEMA_signal_25447) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_7590), .Q (new_AGEMA_signal_25448) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_25449) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_25450) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_25451) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_7593), .Q (new_AGEMA_signal_25452) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_25453) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_6865), .Q (new_AGEMA_signal_25454) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_6866), .Q (new_AGEMA_signal_25455) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_25456) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_25457) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_6877), .Q (new_AGEMA_signal_25458) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_6878), .Q (new_AGEMA_signal_25459) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_25460) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_25461) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_25462) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_25463) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_7617), .Q (new_AGEMA_signal_25464) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_25465) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7618), .Q (new_AGEMA_signal_25466) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_7619), .Q (new_AGEMA_signal_25467) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_25468) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_25469) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_6904), .Q (new_AGEMA_signal_25470) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_6905), .Q (new_AGEMA_signal_25471) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_6906), .Q (new_AGEMA_signal_25472) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_25473) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_6916), .Q (new_AGEMA_signal_25474) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_6917), .Q (new_AGEMA_signal_25475) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_6918), .Q (new_AGEMA_signal_25476) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_25477) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7642), .Q (new_AGEMA_signal_25478) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_7643), .Q (new_AGEMA_signal_25479) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_7644), .Q (new_AGEMA_signal_25480) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_25481) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_25482) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_7646), .Q (new_AGEMA_signal_25483) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_7647), .Q (new_AGEMA_signal_25484) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C (clk), .D (n321), .Q (new_AGEMA_signal_26125) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C (clk), .D (n315), .Q (new_AGEMA_signal_26129) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C (clk), .D (n316), .Q (new_AGEMA_signal_26133) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C (clk), .D (n317), .Q (new_AGEMA_signal_26137) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C (clk), .D (n318), .Q (new_AGEMA_signal_26141) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C (clk), .D (n319), .Q (new_AGEMA_signal_26145) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C (clk), .D (n320), .Q (new_AGEMA_signal_26149) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_26153) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_26157) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_26161) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C (clk), .D (plaintext_s2[0]), .Q (new_AGEMA_signal_26165) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C (clk), .D (plaintext_s3[0]), .Q (new_AGEMA_signal_26169) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_26173) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_26177) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C (clk), .D (plaintext_s2[1]), .Q (new_AGEMA_signal_26181) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C (clk), .D (plaintext_s3[1]), .Q (new_AGEMA_signal_26185) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_26189) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_26193) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C (clk), .D (plaintext_s2[2]), .Q (new_AGEMA_signal_26197) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C (clk), .D (plaintext_s3[2]), .Q (new_AGEMA_signal_26201) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_26205) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_26209) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C (clk), .D (plaintext_s2[3]), .Q (new_AGEMA_signal_26213) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C (clk), .D (plaintext_s3[3]), .Q (new_AGEMA_signal_26217) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_26221) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_26225) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C (clk), .D (plaintext_s2[4]), .Q (new_AGEMA_signal_26229) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C (clk), .D (plaintext_s3[4]), .Q (new_AGEMA_signal_26233) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_26237) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_26241) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C (clk), .D (plaintext_s2[5]), .Q (new_AGEMA_signal_26245) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C (clk), .D (plaintext_s3[5]), .Q (new_AGEMA_signal_26249) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_26253) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_26257) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C (clk), .D (plaintext_s2[6]), .Q (new_AGEMA_signal_26261) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C (clk), .D (plaintext_s3[6]), .Q (new_AGEMA_signal_26265) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_26269) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_26273) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C (clk), .D (plaintext_s2[7]), .Q (new_AGEMA_signal_26277) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C (clk), .D (plaintext_s3[7]), .Q (new_AGEMA_signal_26281) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_26285) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_26289) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C (clk), .D (plaintext_s2[8]), .Q (new_AGEMA_signal_26293) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C (clk), .D (plaintext_s3[8]), .Q (new_AGEMA_signal_26297) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_26301) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_26305) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C (clk), .D (plaintext_s2[9]), .Q (new_AGEMA_signal_26309) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C (clk), .D (plaintext_s3[9]), .Q (new_AGEMA_signal_26313) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_26317) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_26321) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C (clk), .D (plaintext_s2[10]), .Q (new_AGEMA_signal_26325) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C (clk), .D (plaintext_s3[10]), .Q (new_AGEMA_signal_26329) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_26333) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_26337) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C (clk), .D (plaintext_s2[11]), .Q (new_AGEMA_signal_26341) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C (clk), .D (plaintext_s3[11]), .Q (new_AGEMA_signal_26345) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_26349) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_26353) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C (clk), .D (plaintext_s2[12]), .Q (new_AGEMA_signal_26357) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C (clk), .D (plaintext_s3[12]), .Q (new_AGEMA_signal_26361) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_26365) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_26369) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C (clk), .D (plaintext_s2[13]), .Q (new_AGEMA_signal_26373) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C (clk), .D (plaintext_s3[13]), .Q (new_AGEMA_signal_26377) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_26381) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_26385) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C (clk), .D (plaintext_s2[14]), .Q (new_AGEMA_signal_26389) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C (clk), .D (plaintext_s3[14]), .Q (new_AGEMA_signal_26393) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_26397) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_26401) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C (clk), .D (plaintext_s2[15]), .Q (new_AGEMA_signal_26405) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C (clk), .D (plaintext_s3[15]), .Q (new_AGEMA_signal_26409) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_26413) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_26417) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C (clk), .D (plaintext_s2[16]), .Q (new_AGEMA_signal_26421) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C (clk), .D (plaintext_s3[16]), .Q (new_AGEMA_signal_26425) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_26429) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_26433) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C (clk), .D (plaintext_s2[17]), .Q (new_AGEMA_signal_26437) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C (clk), .D (plaintext_s3[17]), .Q (new_AGEMA_signal_26441) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_26445) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_26449) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C (clk), .D (plaintext_s2[18]), .Q (new_AGEMA_signal_26453) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C (clk), .D (plaintext_s3[18]), .Q (new_AGEMA_signal_26457) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_26461) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_26465) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C (clk), .D (plaintext_s2[19]), .Q (new_AGEMA_signal_26469) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C (clk), .D (plaintext_s3[19]), .Q (new_AGEMA_signal_26473) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_26477) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_26481) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C (clk), .D (plaintext_s2[20]), .Q (new_AGEMA_signal_26485) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C (clk), .D (plaintext_s3[20]), .Q (new_AGEMA_signal_26489) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_26493) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_26497) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C (clk), .D (plaintext_s2[21]), .Q (new_AGEMA_signal_26501) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C (clk), .D (plaintext_s3[21]), .Q (new_AGEMA_signal_26505) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_26509) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_26513) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C (clk), .D (plaintext_s2[22]), .Q (new_AGEMA_signal_26517) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C (clk), .D (plaintext_s3[22]), .Q (new_AGEMA_signal_26521) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_26525) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_26529) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C (clk), .D (plaintext_s2[23]), .Q (new_AGEMA_signal_26533) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C (clk), .D (plaintext_s3[23]), .Q (new_AGEMA_signal_26537) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_26541) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_26545) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C (clk), .D (plaintext_s2[24]), .Q (new_AGEMA_signal_26549) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C (clk), .D (plaintext_s3[24]), .Q (new_AGEMA_signal_26553) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_26557) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_26561) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C (clk), .D (plaintext_s2[25]), .Q (new_AGEMA_signal_26565) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C (clk), .D (plaintext_s3[25]), .Q (new_AGEMA_signal_26569) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_26573) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_26577) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C (clk), .D (plaintext_s2[26]), .Q (new_AGEMA_signal_26581) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C (clk), .D (plaintext_s3[26]), .Q (new_AGEMA_signal_26585) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_26589) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_26593) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C (clk), .D (plaintext_s2[27]), .Q (new_AGEMA_signal_26597) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C (clk), .D (plaintext_s3[27]), .Q (new_AGEMA_signal_26601) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_26605) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_26609) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C (clk), .D (plaintext_s2[28]), .Q (new_AGEMA_signal_26613) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C (clk), .D (plaintext_s3[28]), .Q (new_AGEMA_signal_26617) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_26621) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_26625) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C (clk), .D (plaintext_s2[29]), .Q (new_AGEMA_signal_26629) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C (clk), .D (plaintext_s3[29]), .Q (new_AGEMA_signal_26633) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_26637) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_26641) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C (clk), .D (plaintext_s2[30]), .Q (new_AGEMA_signal_26645) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C (clk), .D (plaintext_s3[30]), .Q (new_AGEMA_signal_26649) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_26653) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_26657) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C (clk), .D (plaintext_s2[31]), .Q (new_AGEMA_signal_26661) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C (clk), .D (plaintext_s3[31]), .Q (new_AGEMA_signal_26665) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_26669) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_26673) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C (clk), .D (plaintext_s2[32]), .Q (new_AGEMA_signal_26677) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C (clk), .D (plaintext_s3[32]), .Q (new_AGEMA_signal_26681) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_26685) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_26689) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C (clk), .D (plaintext_s2[33]), .Q (new_AGEMA_signal_26693) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C (clk), .D (plaintext_s3[33]), .Q (new_AGEMA_signal_26697) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_26701) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_26705) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C (clk), .D (plaintext_s2[34]), .Q (new_AGEMA_signal_26709) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C (clk), .D (plaintext_s3[34]), .Q (new_AGEMA_signal_26713) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_26717) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_26721) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C (clk), .D (plaintext_s2[35]), .Q (new_AGEMA_signal_26725) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C (clk), .D (plaintext_s3[35]), .Q (new_AGEMA_signal_26729) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_26733) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_26737) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C (clk), .D (plaintext_s2[36]), .Q (new_AGEMA_signal_26741) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C (clk), .D (plaintext_s3[36]), .Q (new_AGEMA_signal_26745) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_26749) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_26753) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C (clk), .D (plaintext_s2[37]), .Q (new_AGEMA_signal_26757) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C (clk), .D (plaintext_s3[37]), .Q (new_AGEMA_signal_26761) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_26765) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_26769) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C (clk), .D (plaintext_s2[38]), .Q (new_AGEMA_signal_26773) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C (clk), .D (plaintext_s3[38]), .Q (new_AGEMA_signal_26777) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_26781) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_26785) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C (clk), .D (plaintext_s2[39]), .Q (new_AGEMA_signal_26789) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C (clk), .D (plaintext_s3[39]), .Q (new_AGEMA_signal_26793) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_26797) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_26801) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C (clk), .D (plaintext_s2[40]), .Q (new_AGEMA_signal_26805) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C (clk), .D (plaintext_s3[40]), .Q (new_AGEMA_signal_26809) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_26813) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_26817) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C (clk), .D (plaintext_s2[41]), .Q (new_AGEMA_signal_26821) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C (clk), .D (plaintext_s3[41]), .Q (new_AGEMA_signal_26825) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_26829) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_26833) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C (clk), .D (plaintext_s2[42]), .Q (new_AGEMA_signal_26837) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C (clk), .D (plaintext_s3[42]), .Q (new_AGEMA_signal_26841) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_26845) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_26849) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C (clk), .D (plaintext_s2[43]), .Q (new_AGEMA_signal_26853) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C (clk), .D (plaintext_s3[43]), .Q (new_AGEMA_signal_26857) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_26861) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_26865) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C (clk), .D (plaintext_s2[44]), .Q (new_AGEMA_signal_26869) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C (clk), .D (plaintext_s3[44]), .Q (new_AGEMA_signal_26873) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_26877) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_26881) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C (clk), .D (plaintext_s2[45]), .Q (new_AGEMA_signal_26885) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C (clk), .D (plaintext_s3[45]), .Q (new_AGEMA_signal_26889) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_26893) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_26897) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C (clk), .D (plaintext_s2[46]), .Q (new_AGEMA_signal_26901) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C (clk), .D (plaintext_s3[46]), .Q (new_AGEMA_signal_26905) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_26909) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_26913) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C (clk), .D (plaintext_s2[47]), .Q (new_AGEMA_signal_26917) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C (clk), .D (plaintext_s3[47]), .Q (new_AGEMA_signal_26921) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_26925) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_26929) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C (clk), .D (plaintext_s2[48]), .Q (new_AGEMA_signal_26933) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C (clk), .D (plaintext_s3[48]), .Q (new_AGEMA_signal_26937) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_26941) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_26945) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C (clk), .D (plaintext_s2[49]), .Q (new_AGEMA_signal_26949) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C (clk), .D (plaintext_s3[49]), .Q (new_AGEMA_signal_26953) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_26957) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_26961) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C (clk), .D (plaintext_s2[50]), .Q (new_AGEMA_signal_26965) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C (clk), .D (plaintext_s3[50]), .Q (new_AGEMA_signal_26969) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_26973) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_26977) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C (clk), .D (plaintext_s2[51]), .Q (new_AGEMA_signal_26981) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C (clk), .D (plaintext_s3[51]), .Q (new_AGEMA_signal_26985) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_26989) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_26993) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C (clk), .D (plaintext_s2[52]), .Q (new_AGEMA_signal_26997) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C (clk), .D (plaintext_s3[52]), .Q (new_AGEMA_signal_27001) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_27005) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_27009) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C (clk), .D (plaintext_s2[53]), .Q (new_AGEMA_signal_27013) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C (clk), .D (plaintext_s3[53]), .Q (new_AGEMA_signal_27017) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_27021) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_27025) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C (clk), .D (plaintext_s2[54]), .Q (new_AGEMA_signal_27029) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C (clk), .D (plaintext_s3[54]), .Q (new_AGEMA_signal_27033) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_27037) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_27041) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C (clk), .D (plaintext_s2[55]), .Q (new_AGEMA_signal_27045) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C (clk), .D (plaintext_s3[55]), .Q (new_AGEMA_signal_27049) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_27053) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_27057) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C (clk), .D (plaintext_s2[56]), .Q (new_AGEMA_signal_27061) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C (clk), .D (plaintext_s3[56]), .Q (new_AGEMA_signal_27065) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_27069) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_27073) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C (clk), .D (plaintext_s2[57]), .Q (new_AGEMA_signal_27077) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C (clk), .D (plaintext_s3[57]), .Q (new_AGEMA_signal_27081) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_27085) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_27089) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C (clk), .D (plaintext_s2[58]), .Q (new_AGEMA_signal_27093) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C (clk), .D (plaintext_s3[58]), .Q (new_AGEMA_signal_27097) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_27101) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_27105) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C (clk), .D (plaintext_s2[59]), .Q (new_AGEMA_signal_27109) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C (clk), .D (plaintext_s3[59]), .Q (new_AGEMA_signal_27113) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_27117) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_27121) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C (clk), .D (plaintext_s2[60]), .Q (new_AGEMA_signal_27125) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C (clk), .D (plaintext_s3[60]), .Q (new_AGEMA_signal_27129) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_27133) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_27137) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C (clk), .D (plaintext_s2[61]), .Q (new_AGEMA_signal_27141) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C (clk), .D (plaintext_s3[61]), .Q (new_AGEMA_signal_27145) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_27149) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_27153) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C (clk), .D (plaintext_s2[62]), .Q (new_AGEMA_signal_27157) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C (clk), .D (plaintext_s3[62]), .Q (new_AGEMA_signal_27161) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_27165) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_27169) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C (clk), .D (plaintext_s2[63]), .Q (new_AGEMA_signal_27173) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C (clk), .D (plaintext_s3[63]), .Q (new_AGEMA_signal_27177) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C (clk), .D (plaintext_s0[64]), .Q (new_AGEMA_signal_27181) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C (clk), .D (plaintext_s1[64]), .Q (new_AGEMA_signal_27185) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C (clk), .D (plaintext_s2[64]), .Q (new_AGEMA_signal_27189) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C (clk), .D (plaintext_s3[64]), .Q (new_AGEMA_signal_27193) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C (clk), .D (plaintext_s0[65]), .Q (new_AGEMA_signal_27197) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C (clk), .D (plaintext_s1[65]), .Q (new_AGEMA_signal_27201) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C (clk), .D (plaintext_s2[65]), .Q (new_AGEMA_signal_27205) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C (clk), .D (plaintext_s3[65]), .Q (new_AGEMA_signal_27209) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C (clk), .D (plaintext_s0[66]), .Q (new_AGEMA_signal_27213) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C (clk), .D (plaintext_s1[66]), .Q (new_AGEMA_signal_27217) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C (clk), .D (plaintext_s2[66]), .Q (new_AGEMA_signal_27221) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C (clk), .D (plaintext_s3[66]), .Q (new_AGEMA_signal_27225) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C (clk), .D (plaintext_s0[67]), .Q (new_AGEMA_signal_27229) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C (clk), .D (plaintext_s1[67]), .Q (new_AGEMA_signal_27233) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C (clk), .D (plaintext_s2[67]), .Q (new_AGEMA_signal_27237) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C (clk), .D (plaintext_s3[67]), .Q (new_AGEMA_signal_27241) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C (clk), .D (plaintext_s0[68]), .Q (new_AGEMA_signal_27245) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C (clk), .D (plaintext_s1[68]), .Q (new_AGEMA_signal_27249) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C (clk), .D (plaintext_s2[68]), .Q (new_AGEMA_signal_27253) ) ;
    buf_clk new_AGEMA_reg_buffer_6301 ( .C (clk), .D (plaintext_s3[68]), .Q (new_AGEMA_signal_27257) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C (clk), .D (plaintext_s0[69]), .Q (new_AGEMA_signal_27261) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C (clk), .D (plaintext_s1[69]), .Q (new_AGEMA_signal_27265) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C (clk), .D (plaintext_s2[69]), .Q (new_AGEMA_signal_27269) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C (clk), .D (plaintext_s3[69]), .Q (new_AGEMA_signal_27273) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C (clk), .D (plaintext_s0[70]), .Q (new_AGEMA_signal_27277) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C (clk), .D (plaintext_s1[70]), .Q (new_AGEMA_signal_27281) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C (clk), .D (plaintext_s2[70]), .Q (new_AGEMA_signal_27285) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C (clk), .D (plaintext_s3[70]), .Q (new_AGEMA_signal_27289) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C (clk), .D (plaintext_s0[71]), .Q (new_AGEMA_signal_27293) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C (clk), .D (plaintext_s1[71]), .Q (new_AGEMA_signal_27297) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C (clk), .D (plaintext_s2[71]), .Q (new_AGEMA_signal_27301) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C (clk), .D (plaintext_s3[71]), .Q (new_AGEMA_signal_27305) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C (clk), .D (plaintext_s0[72]), .Q (new_AGEMA_signal_27309) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C (clk), .D (plaintext_s1[72]), .Q (new_AGEMA_signal_27313) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C (clk), .D (plaintext_s2[72]), .Q (new_AGEMA_signal_27317) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C (clk), .D (plaintext_s3[72]), .Q (new_AGEMA_signal_27321) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C (clk), .D (plaintext_s0[73]), .Q (new_AGEMA_signal_27325) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C (clk), .D (plaintext_s1[73]), .Q (new_AGEMA_signal_27329) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C (clk), .D (plaintext_s2[73]), .Q (new_AGEMA_signal_27333) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C (clk), .D (plaintext_s3[73]), .Q (new_AGEMA_signal_27337) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C (clk), .D (plaintext_s0[74]), .Q (new_AGEMA_signal_27341) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C (clk), .D (plaintext_s1[74]), .Q (new_AGEMA_signal_27345) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C (clk), .D (plaintext_s2[74]), .Q (new_AGEMA_signal_27349) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C (clk), .D (plaintext_s3[74]), .Q (new_AGEMA_signal_27353) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C (clk), .D (plaintext_s0[75]), .Q (new_AGEMA_signal_27357) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C (clk), .D (plaintext_s1[75]), .Q (new_AGEMA_signal_27361) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C (clk), .D (plaintext_s2[75]), .Q (new_AGEMA_signal_27365) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C (clk), .D (plaintext_s3[75]), .Q (new_AGEMA_signal_27369) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C (clk), .D (plaintext_s0[76]), .Q (new_AGEMA_signal_27373) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C (clk), .D (plaintext_s1[76]), .Q (new_AGEMA_signal_27377) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C (clk), .D (plaintext_s2[76]), .Q (new_AGEMA_signal_27381) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C (clk), .D (plaintext_s3[76]), .Q (new_AGEMA_signal_27385) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C (clk), .D (plaintext_s0[77]), .Q (new_AGEMA_signal_27389) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C (clk), .D (plaintext_s1[77]), .Q (new_AGEMA_signal_27393) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C (clk), .D (plaintext_s2[77]), .Q (new_AGEMA_signal_27397) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C (clk), .D (plaintext_s3[77]), .Q (new_AGEMA_signal_27401) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C (clk), .D (plaintext_s0[78]), .Q (new_AGEMA_signal_27405) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C (clk), .D (plaintext_s1[78]), .Q (new_AGEMA_signal_27409) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C (clk), .D (plaintext_s2[78]), .Q (new_AGEMA_signal_27413) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C (clk), .D (plaintext_s3[78]), .Q (new_AGEMA_signal_27417) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C (clk), .D (plaintext_s0[79]), .Q (new_AGEMA_signal_27421) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C (clk), .D (plaintext_s1[79]), .Q (new_AGEMA_signal_27425) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C (clk), .D (plaintext_s2[79]), .Q (new_AGEMA_signal_27429) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C (clk), .D (plaintext_s3[79]), .Q (new_AGEMA_signal_27433) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C (clk), .D (plaintext_s0[80]), .Q (new_AGEMA_signal_27437) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C (clk), .D (plaintext_s1[80]), .Q (new_AGEMA_signal_27441) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C (clk), .D (plaintext_s2[80]), .Q (new_AGEMA_signal_27445) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C (clk), .D (plaintext_s3[80]), .Q (new_AGEMA_signal_27449) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C (clk), .D (plaintext_s0[81]), .Q (new_AGEMA_signal_27453) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C (clk), .D (plaintext_s1[81]), .Q (new_AGEMA_signal_27457) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C (clk), .D (plaintext_s2[81]), .Q (new_AGEMA_signal_27461) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C (clk), .D (plaintext_s3[81]), .Q (new_AGEMA_signal_27465) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C (clk), .D (plaintext_s0[82]), .Q (new_AGEMA_signal_27469) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C (clk), .D (plaintext_s1[82]), .Q (new_AGEMA_signal_27473) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C (clk), .D (plaintext_s2[82]), .Q (new_AGEMA_signal_27477) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C (clk), .D (plaintext_s3[82]), .Q (new_AGEMA_signal_27481) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C (clk), .D (plaintext_s0[83]), .Q (new_AGEMA_signal_27485) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C (clk), .D (plaintext_s1[83]), .Q (new_AGEMA_signal_27489) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C (clk), .D (plaintext_s2[83]), .Q (new_AGEMA_signal_27493) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C (clk), .D (plaintext_s3[83]), .Q (new_AGEMA_signal_27497) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C (clk), .D (plaintext_s0[84]), .Q (new_AGEMA_signal_27501) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C (clk), .D (plaintext_s1[84]), .Q (new_AGEMA_signal_27505) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C (clk), .D (plaintext_s2[84]), .Q (new_AGEMA_signal_27509) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C (clk), .D (plaintext_s3[84]), .Q (new_AGEMA_signal_27513) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C (clk), .D (plaintext_s0[85]), .Q (new_AGEMA_signal_27517) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C (clk), .D (plaintext_s1[85]), .Q (new_AGEMA_signal_27521) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C (clk), .D (plaintext_s2[85]), .Q (new_AGEMA_signal_27525) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C (clk), .D (plaintext_s3[85]), .Q (new_AGEMA_signal_27529) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C (clk), .D (plaintext_s0[86]), .Q (new_AGEMA_signal_27533) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C (clk), .D (plaintext_s1[86]), .Q (new_AGEMA_signal_27537) ) ;
    buf_clk new_AGEMA_reg_buffer_6585 ( .C (clk), .D (plaintext_s2[86]), .Q (new_AGEMA_signal_27541) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C (clk), .D (plaintext_s3[86]), .Q (new_AGEMA_signal_27545) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C (clk), .D (plaintext_s0[87]), .Q (new_AGEMA_signal_27549) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C (clk), .D (plaintext_s1[87]), .Q (new_AGEMA_signal_27553) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C (clk), .D (plaintext_s2[87]), .Q (new_AGEMA_signal_27557) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C (clk), .D (plaintext_s3[87]), .Q (new_AGEMA_signal_27561) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C (clk), .D (plaintext_s0[88]), .Q (new_AGEMA_signal_27565) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C (clk), .D (plaintext_s1[88]), .Q (new_AGEMA_signal_27569) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C (clk), .D (plaintext_s2[88]), .Q (new_AGEMA_signal_27573) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C (clk), .D (plaintext_s3[88]), .Q (new_AGEMA_signal_27577) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C (clk), .D (plaintext_s0[89]), .Q (new_AGEMA_signal_27581) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C (clk), .D (plaintext_s1[89]), .Q (new_AGEMA_signal_27585) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C (clk), .D (plaintext_s2[89]), .Q (new_AGEMA_signal_27589) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C (clk), .D (plaintext_s3[89]), .Q (new_AGEMA_signal_27593) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C (clk), .D (plaintext_s0[90]), .Q (new_AGEMA_signal_27597) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C (clk), .D (plaintext_s1[90]), .Q (new_AGEMA_signal_27601) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C (clk), .D (plaintext_s2[90]), .Q (new_AGEMA_signal_27605) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C (clk), .D (plaintext_s3[90]), .Q (new_AGEMA_signal_27609) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C (clk), .D (plaintext_s0[91]), .Q (new_AGEMA_signal_27613) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C (clk), .D (plaintext_s1[91]), .Q (new_AGEMA_signal_27617) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C (clk), .D (plaintext_s2[91]), .Q (new_AGEMA_signal_27621) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C (clk), .D (plaintext_s3[91]), .Q (new_AGEMA_signal_27625) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C (clk), .D (plaintext_s0[92]), .Q (new_AGEMA_signal_27629) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C (clk), .D (plaintext_s1[92]), .Q (new_AGEMA_signal_27633) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C (clk), .D (plaintext_s2[92]), .Q (new_AGEMA_signal_27637) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C (clk), .D (plaintext_s3[92]), .Q (new_AGEMA_signal_27641) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C (clk), .D (plaintext_s0[93]), .Q (new_AGEMA_signal_27645) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C (clk), .D (plaintext_s1[93]), .Q (new_AGEMA_signal_27649) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C (clk), .D (plaintext_s2[93]), .Q (new_AGEMA_signal_27653) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C (clk), .D (plaintext_s3[93]), .Q (new_AGEMA_signal_27657) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C (clk), .D (plaintext_s0[94]), .Q (new_AGEMA_signal_27661) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C (clk), .D (plaintext_s1[94]), .Q (new_AGEMA_signal_27665) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C (clk), .D (plaintext_s2[94]), .Q (new_AGEMA_signal_27669) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C (clk), .D (plaintext_s3[94]), .Q (new_AGEMA_signal_27673) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C (clk), .D (plaintext_s0[95]), .Q (new_AGEMA_signal_27677) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C (clk), .D (plaintext_s1[95]), .Q (new_AGEMA_signal_27681) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C (clk), .D (plaintext_s2[95]), .Q (new_AGEMA_signal_27685) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C (clk), .D (plaintext_s3[95]), .Q (new_AGEMA_signal_27689) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C (clk), .D (plaintext_s0[96]), .Q (new_AGEMA_signal_27693) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C (clk), .D (plaintext_s1[96]), .Q (new_AGEMA_signal_27697) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C (clk), .D (plaintext_s2[96]), .Q (new_AGEMA_signal_27701) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C (clk), .D (plaintext_s3[96]), .Q (new_AGEMA_signal_27705) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C (clk), .D (plaintext_s0[97]), .Q (new_AGEMA_signal_27709) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C (clk), .D (plaintext_s1[97]), .Q (new_AGEMA_signal_27713) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C (clk), .D (plaintext_s2[97]), .Q (new_AGEMA_signal_27717) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C (clk), .D (plaintext_s3[97]), .Q (new_AGEMA_signal_27721) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C (clk), .D (plaintext_s0[98]), .Q (new_AGEMA_signal_27725) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C (clk), .D (plaintext_s1[98]), .Q (new_AGEMA_signal_27729) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C (clk), .D (plaintext_s2[98]), .Q (new_AGEMA_signal_27733) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C (clk), .D (plaintext_s3[98]), .Q (new_AGEMA_signal_27737) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C (clk), .D (plaintext_s0[99]), .Q (new_AGEMA_signal_27741) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C (clk), .D (plaintext_s1[99]), .Q (new_AGEMA_signal_27745) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C (clk), .D (plaintext_s2[99]), .Q (new_AGEMA_signal_27749) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C (clk), .D (plaintext_s3[99]), .Q (new_AGEMA_signal_27753) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C (clk), .D (plaintext_s0[100]), .Q (new_AGEMA_signal_27757) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C (clk), .D (plaintext_s1[100]), .Q (new_AGEMA_signal_27761) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C (clk), .D (plaintext_s2[100]), .Q (new_AGEMA_signal_27765) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C (clk), .D (plaintext_s3[100]), .Q (new_AGEMA_signal_27769) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C (clk), .D (plaintext_s0[101]), .Q (new_AGEMA_signal_27773) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C (clk), .D (plaintext_s1[101]), .Q (new_AGEMA_signal_27777) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C (clk), .D (plaintext_s2[101]), .Q (new_AGEMA_signal_27781) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C (clk), .D (plaintext_s3[101]), .Q (new_AGEMA_signal_27785) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C (clk), .D (plaintext_s0[102]), .Q (new_AGEMA_signal_27789) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C (clk), .D (plaintext_s1[102]), .Q (new_AGEMA_signal_27793) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C (clk), .D (plaintext_s2[102]), .Q (new_AGEMA_signal_27797) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C (clk), .D (plaintext_s3[102]), .Q (new_AGEMA_signal_27801) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C (clk), .D (plaintext_s0[103]), .Q (new_AGEMA_signal_27805) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C (clk), .D (plaintext_s1[103]), .Q (new_AGEMA_signal_27809) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C (clk), .D (plaintext_s2[103]), .Q (new_AGEMA_signal_27813) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C (clk), .D (plaintext_s3[103]), .Q (new_AGEMA_signal_27817) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C (clk), .D (plaintext_s0[104]), .Q (new_AGEMA_signal_27821) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C (clk), .D (plaintext_s1[104]), .Q (new_AGEMA_signal_27825) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C (clk), .D (plaintext_s2[104]), .Q (new_AGEMA_signal_27829) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C (clk), .D (plaintext_s3[104]), .Q (new_AGEMA_signal_27833) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C (clk), .D (plaintext_s0[105]), .Q (new_AGEMA_signal_27837) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C (clk), .D (plaintext_s1[105]), .Q (new_AGEMA_signal_27841) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C (clk), .D (plaintext_s2[105]), .Q (new_AGEMA_signal_27845) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C (clk), .D (plaintext_s3[105]), .Q (new_AGEMA_signal_27849) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C (clk), .D (plaintext_s0[106]), .Q (new_AGEMA_signal_27853) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C (clk), .D (plaintext_s1[106]), .Q (new_AGEMA_signal_27857) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C (clk), .D (plaintext_s2[106]), .Q (new_AGEMA_signal_27861) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C (clk), .D (plaintext_s3[106]), .Q (new_AGEMA_signal_27865) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C (clk), .D (plaintext_s0[107]), .Q (new_AGEMA_signal_27869) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C (clk), .D (plaintext_s1[107]), .Q (new_AGEMA_signal_27873) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C (clk), .D (plaintext_s2[107]), .Q (new_AGEMA_signal_27877) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C (clk), .D (plaintext_s3[107]), .Q (new_AGEMA_signal_27881) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C (clk), .D (plaintext_s0[108]), .Q (new_AGEMA_signal_27885) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C (clk), .D (plaintext_s1[108]), .Q (new_AGEMA_signal_27889) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C (clk), .D (plaintext_s2[108]), .Q (new_AGEMA_signal_27893) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C (clk), .D (plaintext_s3[108]), .Q (new_AGEMA_signal_27897) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C (clk), .D (plaintext_s0[109]), .Q (new_AGEMA_signal_27901) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C (clk), .D (plaintext_s1[109]), .Q (new_AGEMA_signal_27905) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C (clk), .D (plaintext_s2[109]), .Q (new_AGEMA_signal_27909) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C (clk), .D (plaintext_s3[109]), .Q (new_AGEMA_signal_27913) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C (clk), .D (plaintext_s0[110]), .Q (new_AGEMA_signal_27917) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C (clk), .D (plaintext_s1[110]), .Q (new_AGEMA_signal_27921) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C (clk), .D (plaintext_s2[110]), .Q (new_AGEMA_signal_27925) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C (clk), .D (plaintext_s3[110]), .Q (new_AGEMA_signal_27929) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C (clk), .D (plaintext_s0[111]), .Q (new_AGEMA_signal_27933) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C (clk), .D (plaintext_s1[111]), .Q (new_AGEMA_signal_27937) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C (clk), .D (plaintext_s2[111]), .Q (new_AGEMA_signal_27941) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C (clk), .D (plaintext_s3[111]), .Q (new_AGEMA_signal_27945) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C (clk), .D (plaintext_s0[112]), .Q (new_AGEMA_signal_27949) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C (clk), .D (plaintext_s1[112]), .Q (new_AGEMA_signal_27953) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C (clk), .D (plaintext_s2[112]), .Q (new_AGEMA_signal_27957) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C (clk), .D (plaintext_s3[112]), .Q (new_AGEMA_signal_27961) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C (clk), .D (plaintext_s0[113]), .Q (new_AGEMA_signal_27965) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C (clk), .D (plaintext_s1[113]), .Q (new_AGEMA_signal_27969) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C (clk), .D (plaintext_s2[113]), .Q (new_AGEMA_signal_27973) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C (clk), .D (plaintext_s3[113]), .Q (new_AGEMA_signal_27977) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C (clk), .D (plaintext_s0[114]), .Q (new_AGEMA_signal_27981) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C (clk), .D (plaintext_s1[114]), .Q (new_AGEMA_signal_27985) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C (clk), .D (plaintext_s2[114]), .Q (new_AGEMA_signal_27989) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C (clk), .D (plaintext_s3[114]), .Q (new_AGEMA_signal_27993) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C (clk), .D (plaintext_s0[115]), .Q (new_AGEMA_signal_27997) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C (clk), .D (plaintext_s1[115]), .Q (new_AGEMA_signal_28001) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C (clk), .D (plaintext_s2[115]), .Q (new_AGEMA_signal_28005) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C (clk), .D (plaintext_s3[115]), .Q (new_AGEMA_signal_28009) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C (clk), .D (plaintext_s0[116]), .Q (new_AGEMA_signal_28013) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C (clk), .D (plaintext_s1[116]), .Q (new_AGEMA_signal_28017) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C (clk), .D (plaintext_s2[116]), .Q (new_AGEMA_signal_28021) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C (clk), .D (plaintext_s3[116]), .Q (new_AGEMA_signal_28025) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C (clk), .D (plaintext_s0[117]), .Q (new_AGEMA_signal_28029) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C (clk), .D (plaintext_s1[117]), .Q (new_AGEMA_signal_28033) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C (clk), .D (plaintext_s2[117]), .Q (new_AGEMA_signal_28037) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C (clk), .D (plaintext_s3[117]), .Q (new_AGEMA_signal_28041) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C (clk), .D (plaintext_s0[118]), .Q (new_AGEMA_signal_28045) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C (clk), .D (plaintext_s1[118]), .Q (new_AGEMA_signal_28049) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C (clk), .D (plaintext_s2[118]), .Q (new_AGEMA_signal_28053) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C (clk), .D (plaintext_s3[118]), .Q (new_AGEMA_signal_28057) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C (clk), .D (plaintext_s0[119]), .Q (new_AGEMA_signal_28061) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C (clk), .D (plaintext_s1[119]), .Q (new_AGEMA_signal_28065) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C (clk), .D (plaintext_s2[119]), .Q (new_AGEMA_signal_28069) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C (clk), .D (plaintext_s3[119]), .Q (new_AGEMA_signal_28073) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C (clk), .D (plaintext_s0[120]), .Q (new_AGEMA_signal_28077) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C (clk), .D (plaintext_s1[120]), .Q (new_AGEMA_signal_28081) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C (clk), .D (plaintext_s2[120]), .Q (new_AGEMA_signal_28085) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C (clk), .D (plaintext_s3[120]), .Q (new_AGEMA_signal_28089) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C (clk), .D (plaintext_s0[121]), .Q (new_AGEMA_signal_28093) ) ;
    buf_clk new_AGEMA_reg_buffer_7141 ( .C (clk), .D (plaintext_s1[121]), .Q (new_AGEMA_signal_28097) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C (clk), .D (plaintext_s2[121]), .Q (new_AGEMA_signal_28101) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C (clk), .D (plaintext_s3[121]), .Q (new_AGEMA_signal_28105) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C (clk), .D (plaintext_s0[122]), .Q (new_AGEMA_signal_28109) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C (clk), .D (plaintext_s1[122]), .Q (new_AGEMA_signal_28113) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C (clk), .D (plaintext_s2[122]), .Q (new_AGEMA_signal_28117) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C (clk), .D (plaintext_s3[122]), .Q (new_AGEMA_signal_28121) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C (clk), .D (plaintext_s0[123]), .Q (new_AGEMA_signal_28125) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C (clk), .D (plaintext_s1[123]), .Q (new_AGEMA_signal_28129) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C (clk), .D (plaintext_s2[123]), .Q (new_AGEMA_signal_28133) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C (clk), .D (plaintext_s3[123]), .Q (new_AGEMA_signal_28137) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C (clk), .D (plaintext_s0[124]), .Q (new_AGEMA_signal_28141) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C (clk), .D (plaintext_s1[124]), .Q (new_AGEMA_signal_28145) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C (clk), .D (plaintext_s2[124]), .Q (new_AGEMA_signal_28149) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C (clk), .D (plaintext_s3[124]), .Q (new_AGEMA_signal_28153) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C (clk), .D (plaintext_s0[125]), .Q (new_AGEMA_signal_28157) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C (clk), .D (plaintext_s1[125]), .Q (new_AGEMA_signal_28161) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C (clk), .D (plaintext_s2[125]), .Q (new_AGEMA_signal_28165) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C (clk), .D (plaintext_s3[125]), .Q (new_AGEMA_signal_28169) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C (clk), .D (plaintext_s0[126]), .Q (new_AGEMA_signal_28173) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C (clk), .D (plaintext_s1[126]), .Q (new_AGEMA_signal_28177) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C (clk), .D (plaintext_s2[126]), .Q (new_AGEMA_signal_28181) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C (clk), .D (plaintext_s3[126]), .Q (new_AGEMA_signal_28185) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C (clk), .D (plaintext_s0[127]), .Q (new_AGEMA_signal_28189) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C (clk), .D (plaintext_s1[127]), .Q (new_AGEMA_signal_28193) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C (clk), .D (plaintext_s2[127]), .Q (new_AGEMA_signal_28197) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C (clk), .D (plaintext_s3[127]), .Q (new_AGEMA_signal_28201) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_28205) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C (clk), .D (new_AGEMA_signal_6397), .Q (new_AGEMA_signal_28208) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_28211) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_28214) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_28217) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C (clk), .D (new_AGEMA_signal_6937), .Q (new_AGEMA_signal_28220) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C (clk), .D (new_AGEMA_signal_6938), .Q (new_AGEMA_signal_28223) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_28226) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_28229) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_28232) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C (clk), .D (ciphertext_s2[0]), .Q (new_AGEMA_signal_28235) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C (clk), .D (ciphertext_s3[0]), .Q (new_AGEMA_signal_28238) ) ;
    buf_clk new_AGEMA_reg_buffer_7285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_28241) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C (clk), .D (new_AGEMA_signal_6409), .Q (new_AGEMA_signal_28244) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_28247) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_28250) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_28253) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_28256) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C (clk), .D (new_AGEMA_signal_6401), .Q (new_AGEMA_signal_28259) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_28262) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_28265) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C (clk), .D (new_AGEMA_signal_6946), .Q (new_AGEMA_signal_28268) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C (clk), .D (new_AGEMA_signal_6947), .Q (new_AGEMA_signal_28271) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C (clk), .D (new_AGEMA_signal_6948), .Q (new_AGEMA_signal_28274) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_28277) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_28280) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_28283) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_28286) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_28289) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C (clk), .D (new_AGEMA_signal_6418), .Q (new_AGEMA_signal_28292) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_28295) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_28298) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_28301) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C (clk), .D (new_AGEMA_signal_6940), .Q (new_AGEMA_signal_28304) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C (clk), .D (new_AGEMA_signal_6941), .Q (new_AGEMA_signal_28307) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C (clk), .D (new_AGEMA_signal_6942), .Q (new_AGEMA_signal_28310) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_28313) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_28316) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_28319) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_28322) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_28325) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C (clk), .D (new_AGEMA_signal_6952), .Q (new_AGEMA_signal_28328) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C (clk), .D (new_AGEMA_signal_6953), .Q (new_AGEMA_signal_28331) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C (clk), .D (new_AGEMA_signal_6954), .Q (new_AGEMA_signal_28334) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_28337) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_28340) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C (clk), .D (new_AGEMA_signal_6413), .Q (new_AGEMA_signal_28343) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_28346) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_28349) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_28352) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_28355) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_28358) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_28361) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C (clk), .D (new_AGEMA_signal_6415), .Q (new_AGEMA_signal_28364) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_28367) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C (clk), .D (new_AGEMA_signal_6417), .Q (new_AGEMA_signal_28370) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_28373) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C (clk), .D (new_AGEMA_signal_6949), .Q (new_AGEMA_signal_28376) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C (clk), .D (new_AGEMA_signal_6950), .Q (new_AGEMA_signal_28379) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_28382) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_28385) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C (clk), .D (new_AGEMA_signal_5821), .Q (new_AGEMA_signal_28388) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_28391) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_28394) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_28397) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_28400) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_28403) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_28406) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_28409) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_28412) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_28415) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_28418) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_28421) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C (clk), .D (new_AGEMA_signal_6421), .Q (new_AGEMA_signal_28424) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_28427) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_28430) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_28433) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C (clk), .D (new_AGEMA_signal_6976), .Q (new_AGEMA_signal_28436) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C (clk), .D (new_AGEMA_signal_6977), .Q (new_AGEMA_signal_28439) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C (clk), .D (new_AGEMA_signal_6978), .Q (new_AGEMA_signal_28442) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_28445) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_28448) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C (clk), .D (ciphertext_s2[8]), .Q (new_AGEMA_signal_28451) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C (clk), .D (ciphertext_s3[8]), .Q (new_AGEMA_signal_28454) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_28457) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C (clk), .D (new_AGEMA_signal_6433), .Q (new_AGEMA_signal_28460) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_28463) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_28466) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_28469) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C (clk), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_28472) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C (clk), .D (new_AGEMA_signal_6425), .Q (new_AGEMA_signal_28475) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C (clk), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_28478) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_28481) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C (clk), .D (new_AGEMA_signal_6985), .Q (new_AGEMA_signal_28484) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C (clk), .D (new_AGEMA_signal_6986), .Q (new_AGEMA_signal_28487) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_28490) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_28493) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_28496) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_28499) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_28502) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_28505) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C (clk), .D (new_AGEMA_signal_6442), .Q (new_AGEMA_signal_28508) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_28511) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_28514) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_28517) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_28520) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C (clk), .D (new_AGEMA_signal_6980), .Q (new_AGEMA_signal_28523) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C (clk), .D (new_AGEMA_signal_6981), .Q (new_AGEMA_signal_28526) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_28529) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_28532) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_28535) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_28538) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_28541) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_28544) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C (clk), .D (new_AGEMA_signal_6992), .Q (new_AGEMA_signal_28547) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C (clk), .D (new_AGEMA_signal_6993), .Q (new_AGEMA_signal_28550) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_28553) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_28556) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C (clk), .D (new_AGEMA_signal_6437), .Q (new_AGEMA_signal_28559) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_28562) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_28565) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_28568) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_28571) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_28574) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_28577) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_28580) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_28583) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_28586) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_28589) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C (clk), .D (new_AGEMA_signal_6988), .Q (new_AGEMA_signal_28592) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C (clk), .D (new_AGEMA_signal_6989), .Q (new_AGEMA_signal_28595) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C (clk), .D (new_AGEMA_signal_6990), .Q (new_AGEMA_signal_28598) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_28601) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_28604) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_28607) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_28610) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_28613) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_28616) ) ;
    buf_clk new_AGEMA_reg_buffer_7663 ( .C (clk), .D (new_AGEMA_signal_5861), .Q (new_AGEMA_signal_28619) ) ;
    buf_clk new_AGEMA_reg_buffer_7666 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_28622) ) ;
    buf_clk new_AGEMA_reg_buffer_7669 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_28625) ) ;
    buf_clk new_AGEMA_reg_buffer_7672 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_28628) ) ;
    buf_clk new_AGEMA_reg_buffer_7675 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_28631) ) ;
    buf_clk new_AGEMA_reg_buffer_7678 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_28634) ) ;
    buf_clk new_AGEMA_reg_buffer_7681 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_28637) ) ;
    buf_clk new_AGEMA_reg_buffer_7684 ( .C (clk), .D (new_AGEMA_signal_6445), .Q (new_AGEMA_signal_28640) ) ;
    buf_clk new_AGEMA_reg_buffer_7687 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_28643) ) ;
    buf_clk new_AGEMA_reg_buffer_7690 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_28646) ) ;
    buf_clk new_AGEMA_reg_buffer_7693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_28649) ) ;
    buf_clk new_AGEMA_reg_buffer_7696 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_28652) ) ;
    buf_clk new_AGEMA_reg_buffer_7699 ( .C (clk), .D (new_AGEMA_signal_7016), .Q (new_AGEMA_signal_28655) ) ;
    buf_clk new_AGEMA_reg_buffer_7702 ( .C (clk), .D (new_AGEMA_signal_7017), .Q (new_AGEMA_signal_28658) ) ;
    buf_clk new_AGEMA_reg_buffer_7705 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_28661) ) ;
    buf_clk new_AGEMA_reg_buffer_7708 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_28664) ) ;
    buf_clk new_AGEMA_reg_buffer_7711 ( .C (clk), .D (ciphertext_s2[16]), .Q (new_AGEMA_signal_28667) ) ;
    buf_clk new_AGEMA_reg_buffer_7714 ( .C (clk), .D (ciphertext_s3[16]), .Q (new_AGEMA_signal_28670) ) ;
    buf_clk new_AGEMA_reg_buffer_7717 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_28673) ) ;
    buf_clk new_AGEMA_reg_buffer_7720 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_28676) ) ;
    buf_clk new_AGEMA_reg_buffer_7723 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_28679) ) ;
    buf_clk new_AGEMA_reg_buffer_7726 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_28682) ) ;
    buf_clk new_AGEMA_reg_buffer_7729 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_28685) ) ;
    buf_clk new_AGEMA_reg_buffer_7732 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_28688) ) ;
    buf_clk new_AGEMA_reg_buffer_7735 ( .C (clk), .D (new_AGEMA_signal_6449), .Q (new_AGEMA_signal_28691) ) ;
    buf_clk new_AGEMA_reg_buffer_7738 ( .C (clk), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_28694) ) ;
    buf_clk new_AGEMA_reg_buffer_7741 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_28697) ) ;
    buf_clk new_AGEMA_reg_buffer_7744 ( .C (clk), .D (new_AGEMA_signal_7024), .Q (new_AGEMA_signal_28700) ) ;
    buf_clk new_AGEMA_reg_buffer_7747 ( .C (clk), .D (new_AGEMA_signal_7025), .Q (new_AGEMA_signal_28703) ) ;
    buf_clk new_AGEMA_reg_buffer_7750 ( .C (clk), .D (new_AGEMA_signal_7026), .Q (new_AGEMA_signal_28706) ) ;
    buf_clk new_AGEMA_reg_buffer_7753 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_28709) ) ;
    buf_clk new_AGEMA_reg_buffer_7756 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_28712) ) ;
    buf_clk new_AGEMA_reg_buffer_7759 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_28715) ) ;
    buf_clk new_AGEMA_reg_buffer_7762 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_28718) ) ;
    buf_clk new_AGEMA_reg_buffer_7765 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_28721) ) ;
    buf_clk new_AGEMA_reg_buffer_7768 ( .C (clk), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_28724) ) ;
    buf_clk new_AGEMA_reg_buffer_7771 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_28727) ) ;
    buf_clk new_AGEMA_reg_buffer_7774 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_28730) ) ;
    buf_clk new_AGEMA_reg_buffer_7777 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_28733) ) ;
    buf_clk new_AGEMA_reg_buffer_7780 ( .C (clk), .D (new_AGEMA_signal_7018), .Q (new_AGEMA_signal_28736) ) ;
    buf_clk new_AGEMA_reg_buffer_7783 ( .C (clk), .D (new_AGEMA_signal_7019), .Q (new_AGEMA_signal_28739) ) ;
    buf_clk new_AGEMA_reg_buffer_7786 ( .C (clk), .D (new_AGEMA_signal_7020), .Q (new_AGEMA_signal_28742) ) ;
    buf_clk new_AGEMA_reg_buffer_7789 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_28745) ) ;
    buf_clk new_AGEMA_reg_buffer_7792 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_28748) ) ;
    buf_clk new_AGEMA_reg_buffer_7795 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_28751) ) ;
    buf_clk new_AGEMA_reg_buffer_7798 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_28754) ) ;
    buf_clk new_AGEMA_reg_buffer_7801 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_28757) ) ;
    buf_clk new_AGEMA_reg_buffer_7804 ( .C (clk), .D (new_AGEMA_signal_7030), .Q (new_AGEMA_signal_28760) ) ;
    buf_clk new_AGEMA_reg_buffer_7807 ( .C (clk), .D (new_AGEMA_signal_7031), .Q (new_AGEMA_signal_28763) ) ;
    buf_clk new_AGEMA_reg_buffer_7810 ( .C (clk), .D (new_AGEMA_signal_7032), .Q (new_AGEMA_signal_28766) ) ;
    buf_clk new_AGEMA_reg_buffer_7813 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_28769) ) ;
    buf_clk new_AGEMA_reg_buffer_7816 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_28772) ) ;
    buf_clk new_AGEMA_reg_buffer_7819 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_28775) ) ;
    buf_clk new_AGEMA_reg_buffer_7822 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_28778) ) ;
    buf_clk new_AGEMA_reg_buffer_7825 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_28781) ) ;
    buf_clk new_AGEMA_reg_buffer_7828 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_28784) ) ;
    buf_clk new_AGEMA_reg_buffer_7831 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_28787) ) ;
    buf_clk new_AGEMA_reg_buffer_7834 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_28790) ) ;
    buf_clk new_AGEMA_reg_buffer_7837 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_28793) ) ;
    buf_clk new_AGEMA_reg_buffer_7840 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_28796) ) ;
    buf_clk new_AGEMA_reg_buffer_7843 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_28799) ) ;
    buf_clk new_AGEMA_reg_buffer_7846 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_28802) ) ;
    buf_clk new_AGEMA_reg_buffer_7849 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_28805) ) ;
    buf_clk new_AGEMA_reg_buffer_7852 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_28808) ) ;
    buf_clk new_AGEMA_reg_buffer_7855 ( .C (clk), .D (new_AGEMA_signal_7028), .Q (new_AGEMA_signal_28811) ) ;
    buf_clk new_AGEMA_reg_buffer_7858 ( .C (clk), .D (new_AGEMA_signal_7029), .Q (new_AGEMA_signal_28814) ) ;
    buf_clk new_AGEMA_reg_buffer_7861 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_28817) ) ;
    buf_clk new_AGEMA_reg_buffer_7864 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_28820) ) ;
    buf_clk new_AGEMA_reg_buffer_7867 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_28823) ) ;
    buf_clk new_AGEMA_reg_buffer_7870 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_28826) ) ;
    buf_clk new_AGEMA_reg_buffer_7873 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_28829) ) ;
    buf_clk new_AGEMA_reg_buffer_7876 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_28832) ) ;
    buf_clk new_AGEMA_reg_buffer_7879 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_28835) ) ;
    buf_clk new_AGEMA_reg_buffer_7882 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_28838) ) ;
    buf_clk new_AGEMA_reg_buffer_7885 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_28841) ) ;
    buf_clk new_AGEMA_reg_buffer_7888 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_28844) ) ;
    buf_clk new_AGEMA_reg_buffer_7891 ( .C (clk), .D (new_AGEMA_signal_5885), .Q (new_AGEMA_signal_28847) ) ;
    buf_clk new_AGEMA_reg_buffer_7894 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_28850) ) ;
    buf_clk new_AGEMA_reg_buffer_7897 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_28853) ) ;
    buf_clk new_AGEMA_reg_buffer_7900 ( .C (clk), .D (new_AGEMA_signal_6469), .Q (new_AGEMA_signal_28856) ) ;
    buf_clk new_AGEMA_reg_buffer_7903 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_28859) ) ;
    buf_clk new_AGEMA_reg_buffer_7906 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_28862) ) ;
    buf_clk new_AGEMA_reg_buffer_7909 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_28865) ) ;
    buf_clk new_AGEMA_reg_buffer_7912 ( .C (clk), .D (new_AGEMA_signal_7054), .Q (new_AGEMA_signal_28868) ) ;
    buf_clk new_AGEMA_reg_buffer_7915 ( .C (clk), .D (new_AGEMA_signal_7055), .Q (new_AGEMA_signal_28871) ) ;
    buf_clk new_AGEMA_reg_buffer_7918 ( .C (clk), .D (new_AGEMA_signal_7056), .Q (new_AGEMA_signal_28874) ) ;
    buf_clk new_AGEMA_reg_buffer_7921 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_28877) ) ;
    buf_clk new_AGEMA_reg_buffer_7924 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_28880) ) ;
    buf_clk new_AGEMA_reg_buffer_7927 ( .C (clk), .D (ciphertext_s2[24]), .Q (new_AGEMA_signal_28883) ) ;
    buf_clk new_AGEMA_reg_buffer_7930 ( .C (clk), .D (ciphertext_s3[24]), .Q (new_AGEMA_signal_28886) ) ;
    buf_clk new_AGEMA_reg_buffer_7933 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_28889) ) ;
    buf_clk new_AGEMA_reg_buffer_7936 ( .C (clk), .D (new_AGEMA_signal_6481), .Q (new_AGEMA_signal_28892) ) ;
    buf_clk new_AGEMA_reg_buffer_7939 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_28895) ) ;
    buf_clk new_AGEMA_reg_buffer_7942 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_28898) ) ;
    buf_clk new_AGEMA_reg_buffer_7945 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_28901) ) ;
    buf_clk new_AGEMA_reg_buffer_7948 ( .C (clk), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_28904) ) ;
    buf_clk new_AGEMA_reg_buffer_7951 ( .C (clk), .D (new_AGEMA_signal_6473), .Q (new_AGEMA_signal_28907) ) ;
    buf_clk new_AGEMA_reg_buffer_7954 ( .C (clk), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_28910) ) ;
    buf_clk new_AGEMA_reg_buffer_7957 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_28913) ) ;
    buf_clk new_AGEMA_reg_buffer_7960 ( .C (clk), .D (new_AGEMA_signal_7063), .Q (new_AGEMA_signal_28916) ) ;
    buf_clk new_AGEMA_reg_buffer_7963 ( .C (clk), .D (new_AGEMA_signal_7064), .Q (new_AGEMA_signal_28919) ) ;
    buf_clk new_AGEMA_reg_buffer_7966 ( .C (clk), .D (new_AGEMA_signal_7065), .Q (new_AGEMA_signal_28922) ) ;
    buf_clk new_AGEMA_reg_buffer_7969 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_28925) ) ;
    buf_clk new_AGEMA_reg_buffer_7972 ( .C (clk), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_28928) ) ;
    buf_clk new_AGEMA_reg_buffer_7975 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_28931) ) ;
    buf_clk new_AGEMA_reg_buffer_7978 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_28934) ) ;
    buf_clk new_AGEMA_reg_buffer_7981 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_28937) ) ;
    buf_clk new_AGEMA_reg_buffer_7984 ( .C (clk), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_28940) ) ;
    buf_clk new_AGEMA_reg_buffer_7987 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_28943) ) ;
    buf_clk new_AGEMA_reg_buffer_7990 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_28946) ) ;
    buf_clk new_AGEMA_reg_buffer_7993 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_28949) ) ;
    buf_clk new_AGEMA_reg_buffer_7996 ( .C (clk), .D (new_AGEMA_signal_7057), .Q (new_AGEMA_signal_28952) ) ;
    buf_clk new_AGEMA_reg_buffer_7999 ( .C (clk), .D (new_AGEMA_signal_7058), .Q (new_AGEMA_signal_28955) ) ;
    buf_clk new_AGEMA_reg_buffer_8002 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_28958) ) ;
    buf_clk new_AGEMA_reg_buffer_8005 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_28961) ) ;
    buf_clk new_AGEMA_reg_buffer_8008 ( .C (clk), .D (new_AGEMA_signal_6475), .Q (new_AGEMA_signal_28964) ) ;
    buf_clk new_AGEMA_reg_buffer_8011 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_28967) ) ;
    buf_clk new_AGEMA_reg_buffer_8014 ( .C (clk), .D (new_AGEMA_signal_6477), .Q (new_AGEMA_signal_28970) ) ;
    buf_clk new_AGEMA_reg_buffer_8017 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_28973) ) ;
    buf_clk new_AGEMA_reg_buffer_8020 ( .C (clk), .D (new_AGEMA_signal_7069), .Q (new_AGEMA_signal_28976) ) ;
    buf_clk new_AGEMA_reg_buffer_8023 ( .C (clk), .D (new_AGEMA_signal_7070), .Q (new_AGEMA_signal_28979) ) ;
    buf_clk new_AGEMA_reg_buffer_8026 ( .C (clk), .D (new_AGEMA_signal_7071), .Q (new_AGEMA_signal_28982) ) ;
    buf_clk new_AGEMA_reg_buffer_8029 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_28985) ) ;
    buf_clk new_AGEMA_reg_buffer_8032 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_28988) ) ;
    buf_clk new_AGEMA_reg_buffer_8035 ( .C (clk), .D (new_AGEMA_signal_6485), .Q (new_AGEMA_signal_28991) ) ;
    buf_clk new_AGEMA_reg_buffer_8038 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_28994) ) ;
    buf_clk new_AGEMA_reg_buffer_8041 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_28997) ) ;
    buf_clk new_AGEMA_reg_buffer_8044 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_29000) ) ;
    buf_clk new_AGEMA_reg_buffer_8047 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_29003) ) ;
    buf_clk new_AGEMA_reg_buffer_8050 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_29006) ) ;
    buf_clk new_AGEMA_reg_buffer_8053 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_29009) ) ;
    buf_clk new_AGEMA_reg_buffer_8056 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_29012) ) ;
    buf_clk new_AGEMA_reg_buffer_8059 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_29015) ) ;
    buf_clk new_AGEMA_reg_buffer_8062 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_29018) ) ;
    buf_clk new_AGEMA_reg_buffer_8065 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_29021) ) ;
    buf_clk new_AGEMA_reg_buffer_8068 ( .C (clk), .D (new_AGEMA_signal_7066), .Q (new_AGEMA_signal_29024) ) ;
    buf_clk new_AGEMA_reg_buffer_8071 ( .C (clk), .D (new_AGEMA_signal_7067), .Q (new_AGEMA_signal_29027) ) ;
    buf_clk new_AGEMA_reg_buffer_8074 ( .C (clk), .D (new_AGEMA_signal_7068), .Q (new_AGEMA_signal_29030) ) ;
    buf_clk new_AGEMA_reg_buffer_8077 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_29033) ) ;
    buf_clk new_AGEMA_reg_buffer_8080 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_29036) ) ;
    buf_clk new_AGEMA_reg_buffer_8083 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_29039) ) ;
    buf_clk new_AGEMA_reg_buffer_8086 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_29042) ) ;
    buf_clk new_AGEMA_reg_buffer_8089 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_29045) ) ;
    buf_clk new_AGEMA_reg_buffer_8092 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_29048) ) ;
    buf_clk new_AGEMA_reg_buffer_8095 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_29051) ) ;
    buf_clk new_AGEMA_reg_buffer_8098 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_29054) ) ;
    buf_clk new_AGEMA_reg_buffer_8101 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_29057) ) ;
    buf_clk new_AGEMA_reg_buffer_8104 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_29060) ) ;
    buf_clk new_AGEMA_reg_buffer_8107 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_29063) ) ;
    buf_clk new_AGEMA_reg_buffer_8110 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_29066) ) ;
    buf_clk new_AGEMA_reg_buffer_8113 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T6), .Q (new_AGEMA_signal_29069) ) ;
    buf_clk new_AGEMA_reg_buffer_8116 ( .C (clk), .D (new_AGEMA_signal_6493), .Q (new_AGEMA_signal_29072) ) ;
    buf_clk new_AGEMA_reg_buffer_8119 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_29075) ) ;
    buf_clk new_AGEMA_reg_buffer_8122 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_29078) ) ;
    buf_clk new_AGEMA_reg_buffer_8125 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T8), .Q (new_AGEMA_signal_29081) ) ;
    buf_clk new_AGEMA_reg_buffer_8128 ( .C (clk), .D (new_AGEMA_signal_7093), .Q (new_AGEMA_signal_29084) ) ;
    buf_clk new_AGEMA_reg_buffer_8131 ( .C (clk), .D (new_AGEMA_signal_7094), .Q (new_AGEMA_signal_29087) ) ;
    buf_clk new_AGEMA_reg_buffer_8134 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_29090) ) ;
    buf_clk new_AGEMA_reg_buffer_8137 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_29093) ) ;
    buf_clk new_AGEMA_reg_buffer_8140 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_29096) ) ;
    buf_clk new_AGEMA_reg_buffer_8143 ( .C (clk), .D (ciphertext_s2[32]), .Q (new_AGEMA_signal_29099) ) ;
    buf_clk new_AGEMA_reg_buffer_8146 ( .C (clk), .D (ciphertext_s3[32]), .Q (new_AGEMA_signal_29102) ) ;
    buf_clk new_AGEMA_reg_buffer_8149 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T16), .Q (new_AGEMA_signal_29105) ) ;
    buf_clk new_AGEMA_reg_buffer_8152 ( .C (clk), .D (new_AGEMA_signal_6505), .Q (new_AGEMA_signal_29108) ) ;
    buf_clk new_AGEMA_reg_buffer_8155 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_29111) ) ;
    buf_clk new_AGEMA_reg_buffer_8158 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_29114) ) ;
    buf_clk new_AGEMA_reg_buffer_8161 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T9), .Q (new_AGEMA_signal_29117) ) ;
    buf_clk new_AGEMA_reg_buffer_8164 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_29120) ) ;
    buf_clk new_AGEMA_reg_buffer_8167 ( .C (clk), .D (new_AGEMA_signal_6497), .Q (new_AGEMA_signal_29123) ) ;
    buf_clk new_AGEMA_reg_buffer_8170 ( .C (clk), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_29126) ) ;
    buf_clk new_AGEMA_reg_buffer_8173 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T17), .Q (new_AGEMA_signal_29129) ) ;
    buf_clk new_AGEMA_reg_buffer_8176 ( .C (clk), .D (new_AGEMA_signal_7102), .Q (new_AGEMA_signal_29132) ) ;
    buf_clk new_AGEMA_reg_buffer_8179 ( .C (clk), .D (new_AGEMA_signal_7103), .Q (new_AGEMA_signal_29135) ) ;
    buf_clk new_AGEMA_reg_buffer_8182 ( .C (clk), .D (new_AGEMA_signal_7104), .Q (new_AGEMA_signal_29138) ) ;
    buf_clk new_AGEMA_reg_buffer_8185 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T15), .Q (new_AGEMA_signal_29141) ) ;
    buf_clk new_AGEMA_reg_buffer_8188 ( .C (clk), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_29144) ) ;
    buf_clk new_AGEMA_reg_buffer_8191 ( .C (clk), .D (new_AGEMA_signal_6503), .Q (new_AGEMA_signal_29147) ) ;
    buf_clk new_AGEMA_reg_buffer_8194 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_29150) ) ;
    buf_clk new_AGEMA_reg_buffer_8197 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T27), .Q (new_AGEMA_signal_29153) ) ;
    buf_clk new_AGEMA_reg_buffer_8200 ( .C (clk), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_29156) ) ;
    buf_clk new_AGEMA_reg_buffer_8203 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_29159) ) ;
    buf_clk new_AGEMA_reg_buffer_8206 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_29162) ) ;
    buf_clk new_AGEMA_reg_buffer_8209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T10), .Q (new_AGEMA_signal_29165) ) ;
    buf_clk new_AGEMA_reg_buffer_8212 ( .C (clk), .D (new_AGEMA_signal_7096), .Q (new_AGEMA_signal_29168) ) ;
    buf_clk new_AGEMA_reg_buffer_8215 ( .C (clk), .D (new_AGEMA_signal_7097), .Q (new_AGEMA_signal_29171) ) ;
    buf_clk new_AGEMA_reg_buffer_8218 ( .C (clk), .D (new_AGEMA_signal_7098), .Q (new_AGEMA_signal_29174) ) ;
    buf_clk new_AGEMA_reg_buffer_8221 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T13), .Q (new_AGEMA_signal_29177) ) ;
    buf_clk new_AGEMA_reg_buffer_8224 ( .C (clk), .D (new_AGEMA_signal_6499), .Q (new_AGEMA_signal_29180) ) ;
    buf_clk new_AGEMA_reg_buffer_8227 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_29183) ) ;
    buf_clk new_AGEMA_reg_buffer_8230 ( .C (clk), .D (new_AGEMA_signal_6501), .Q (new_AGEMA_signal_29186) ) ;
    buf_clk new_AGEMA_reg_buffer_8233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T23), .Q (new_AGEMA_signal_29189) ) ;
    buf_clk new_AGEMA_reg_buffer_8236 ( .C (clk), .D (new_AGEMA_signal_7108), .Q (new_AGEMA_signal_29192) ) ;
    buf_clk new_AGEMA_reg_buffer_8239 ( .C (clk), .D (new_AGEMA_signal_7109), .Q (new_AGEMA_signal_29195) ) ;
    buf_clk new_AGEMA_reg_buffer_8242 ( .C (clk), .D (new_AGEMA_signal_7110), .Q (new_AGEMA_signal_29198) ) ;
    buf_clk new_AGEMA_reg_buffer_8245 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T19), .Q (new_AGEMA_signal_29201) ) ;
    buf_clk new_AGEMA_reg_buffer_8248 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_29204) ) ;
    buf_clk new_AGEMA_reg_buffer_8251 ( .C (clk), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_29207) ) ;
    buf_clk new_AGEMA_reg_buffer_8254 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_29210) ) ;
    buf_clk new_AGEMA_reg_buffer_8257 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T3), .Q (new_AGEMA_signal_29213) ) ;
    buf_clk new_AGEMA_reg_buffer_8260 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_29216) ) ;
    buf_clk new_AGEMA_reg_buffer_8263 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_29219) ) ;
    buf_clk new_AGEMA_reg_buffer_8266 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_29222) ) ;
    buf_clk new_AGEMA_reg_buffer_8269 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T22), .Q (new_AGEMA_signal_29225) ) ;
    buf_clk new_AGEMA_reg_buffer_8272 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_29228) ) ;
    buf_clk new_AGEMA_reg_buffer_8275 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_29231) ) ;
    buf_clk new_AGEMA_reg_buffer_8278 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_29234) ) ;
    buf_clk new_AGEMA_reg_buffer_8281 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T20), .Q (new_AGEMA_signal_29237) ) ;
    buf_clk new_AGEMA_reg_buffer_8284 ( .C (clk), .D (new_AGEMA_signal_7105), .Q (new_AGEMA_signal_29240) ) ;
    buf_clk new_AGEMA_reg_buffer_8287 ( .C (clk), .D (new_AGEMA_signal_7106), .Q (new_AGEMA_signal_29243) ) ;
    buf_clk new_AGEMA_reg_buffer_8290 ( .C (clk), .D (new_AGEMA_signal_7107), .Q (new_AGEMA_signal_29246) ) ;
    buf_clk new_AGEMA_reg_buffer_8293 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T1), .Q (new_AGEMA_signal_29249) ) ;
    buf_clk new_AGEMA_reg_buffer_8296 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_29252) ) ;
    buf_clk new_AGEMA_reg_buffer_8299 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_29255) ) ;
    buf_clk new_AGEMA_reg_buffer_8302 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_29258) ) ;
    buf_clk new_AGEMA_reg_buffer_8305 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T4), .Q (new_AGEMA_signal_29261) ) ;
    buf_clk new_AGEMA_reg_buffer_8308 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_29264) ) ;
    buf_clk new_AGEMA_reg_buffer_8311 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_29267) ) ;
    buf_clk new_AGEMA_reg_buffer_8314 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_29270) ) ;
    buf_clk new_AGEMA_reg_buffer_8317 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T2), .Q (new_AGEMA_signal_29273) ) ;
    buf_clk new_AGEMA_reg_buffer_8320 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_29276) ) ;
    buf_clk new_AGEMA_reg_buffer_8323 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_29279) ) ;
    buf_clk new_AGEMA_reg_buffer_8326 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_29282) ) ;
    buf_clk new_AGEMA_reg_buffer_8329 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T6), .Q (new_AGEMA_signal_29285) ) ;
    buf_clk new_AGEMA_reg_buffer_8332 ( .C (clk), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_29288) ) ;
    buf_clk new_AGEMA_reg_buffer_8335 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_29291) ) ;
    buf_clk new_AGEMA_reg_buffer_8338 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_29294) ) ;
    buf_clk new_AGEMA_reg_buffer_8341 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T8), .Q (new_AGEMA_signal_29297) ) ;
    buf_clk new_AGEMA_reg_buffer_8344 ( .C (clk), .D (new_AGEMA_signal_7132), .Q (new_AGEMA_signal_29300) ) ;
    buf_clk new_AGEMA_reg_buffer_8347 ( .C (clk), .D (new_AGEMA_signal_7133), .Q (new_AGEMA_signal_29303) ) ;
    buf_clk new_AGEMA_reg_buffer_8350 ( .C (clk), .D (new_AGEMA_signal_7134), .Q (new_AGEMA_signal_29306) ) ;
    buf_clk new_AGEMA_reg_buffer_8353 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_29309) ) ;
    buf_clk new_AGEMA_reg_buffer_8356 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_29312) ) ;
    buf_clk new_AGEMA_reg_buffer_8359 ( .C (clk), .D (ciphertext_s2[40]), .Q (new_AGEMA_signal_29315) ) ;
    buf_clk new_AGEMA_reg_buffer_8362 ( .C (clk), .D (ciphertext_s3[40]), .Q (new_AGEMA_signal_29318) ) ;
    buf_clk new_AGEMA_reg_buffer_8365 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T16), .Q (new_AGEMA_signal_29321) ) ;
    buf_clk new_AGEMA_reg_buffer_8368 ( .C (clk), .D (new_AGEMA_signal_6529), .Q (new_AGEMA_signal_29324) ) ;
    buf_clk new_AGEMA_reg_buffer_8371 ( .C (clk), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_29327) ) ;
    buf_clk new_AGEMA_reg_buffer_8374 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_29330) ) ;
    buf_clk new_AGEMA_reg_buffer_8377 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T9), .Q (new_AGEMA_signal_29333) ) ;
    buf_clk new_AGEMA_reg_buffer_8380 ( .C (clk), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_29336) ) ;
    buf_clk new_AGEMA_reg_buffer_8383 ( .C (clk), .D (new_AGEMA_signal_6521), .Q (new_AGEMA_signal_29339) ) ;
    buf_clk new_AGEMA_reg_buffer_8386 ( .C (clk), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_29342) ) ;
    buf_clk new_AGEMA_reg_buffer_8389 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T17), .Q (new_AGEMA_signal_29345) ) ;
    buf_clk new_AGEMA_reg_buffer_8392 ( .C (clk), .D (new_AGEMA_signal_7141), .Q (new_AGEMA_signal_29348) ) ;
    buf_clk new_AGEMA_reg_buffer_8395 ( .C (clk), .D (new_AGEMA_signal_7142), .Q (new_AGEMA_signal_29351) ) ;
    buf_clk new_AGEMA_reg_buffer_8398 ( .C (clk), .D (new_AGEMA_signal_7143), .Q (new_AGEMA_signal_29354) ) ;
    buf_clk new_AGEMA_reg_buffer_8401 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T15), .Q (new_AGEMA_signal_29357) ) ;
    buf_clk new_AGEMA_reg_buffer_8404 ( .C (clk), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_29360) ) ;
    buf_clk new_AGEMA_reg_buffer_8407 ( .C (clk), .D (new_AGEMA_signal_6527), .Q (new_AGEMA_signal_29363) ) ;
    buf_clk new_AGEMA_reg_buffer_8410 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_29366) ) ;
    buf_clk new_AGEMA_reg_buffer_8413 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T27), .Q (new_AGEMA_signal_29369) ) ;
    buf_clk new_AGEMA_reg_buffer_8416 ( .C (clk), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_29372) ) ;
    buf_clk new_AGEMA_reg_buffer_8419 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_29375) ) ;
    buf_clk new_AGEMA_reg_buffer_8422 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_29378) ) ;
    buf_clk new_AGEMA_reg_buffer_8425 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T10), .Q (new_AGEMA_signal_29381) ) ;
    buf_clk new_AGEMA_reg_buffer_8428 ( .C (clk), .D (new_AGEMA_signal_7135), .Q (new_AGEMA_signal_29384) ) ;
    buf_clk new_AGEMA_reg_buffer_8431 ( .C (clk), .D (new_AGEMA_signal_7136), .Q (new_AGEMA_signal_29387) ) ;
    buf_clk new_AGEMA_reg_buffer_8434 ( .C (clk), .D (new_AGEMA_signal_7137), .Q (new_AGEMA_signal_29390) ) ;
    buf_clk new_AGEMA_reg_buffer_8437 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T13), .Q (new_AGEMA_signal_29393) ) ;
    buf_clk new_AGEMA_reg_buffer_8440 ( .C (clk), .D (new_AGEMA_signal_6523), .Q (new_AGEMA_signal_29396) ) ;
    buf_clk new_AGEMA_reg_buffer_8443 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_29399) ) ;
    buf_clk new_AGEMA_reg_buffer_8446 ( .C (clk), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_29402) ) ;
    buf_clk new_AGEMA_reg_buffer_8449 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T23), .Q (new_AGEMA_signal_29405) ) ;
    buf_clk new_AGEMA_reg_buffer_8452 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_29408) ) ;
    buf_clk new_AGEMA_reg_buffer_8455 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_29411) ) ;
    buf_clk new_AGEMA_reg_buffer_8458 ( .C (clk), .D (new_AGEMA_signal_7149), .Q (new_AGEMA_signal_29414) ) ;
    buf_clk new_AGEMA_reg_buffer_8461 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T19), .Q (new_AGEMA_signal_29417) ) ;
    buf_clk new_AGEMA_reg_buffer_8464 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_29420) ) ;
    buf_clk new_AGEMA_reg_buffer_8467 ( .C (clk), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_29423) ) ;
    buf_clk new_AGEMA_reg_buffer_8470 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_29426) ) ;
    buf_clk new_AGEMA_reg_buffer_8473 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T3), .Q (new_AGEMA_signal_29429) ) ;
    buf_clk new_AGEMA_reg_buffer_8476 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_29432) ) ;
    buf_clk new_AGEMA_reg_buffer_8479 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_29435) ) ;
    buf_clk new_AGEMA_reg_buffer_8482 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_29438) ) ;
    buf_clk new_AGEMA_reg_buffer_8485 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T22), .Q (new_AGEMA_signal_29441) ) ;
    buf_clk new_AGEMA_reg_buffer_8488 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_29444) ) ;
    buf_clk new_AGEMA_reg_buffer_8491 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_29447) ) ;
    buf_clk new_AGEMA_reg_buffer_8494 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_29450) ) ;
    buf_clk new_AGEMA_reg_buffer_8497 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T20), .Q (new_AGEMA_signal_29453) ) ;
    buf_clk new_AGEMA_reg_buffer_8500 ( .C (clk), .D (new_AGEMA_signal_7144), .Q (new_AGEMA_signal_29456) ) ;
    buf_clk new_AGEMA_reg_buffer_8503 ( .C (clk), .D (new_AGEMA_signal_7145), .Q (new_AGEMA_signal_29459) ) ;
    buf_clk new_AGEMA_reg_buffer_8506 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_29462) ) ;
    buf_clk new_AGEMA_reg_buffer_8509 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T1), .Q (new_AGEMA_signal_29465) ) ;
    buf_clk new_AGEMA_reg_buffer_8512 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_29468) ) ;
    buf_clk new_AGEMA_reg_buffer_8515 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_29471) ) ;
    buf_clk new_AGEMA_reg_buffer_8518 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_29474) ) ;
    buf_clk new_AGEMA_reg_buffer_8521 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T4), .Q (new_AGEMA_signal_29477) ) ;
    buf_clk new_AGEMA_reg_buffer_8524 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_29480) ) ;
    buf_clk new_AGEMA_reg_buffer_8527 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_29483) ) ;
    buf_clk new_AGEMA_reg_buffer_8530 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_29486) ) ;
    buf_clk new_AGEMA_reg_buffer_8533 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T2), .Q (new_AGEMA_signal_29489) ) ;
    buf_clk new_AGEMA_reg_buffer_8536 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_29492) ) ;
    buf_clk new_AGEMA_reg_buffer_8539 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_29495) ) ;
    buf_clk new_AGEMA_reg_buffer_8542 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_29498) ) ;
    buf_clk new_AGEMA_reg_buffer_8545 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T6), .Q (new_AGEMA_signal_29501) ) ;
    buf_clk new_AGEMA_reg_buffer_8548 ( .C (clk), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_29504) ) ;
    buf_clk new_AGEMA_reg_buffer_8551 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_29507) ) ;
    buf_clk new_AGEMA_reg_buffer_8554 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_29510) ) ;
    buf_clk new_AGEMA_reg_buffer_8557 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T8), .Q (new_AGEMA_signal_29513) ) ;
    buf_clk new_AGEMA_reg_buffer_8560 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_29516) ) ;
    buf_clk new_AGEMA_reg_buffer_8563 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_29519) ) ;
    buf_clk new_AGEMA_reg_buffer_8566 ( .C (clk), .D (new_AGEMA_signal_7173), .Q (new_AGEMA_signal_29522) ) ;
    buf_clk new_AGEMA_reg_buffer_8569 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_29525) ) ;
    buf_clk new_AGEMA_reg_buffer_8572 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_29528) ) ;
    buf_clk new_AGEMA_reg_buffer_8575 ( .C (clk), .D (ciphertext_s2[48]), .Q (new_AGEMA_signal_29531) ) ;
    buf_clk new_AGEMA_reg_buffer_8578 ( .C (clk), .D (ciphertext_s3[48]), .Q (new_AGEMA_signal_29534) ) ;
    buf_clk new_AGEMA_reg_buffer_8581 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T16), .Q (new_AGEMA_signal_29537) ) ;
    buf_clk new_AGEMA_reg_buffer_8584 ( .C (clk), .D (new_AGEMA_signal_6553), .Q (new_AGEMA_signal_29540) ) ;
    buf_clk new_AGEMA_reg_buffer_8587 ( .C (clk), .D (new_AGEMA_signal_6554), .Q (new_AGEMA_signal_29543) ) ;
    buf_clk new_AGEMA_reg_buffer_8590 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_29546) ) ;
    buf_clk new_AGEMA_reg_buffer_8593 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T9), .Q (new_AGEMA_signal_29549) ) ;
    buf_clk new_AGEMA_reg_buffer_8596 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_29552) ) ;
    buf_clk new_AGEMA_reg_buffer_8599 ( .C (clk), .D (new_AGEMA_signal_6545), .Q (new_AGEMA_signal_29555) ) ;
    buf_clk new_AGEMA_reg_buffer_8602 ( .C (clk), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_29558) ) ;
    buf_clk new_AGEMA_reg_buffer_8605 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T17), .Q (new_AGEMA_signal_29561) ) ;
    buf_clk new_AGEMA_reg_buffer_8608 ( .C (clk), .D (new_AGEMA_signal_7180), .Q (new_AGEMA_signal_29564) ) ;
    buf_clk new_AGEMA_reg_buffer_8611 ( .C (clk), .D (new_AGEMA_signal_7181), .Q (new_AGEMA_signal_29567) ) ;
    buf_clk new_AGEMA_reg_buffer_8614 ( .C (clk), .D (new_AGEMA_signal_7182), .Q (new_AGEMA_signal_29570) ) ;
    buf_clk new_AGEMA_reg_buffer_8617 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T15), .Q (new_AGEMA_signal_29573) ) ;
    buf_clk new_AGEMA_reg_buffer_8620 ( .C (clk), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_29576) ) ;
    buf_clk new_AGEMA_reg_buffer_8623 ( .C (clk), .D (new_AGEMA_signal_6551), .Q (new_AGEMA_signal_29579) ) ;
    buf_clk new_AGEMA_reg_buffer_8626 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_29582) ) ;
    buf_clk new_AGEMA_reg_buffer_8629 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T27), .Q (new_AGEMA_signal_29585) ) ;
    buf_clk new_AGEMA_reg_buffer_8632 ( .C (clk), .D (new_AGEMA_signal_6562), .Q (new_AGEMA_signal_29588) ) ;
    buf_clk new_AGEMA_reg_buffer_8635 ( .C (clk), .D (new_AGEMA_signal_6563), .Q (new_AGEMA_signal_29591) ) ;
    buf_clk new_AGEMA_reg_buffer_8638 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_29594) ) ;
    buf_clk new_AGEMA_reg_buffer_8641 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T10), .Q (new_AGEMA_signal_29597) ) ;
    buf_clk new_AGEMA_reg_buffer_8644 ( .C (clk), .D (new_AGEMA_signal_7174), .Q (new_AGEMA_signal_29600) ) ;
    buf_clk new_AGEMA_reg_buffer_8647 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_29603) ) ;
    buf_clk new_AGEMA_reg_buffer_8650 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_29606) ) ;
    buf_clk new_AGEMA_reg_buffer_8653 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T13), .Q (new_AGEMA_signal_29609) ) ;
    buf_clk new_AGEMA_reg_buffer_8656 ( .C (clk), .D (new_AGEMA_signal_6547), .Q (new_AGEMA_signal_29612) ) ;
    buf_clk new_AGEMA_reg_buffer_8659 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_29615) ) ;
    buf_clk new_AGEMA_reg_buffer_8662 ( .C (clk), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_29618) ) ;
    buf_clk new_AGEMA_reg_buffer_8665 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T23), .Q (new_AGEMA_signal_29621) ) ;
    buf_clk new_AGEMA_reg_buffer_8668 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_29624) ) ;
    buf_clk new_AGEMA_reg_buffer_8671 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_29627) ) ;
    buf_clk new_AGEMA_reg_buffer_8674 ( .C (clk), .D (new_AGEMA_signal_7188), .Q (new_AGEMA_signal_29630) ) ;
    buf_clk new_AGEMA_reg_buffer_8677 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T19), .Q (new_AGEMA_signal_29633) ) ;
    buf_clk new_AGEMA_reg_buffer_8680 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_29636) ) ;
    buf_clk new_AGEMA_reg_buffer_8683 ( .C (clk), .D (new_AGEMA_signal_6557), .Q (new_AGEMA_signal_29639) ) ;
    buf_clk new_AGEMA_reg_buffer_8686 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_29642) ) ;
    buf_clk new_AGEMA_reg_buffer_8689 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T3), .Q (new_AGEMA_signal_29645) ) ;
    buf_clk new_AGEMA_reg_buffer_8692 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_29648) ) ;
    buf_clk new_AGEMA_reg_buffer_8695 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_29651) ) ;
    buf_clk new_AGEMA_reg_buffer_8698 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_29654) ) ;
    buf_clk new_AGEMA_reg_buffer_8701 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T22), .Q (new_AGEMA_signal_29657) ) ;
    buf_clk new_AGEMA_reg_buffer_8704 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_29660) ) ;
    buf_clk new_AGEMA_reg_buffer_8707 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_29663) ) ;
    buf_clk new_AGEMA_reg_buffer_8710 ( .C (clk), .D (new_AGEMA_signal_6561), .Q (new_AGEMA_signal_29666) ) ;
    buf_clk new_AGEMA_reg_buffer_8713 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T20), .Q (new_AGEMA_signal_29669) ) ;
    buf_clk new_AGEMA_reg_buffer_8716 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_29672) ) ;
    buf_clk new_AGEMA_reg_buffer_8719 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_29675) ) ;
    buf_clk new_AGEMA_reg_buffer_8722 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_29678) ) ;
    buf_clk new_AGEMA_reg_buffer_8725 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T1), .Q (new_AGEMA_signal_29681) ) ;
    buf_clk new_AGEMA_reg_buffer_8728 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_29684) ) ;
    buf_clk new_AGEMA_reg_buffer_8731 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_29687) ) ;
    buf_clk new_AGEMA_reg_buffer_8734 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_29690) ) ;
    buf_clk new_AGEMA_reg_buffer_8737 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T4), .Q (new_AGEMA_signal_29693) ) ;
    buf_clk new_AGEMA_reg_buffer_8740 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_29696) ) ;
    buf_clk new_AGEMA_reg_buffer_8743 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_29699) ) ;
    buf_clk new_AGEMA_reg_buffer_8746 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_29702) ) ;
    buf_clk new_AGEMA_reg_buffer_8749 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T2), .Q (new_AGEMA_signal_29705) ) ;
    buf_clk new_AGEMA_reg_buffer_8752 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_29708) ) ;
    buf_clk new_AGEMA_reg_buffer_8755 ( .C (clk), .D (new_AGEMA_signal_6005), .Q (new_AGEMA_signal_29711) ) ;
    buf_clk new_AGEMA_reg_buffer_8758 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_29714) ) ;
    buf_clk new_AGEMA_reg_buffer_8761 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T6), .Q (new_AGEMA_signal_29717) ) ;
    buf_clk new_AGEMA_reg_buffer_8764 ( .C (clk), .D (new_AGEMA_signal_6565), .Q (new_AGEMA_signal_29720) ) ;
    buf_clk new_AGEMA_reg_buffer_8767 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_29723) ) ;
    buf_clk new_AGEMA_reg_buffer_8770 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_29726) ) ;
    buf_clk new_AGEMA_reg_buffer_8773 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T8), .Q (new_AGEMA_signal_29729) ) ;
    buf_clk new_AGEMA_reg_buffer_8776 ( .C (clk), .D (new_AGEMA_signal_7210), .Q (new_AGEMA_signal_29732) ) ;
    buf_clk new_AGEMA_reg_buffer_8779 ( .C (clk), .D (new_AGEMA_signal_7211), .Q (new_AGEMA_signal_29735) ) ;
    buf_clk new_AGEMA_reg_buffer_8782 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_29738) ) ;
    buf_clk new_AGEMA_reg_buffer_8785 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_29741) ) ;
    buf_clk new_AGEMA_reg_buffer_8788 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_29744) ) ;
    buf_clk new_AGEMA_reg_buffer_8791 ( .C (clk), .D (ciphertext_s2[56]), .Q (new_AGEMA_signal_29747) ) ;
    buf_clk new_AGEMA_reg_buffer_8794 ( .C (clk), .D (ciphertext_s3[56]), .Q (new_AGEMA_signal_29750) ) ;
    buf_clk new_AGEMA_reg_buffer_8797 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T16), .Q (new_AGEMA_signal_29753) ) ;
    buf_clk new_AGEMA_reg_buffer_8800 ( .C (clk), .D (new_AGEMA_signal_6577), .Q (new_AGEMA_signal_29756) ) ;
    buf_clk new_AGEMA_reg_buffer_8803 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_29759) ) ;
    buf_clk new_AGEMA_reg_buffer_8806 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_29762) ) ;
    buf_clk new_AGEMA_reg_buffer_8809 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T9), .Q (new_AGEMA_signal_29765) ) ;
    buf_clk new_AGEMA_reg_buffer_8812 ( .C (clk), .D (new_AGEMA_signal_6568), .Q (new_AGEMA_signal_29768) ) ;
    buf_clk new_AGEMA_reg_buffer_8815 ( .C (clk), .D (new_AGEMA_signal_6569), .Q (new_AGEMA_signal_29771) ) ;
    buf_clk new_AGEMA_reg_buffer_8818 ( .C (clk), .D (new_AGEMA_signal_6570), .Q (new_AGEMA_signal_29774) ) ;
    buf_clk new_AGEMA_reg_buffer_8821 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T17), .Q (new_AGEMA_signal_29777) ) ;
    buf_clk new_AGEMA_reg_buffer_8824 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_29780) ) ;
    buf_clk new_AGEMA_reg_buffer_8827 ( .C (clk), .D (new_AGEMA_signal_7220), .Q (new_AGEMA_signal_29783) ) ;
    buf_clk new_AGEMA_reg_buffer_8830 ( .C (clk), .D (new_AGEMA_signal_7221), .Q (new_AGEMA_signal_29786) ) ;
    buf_clk new_AGEMA_reg_buffer_8833 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T15), .Q (new_AGEMA_signal_29789) ) ;
    buf_clk new_AGEMA_reg_buffer_8836 ( .C (clk), .D (new_AGEMA_signal_6574), .Q (new_AGEMA_signal_29792) ) ;
    buf_clk new_AGEMA_reg_buffer_8839 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_29795) ) ;
    buf_clk new_AGEMA_reg_buffer_8842 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_29798) ) ;
    buf_clk new_AGEMA_reg_buffer_8845 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T27), .Q (new_AGEMA_signal_29801) ) ;
    buf_clk new_AGEMA_reg_buffer_8848 ( .C (clk), .D (new_AGEMA_signal_6586), .Q (new_AGEMA_signal_29804) ) ;
    buf_clk new_AGEMA_reg_buffer_8851 ( .C (clk), .D (new_AGEMA_signal_6587), .Q (new_AGEMA_signal_29807) ) ;
    buf_clk new_AGEMA_reg_buffer_8854 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_29810) ) ;
    buf_clk new_AGEMA_reg_buffer_8857 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T10), .Q (new_AGEMA_signal_29813) ) ;
    buf_clk new_AGEMA_reg_buffer_8860 ( .C (clk), .D (new_AGEMA_signal_7213), .Q (new_AGEMA_signal_29816) ) ;
    buf_clk new_AGEMA_reg_buffer_8863 ( .C (clk), .D (new_AGEMA_signal_7214), .Q (new_AGEMA_signal_29819) ) ;
    buf_clk new_AGEMA_reg_buffer_8866 ( .C (clk), .D (new_AGEMA_signal_7215), .Q (new_AGEMA_signal_29822) ) ;
    buf_clk new_AGEMA_reg_buffer_8869 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T13), .Q (new_AGEMA_signal_29825) ) ;
    buf_clk new_AGEMA_reg_buffer_8872 ( .C (clk), .D (new_AGEMA_signal_6571), .Q (new_AGEMA_signal_29828) ) ;
    buf_clk new_AGEMA_reg_buffer_8875 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_29831) ) ;
    buf_clk new_AGEMA_reg_buffer_8878 ( .C (clk), .D (new_AGEMA_signal_6573), .Q (new_AGEMA_signal_29834) ) ;
    buf_clk new_AGEMA_reg_buffer_8881 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T23), .Q (new_AGEMA_signal_29837) ) ;
    buf_clk new_AGEMA_reg_buffer_8884 ( .C (clk), .D (new_AGEMA_signal_7225), .Q (new_AGEMA_signal_29840) ) ;
    buf_clk new_AGEMA_reg_buffer_8887 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_29843) ) ;
    buf_clk new_AGEMA_reg_buffer_8890 ( .C (clk), .D (new_AGEMA_signal_7227), .Q (new_AGEMA_signal_29846) ) ;
    buf_clk new_AGEMA_reg_buffer_8893 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T19), .Q (new_AGEMA_signal_29849) ) ;
    buf_clk new_AGEMA_reg_buffer_8896 ( .C (clk), .D (new_AGEMA_signal_6580), .Q (new_AGEMA_signal_29852) ) ;
    buf_clk new_AGEMA_reg_buffer_8899 ( .C (clk), .D (new_AGEMA_signal_6581), .Q (new_AGEMA_signal_29855) ) ;
    buf_clk new_AGEMA_reg_buffer_8902 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_29858) ) ;
    buf_clk new_AGEMA_reg_buffer_8905 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T3), .Q (new_AGEMA_signal_29861) ) ;
    buf_clk new_AGEMA_reg_buffer_8908 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_29864) ) ;
    buf_clk new_AGEMA_reg_buffer_8911 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_29867) ) ;
    buf_clk new_AGEMA_reg_buffer_8914 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_29870) ) ;
    buf_clk new_AGEMA_reg_buffer_8917 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T22), .Q (new_AGEMA_signal_29873) ) ;
    buf_clk new_AGEMA_reg_buffer_8920 ( .C (clk), .D (new_AGEMA_signal_6583), .Q (new_AGEMA_signal_29876) ) ;
    buf_clk new_AGEMA_reg_buffer_8923 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_29879) ) ;
    buf_clk new_AGEMA_reg_buffer_8926 ( .C (clk), .D (new_AGEMA_signal_6585), .Q (new_AGEMA_signal_29882) ) ;
    buf_clk new_AGEMA_reg_buffer_8929 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T20), .Q (new_AGEMA_signal_29885) ) ;
    buf_clk new_AGEMA_reg_buffer_8932 ( .C (clk), .D (new_AGEMA_signal_7222), .Q (new_AGEMA_signal_29888) ) ;
    buf_clk new_AGEMA_reg_buffer_8935 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_29891) ) ;
    buf_clk new_AGEMA_reg_buffer_8938 ( .C (clk), .D (new_AGEMA_signal_7224), .Q (new_AGEMA_signal_29894) ) ;
    buf_clk new_AGEMA_reg_buffer_8941 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T1), .Q (new_AGEMA_signal_29897) ) ;
    buf_clk new_AGEMA_reg_buffer_8944 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_29900) ) ;
    buf_clk new_AGEMA_reg_buffer_8947 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_29903) ) ;
    buf_clk new_AGEMA_reg_buffer_8950 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_29906) ) ;
    buf_clk new_AGEMA_reg_buffer_8953 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T4), .Q (new_AGEMA_signal_29909) ) ;
    buf_clk new_AGEMA_reg_buffer_8956 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_29912) ) ;
    buf_clk new_AGEMA_reg_buffer_8959 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_29915) ) ;
    buf_clk new_AGEMA_reg_buffer_8962 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_29918) ) ;
    buf_clk new_AGEMA_reg_buffer_8965 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T2), .Q (new_AGEMA_signal_29921) ) ;
    buf_clk new_AGEMA_reg_buffer_8968 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_29924) ) ;
    buf_clk new_AGEMA_reg_buffer_8971 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_29927) ) ;
    buf_clk new_AGEMA_reg_buffer_8974 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_29930) ) ;
    buf_clk new_AGEMA_reg_buffer_8977 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T6), .Q (new_AGEMA_signal_29933) ) ;
    buf_clk new_AGEMA_reg_buffer_8980 ( .C (clk), .D (new_AGEMA_signal_6589), .Q (new_AGEMA_signal_29936) ) ;
    buf_clk new_AGEMA_reg_buffer_8983 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_29939) ) ;
    buf_clk new_AGEMA_reg_buffer_8986 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_29942) ) ;
    buf_clk new_AGEMA_reg_buffer_8989 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T8), .Q (new_AGEMA_signal_29945) ) ;
    buf_clk new_AGEMA_reg_buffer_8992 ( .C (clk), .D (new_AGEMA_signal_7249), .Q (new_AGEMA_signal_29948) ) ;
    buf_clk new_AGEMA_reg_buffer_8995 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_29951) ) ;
    buf_clk new_AGEMA_reg_buffer_8998 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_29954) ) ;
    buf_clk new_AGEMA_reg_buffer_9001 ( .C (clk), .D (ciphertext_s0[64]), .Q (new_AGEMA_signal_29957) ) ;
    buf_clk new_AGEMA_reg_buffer_9004 ( .C (clk), .D (ciphertext_s1[64]), .Q (new_AGEMA_signal_29960) ) ;
    buf_clk new_AGEMA_reg_buffer_9007 ( .C (clk), .D (ciphertext_s2[64]), .Q (new_AGEMA_signal_29963) ) ;
    buf_clk new_AGEMA_reg_buffer_9010 ( .C (clk), .D (ciphertext_s3[64]), .Q (new_AGEMA_signal_29966) ) ;
    buf_clk new_AGEMA_reg_buffer_9013 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T16), .Q (new_AGEMA_signal_29969) ) ;
    buf_clk new_AGEMA_reg_buffer_9016 ( .C (clk), .D (new_AGEMA_signal_6601), .Q (new_AGEMA_signal_29972) ) ;
    buf_clk new_AGEMA_reg_buffer_9019 ( .C (clk), .D (new_AGEMA_signal_6602), .Q (new_AGEMA_signal_29975) ) ;
    buf_clk new_AGEMA_reg_buffer_9022 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_29978) ) ;
    buf_clk new_AGEMA_reg_buffer_9025 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T9), .Q (new_AGEMA_signal_29981) ) ;
    buf_clk new_AGEMA_reg_buffer_9028 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_29984) ) ;
    buf_clk new_AGEMA_reg_buffer_9031 ( .C (clk), .D (new_AGEMA_signal_6593), .Q (new_AGEMA_signal_29987) ) ;
    buf_clk new_AGEMA_reg_buffer_9034 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_29990) ) ;
    buf_clk new_AGEMA_reg_buffer_9037 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T17), .Q (new_AGEMA_signal_29993) ) ;
    buf_clk new_AGEMA_reg_buffer_9040 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_29996) ) ;
    buf_clk new_AGEMA_reg_buffer_9043 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_29999) ) ;
    buf_clk new_AGEMA_reg_buffer_9046 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_30002) ) ;
    buf_clk new_AGEMA_reg_buffer_9049 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T15), .Q (new_AGEMA_signal_30005) ) ;
    buf_clk new_AGEMA_reg_buffer_9052 ( .C (clk), .D (new_AGEMA_signal_6598), .Q (new_AGEMA_signal_30008) ) ;
    buf_clk new_AGEMA_reg_buffer_9055 ( .C (clk), .D (new_AGEMA_signal_6599), .Q (new_AGEMA_signal_30011) ) ;
    buf_clk new_AGEMA_reg_buffer_9058 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_30014) ) ;
    buf_clk new_AGEMA_reg_buffer_9061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T27), .Q (new_AGEMA_signal_30017) ) ;
    buf_clk new_AGEMA_reg_buffer_9064 ( .C (clk), .D (new_AGEMA_signal_6610), .Q (new_AGEMA_signal_30020) ) ;
    buf_clk new_AGEMA_reg_buffer_9067 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_30023) ) ;
    buf_clk new_AGEMA_reg_buffer_9070 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_30026) ) ;
    buf_clk new_AGEMA_reg_buffer_9073 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T10), .Q (new_AGEMA_signal_30029) ) ;
    buf_clk new_AGEMA_reg_buffer_9076 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_30032) ) ;
    buf_clk new_AGEMA_reg_buffer_9079 ( .C (clk), .D (new_AGEMA_signal_7253), .Q (new_AGEMA_signal_30035) ) ;
    buf_clk new_AGEMA_reg_buffer_9082 ( .C (clk), .D (new_AGEMA_signal_7254), .Q (new_AGEMA_signal_30038) ) ;
    buf_clk new_AGEMA_reg_buffer_9085 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T13), .Q (new_AGEMA_signal_30041) ) ;
    buf_clk new_AGEMA_reg_buffer_9088 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_30044) ) ;
    buf_clk new_AGEMA_reg_buffer_9091 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_30047) ) ;
    buf_clk new_AGEMA_reg_buffer_9094 ( .C (clk), .D (new_AGEMA_signal_6597), .Q (new_AGEMA_signal_30050) ) ;
    buf_clk new_AGEMA_reg_buffer_9097 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T23), .Q (new_AGEMA_signal_30053) ) ;
    buf_clk new_AGEMA_reg_buffer_9100 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_30056) ) ;
    buf_clk new_AGEMA_reg_buffer_9103 ( .C (clk), .D (new_AGEMA_signal_7265), .Q (new_AGEMA_signal_30059) ) ;
    buf_clk new_AGEMA_reg_buffer_9106 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_30062) ) ;
    buf_clk new_AGEMA_reg_buffer_9109 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T19), .Q (new_AGEMA_signal_30065) ) ;
    buf_clk new_AGEMA_reg_buffer_9112 ( .C (clk), .D (new_AGEMA_signal_6604), .Q (new_AGEMA_signal_30068) ) ;
    buf_clk new_AGEMA_reg_buffer_9115 ( .C (clk), .D (new_AGEMA_signal_6605), .Q (new_AGEMA_signal_30071) ) ;
    buf_clk new_AGEMA_reg_buffer_9118 ( .C (clk), .D (new_AGEMA_signal_6606), .Q (new_AGEMA_signal_30074) ) ;
    buf_clk new_AGEMA_reg_buffer_9121 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T3), .Q (new_AGEMA_signal_30077) ) ;
    buf_clk new_AGEMA_reg_buffer_9124 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_30080) ) ;
    buf_clk new_AGEMA_reg_buffer_9127 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_30083) ) ;
    buf_clk new_AGEMA_reg_buffer_9130 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_30086) ) ;
    buf_clk new_AGEMA_reg_buffer_9133 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T22), .Q (new_AGEMA_signal_30089) ) ;
    buf_clk new_AGEMA_reg_buffer_9136 ( .C (clk), .D (new_AGEMA_signal_6607), .Q (new_AGEMA_signal_30092) ) ;
    buf_clk new_AGEMA_reg_buffer_9139 ( .C (clk), .D (new_AGEMA_signal_6608), .Q (new_AGEMA_signal_30095) ) ;
    buf_clk new_AGEMA_reg_buffer_9142 ( .C (clk), .D (new_AGEMA_signal_6609), .Q (new_AGEMA_signal_30098) ) ;
    buf_clk new_AGEMA_reg_buffer_9145 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T20), .Q (new_AGEMA_signal_30101) ) ;
    buf_clk new_AGEMA_reg_buffer_9148 ( .C (clk), .D (new_AGEMA_signal_7261), .Q (new_AGEMA_signal_30104) ) ;
    buf_clk new_AGEMA_reg_buffer_9151 ( .C (clk), .D (new_AGEMA_signal_7262), .Q (new_AGEMA_signal_30107) ) ;
    buf_clk new_AGEMA_reg_buffer_9154 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_30110) ) ;
    buf_clk new_AGEMA_reg_buffer_9157 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T1), .Q (new_AGEMA_signal_30113) ) ;
    buf_clk new_AGEMA_reg_buffer_9160 ( .C (clk), .D (new_AGEMA_signal_6061), .Q (new_AGEMA_signal_30116) ) ;
    buf_clk new_AGEMA_reg_buffer_9163 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_30119) ) ;
    buf_clk new_AGEMA_reg_buffer_9166 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_30122) ) ;
    buf_clk new_AGEMA_reg_buffer_9169 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T4), .Q (new_AGEMA_signal_30125) ) ;
    buf_clk new_AGEMA_reg_buffer_9172 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_30128) ) ;
    buf_clk new_AGEMA_reg_buffer_9175 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_30131) ) ;
    buf_clk new_AGEMA_reg_buffer_9178 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_30134) ) ;
    buf_clk new_AGEMA_reg_buffer_9181 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T2), .Q (new_AGEMA_signal_30137) ) ;
    buf_clk new_AGEMA_reg_buffer_9184 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_30140) ) ;
    buf_clk new_AGEMA_reg_buffer_9187 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_30143) ) ;
    buf_clk new_AGEMA_reg_buffer_9190 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_30146) ) ;
    buf_clk new_AGEMA_reg_buffer_9193 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T6), .Q (new_AGEMA_signal_30149) ) ;
    buf_clk new_AGEMA_reg_buffer_9196 ( .C (clk), .D (new_AGEMA_signal_6613), .Q (new_AGEMA_signal_30152) ) ;
    buf_clk new_AGEMA_reg_buffer_9199 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_30155) ) ;
    buf_clk new_AGEMA_reg_buffer_9202 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_30158) ) ;
    buf_clk new_AGEMA_reg_buffer_9205 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T8), .Q (new_AGEMA_signal_30161) ) ;
    buf_clk new_AGEMA_reg_buffer_9208 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_30164) ) ;
    buf_clk new_AGEMA_reg_buffer_9211 ( .C (clk), .D (new_AGEMA_signal_7289), .Q (new_AGEMA_signal_30167) ) ;
    buf_clk new_AGEMA_reg_buffer_9214 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_30170) ) ;
    buf_clk new_AGEMA_reg_buffer_9217 ( .C (clk), .D (ciphertext_s0[72]), .Q (new_AGEMA_signal_30173) ) ;
    buf_clk new_AGEMA_reg_buffer_9220 ( .C (clk), .D (ciphertext_s1[72]), .Q (new_AGEMA_signal_30176) ) ;
    buf_clk new_AGEMA_reg_buffer_9223 ( .C (clk), .D (ciphertext_s2[72]), .Q (new_AGEMA_signal_30179) ) ;
    buf_clk new_AGEMA_reg_buffer_9226 ( .C (clk), .D (ciphertext_s3[72]), .Q (new_AGEMA_signal_30182) ) ;
    buf_clk new_AGEMA_reg_buffer_9229 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T16), .Q (new_AGEMA_signal_30185) ) ;
    buf_clk new_AGEMA_reg_buffer_9232 ( .C (clk), .D (new_AGEMA_signal_6625), .Q (new_AGEMA_signal_30188) ) ;
    buf_clk new_AGEMA_reg_buffer_9235 ( .C (clk), .D (new_AGEMA_signal_6626), .Q (new_AGEMA_signal_30191) ) ;
    buf_clk new_AGEMA_reg_buffer_9238 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_30194) ) ;
    buf_clk new_AGEMA_reg_buffer_9241 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T9), .Q (new_AGEMA_signal_30197) ) ;
    buf_clk new_AGEMA_reg_buffer_9244 ( .C (clk), .D (new_AGEMA_signal_6616), .Q (new_AGEMA_signal_30200) ) ;
    buf_clk new_AGEMA_reg_buffer_9247 ( .C (clk), .D (new_AGEMA_signal_6617), .Q (new_AGEMA_signal_30203) ) ;
    buf_clk new_AGEMA_reg_buffer_9250 ( .C (clk), .D (new_AGEMA_signal_6618), .Q (new_AGEMA_signal_30206) ) ;
    buf_clk new_AGEMA_reg_buffer_9253 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T17), .Q (new_AGEMA_signal_30209) ) ;
    buf_clk new_AGEMA_reg_buffer_9256 ( .C (clk), .D (new_AGEMA_signal_7297), .Q (new_AGEMA_signal_30212) ) ;
    buf_clk new_AGEMA_reg_buffer_9259 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_30215) ) ;
    buf_clk new_AGEMA_reg_buffer_9262 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_30218) ) ;
    buf_clk new_AGEMA_reg_buffer_9265 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T15), .Q (new_AGEMA_signal_30221) ) ;
    buf_clk new_AGEMA_reg_buffer_9268 ( .C (clk), .D (new_AGEMA_signal_6622), .Q (new_AGEMA_signal_30224) ) ;
    buf_clk new_AGEMA_reg_buffer_9271 ( .C (clk), .D (new_AGEMA_signal_6623), .Q (new_AGEMA_signal_30227) ) ;
    buf_clk new_AGEMA_reg_buffer_9274 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_30230) ) ;
    buf_clk new_AGEMA_reg_buffer_9277 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T27), .Q (new_AGEMA_signal_30233) ) ;
    buf_clk new_AGEMA_reg_buffer_9280 ( .C (clk), .D (new_AGEMA_signal_6634), .Q (new_AGEMA_signal_30236) ) ;
    buf_clk new_AGEMA_reg_buffer_9283 ( .C (clk), .D (new_AGEMA_signal_6635), .Q (new_AGEMA_signal_30239) ) ;
    buf_clk new_AGEMA_reg_buffer_9286 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_30242) ) ;
    buf_clk new_AGEMA_reg_buffer_9289 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T10), .Q (new_AGEMA_signal_30245) ) ;
    buf_clk new_AGEMA_reg_buffer_9292 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_30248) ) ;
    buf_clk new_AGEMA_reg_buffer_9295 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_30251) ) ;
    buf_clk new_AGEMA_reg_buffer_9298 ( .C (clk), .D (new_AGEMA_signal_7293), .Q (new_AGEMA_signal_30254) ) ;
    buf_clk new_AGEMA_reg_buffer_9301 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T13), .Q (new_AGEMA_signal_30257) ) ;
    buf_clk new_AGEMA_reg_buffer_9304 ( .C (clk), .D (new_AGEMA_signal_6619), .Q (new_AGEMA_signal_30260) ) ;
    buf_clk new_AGEMA_reg_buffer_9307 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_30263) ) ;
    buf_clk new_AGEMA_reg_buffer_9310 ( .C (clk), .D (new_AGEMA_signal_6621), .Q (new_AGEMA_signal_30266) ) ;
    buf_clk new_AGEMA_reg_buffer_9313 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T23), .Q (new_AGEMA_signal_30269) ) ;
    buf_clk new_AGEMA_reg_buffer_9316 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_30272) ) ;
    buf_clk new_AGEMA_reg_buffer_9319 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_30275) ) ;
    buf_clk new_AGEMA_reg_buffer_9322 ( .C (clk), .D (new_AGEMA_signal_7305), .Q (new_AGEMA_signal_30278) ) ;
    buf_clk new_AGEMA_reg_buffer_9325 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T19), .Q (new_AGEMA_signal_30281) ) ;
    buf_clk new_AGEMA_reg_buffer_9328 ( .C (clk), .D (new_AGEMA_signal_6628), .Q (new_AGEMA_signal_30284) ) ;
    buf_clk new_AGEMA_reg_buffer_9331 ( .C (clk), .D (new_AGEMA_signal_6629), .Q (new_AGEMA_signal_30287) ) ;
    buf_clk new_AGEMA_reg_buffer_9334 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_30290) ) ;
    buf_clk new_AGEMA_reg_buffer_9337 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T3), .Q (new_AGEMA_signal_30293) ) ;
    buf_clk new_AGEMA_reg_buffer_9340 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_30296) ) ;
    buf_clk new_AGEMA_reg_buffer_9343 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_30299) ) ;
    buf_clk new_AGEMA_reg_buffer_9346 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_30302) ) ;
    buf_clk new_AGEMA_reg_buffer_9349 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T22), .Q (new_AGEMA_signal_30305) ) ;
    buf_clk new_AGEMA_reg_buffer_9352 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_30308) ) ;
    buf_clk new_AGEMA_reg_buffer_9355 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_30311) ) ;
    buf_clk new_AGEMA_reg_buffer_9358 ( .C (clk), .D (new_AGEMA_signal_6633), .Q (new_AGEMA_signal_30314) ) ;
    buf_clk new_AGEMA_reg_buffer_9361 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T20), .Q (new_AGEMA_signal_30317) ) ;
    buf_clk new_AGEMA_reg_buffer_9364 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_30320) ) ;
    buf_clk new_AGEMA_reg_buffer_9367 ( .C (clk), .D (new_AGEMA_signal_7301), .Q (new_AGEMA_signal_30323) ) ;
    buf_clk new_AGEMA_reg_buffer_9370 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_30326) ) ;
    buf_clk new_AGEMA_reg_buffer_9373 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T1), .Q (new_AGEMA_signal_30329) ) ;
    buf_clk new_AGEMA_reg_buffer_9376 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_30332) ) ;
    buf_clk new_AGEMA_reg_buffer_9379 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_30335) ) ;
    buf_clk new_AGEMA_reg_buffer_9382 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_30338) ) ;
    buf_clk new_AGEMA_reg_buffer_9385 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T4), .Q (new_AGEMA_signal_30341) ) ;
    buf_clk new_AGEMA_reg_buffer_9388 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_30344) ) ;
    buf_clk new_AGEMA_reg_buffer_9391 ( .C (clk), .D (new_AGEMA_signal_6101), .Q (new_AGEMA_signal_30347) ) ;
    buf_clk new_AGEMA_reg_buffer_9394 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_30350) ) ;
    buf_clk new_AGEMA_reg_buffer_9397 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T2), .Q (new_AGEMA_signal_30353) ) ;
    buf_clk new_AGEMA_reg_buffer_9400 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_30356) ) ;
    buf_clk new_AGEMA_reg_buffer_9403 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_30359) ) ;
    buf_clk new_AGEMA_reg_buffer_9406 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_30362) ) ;
    buf_clk new_AGEMA_reg_buffer_9409 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T6), .Q (new_AGEMA_signal_30365) ) ;
    buf_clk new_AGEMA_reg_buffer_9412 ( .C (clk), .D (new_AGEMA_signal_6637), .Q (new_AGEMA_signal_30368) ) ;
    buf_clk new_AGEMA_reg_buffer_9415 ( .C (clk), .D (new_AGEMA_signal_6638), .Q (new_AGEMA_signal_30371) ) ;
    buf_clk new_AGEMA_reg_buffer_9418 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_30374) ) ;
    buf_clk new_AGEMA_reg_buffer_9421 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T8), .Q (new_AGEMA_signal_30377) ) ;
    buf_clk new_AGEMA_reg_buffer_9424 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_30380) ) ;
    buf_clk new_AGEMA_reg_buffer_9427 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_30383) ) ;
    buf_clk new_AGEMA_reg_buffer_9430 ( .C (clk), .D (new_AGEMA_signal_7329), .Q (new_AGEMA_signal_30386) ) ;
    buf_clk new_AGEMA_reg_buffer_9433 ( .C (clk), .D (ciphertext_s0[80]), .Q (new_AGEMA_signal_30389) ) ;
    buf_clk new_AGEMA_reg_buffer_9436 ( .C (clk), .D (ciphertext_s1[80]), .Q (new_AGEMA_signal_30392) ) ;
    buf_clk new_AGEMA_reg_buffer_9439 ( .C (clk), .D (ciphertext_s2[80]), .Q (new_AGEMA_signal_30395) ) ;
    buf_clk new_AGEMA_reg_buffer_9442 ( .C (clk), .D (ciphertext_s3[80]), .Q (new_AGEMA_signal_30398) ) ;
    buf_clk new_AGEMA_reg_buffer_9445 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T16), .Q (new_AGEMA_signal_30401) ) ;
    buf_clk new_AGEMA_reg_buffer_9448 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_30404) ) ;
    buf_clk new_AGEMA_reg_buffer_9451 ( .C (clk), .D (new_AGEMA_signal_6650), .Q (new_AGEMA_signal_30407) ) ;
    buf_clk new_AGEMA_reg_buffer_9454 ( .C (clk), .D (new_AGEMA_signal_6651), .Q (new_AGEMA_signal_30410) ) ;
    buf_clk new_AGEMA_reg_buffer_9457 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T9), .Q (new_AGEMA_signal_30413) ) ;
    buf_clk new_AGEMA_reg_buffer_9460 ( .C (clk), .D (new_AGEMA_signal_6640), .Q (new_AGEMA_signal_30416) ) ;
    buf_clk new_AGEMA_reg_buffer_9463 ( .C (clk), .D (new_AGEMA_signal_6641), .Q (new_AGEMA_signal_30419) ) ;
    buf_clk new_AGEMA_reg_buffer_9466 ( .C (clk), .D (new_AGEMA_signal_6642), .Q (new_AGEMA_signal_30422) ) ;
    buf_clk new_AGEMA_reg_buffer_9469 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T17), .Q (new_AGEMA_signal_30425) ) ;
    buf_clk new_AGEMA_reg_buffer_9472 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_30428) ) ;
    buf_clk new_AGEMA_reg_buffer_9475 ( .C (clk), .D (new_AGEMA_signal_7337), .Q (new_AGEMA_signal_30431) ) ;
    buf_clk new_AGEMA_reg_buffer_9478 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_30434) ) ;
    buf_clk new_AGEMA_reg_buffer_9481 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T15), .Q (new_AGEMA_signal_30437) ) ;
    buf_clk new_AGEMA_reg_buffer_9484 ( .C (clk), .D (new_AGEMA_signal_6646), .Q (new_AGEMA_signal_30440) ) ;
    buf_clk new_AGEMA_reg_buffer_9487 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_30443) ) ;
    buf_clk new_AGEMA_reg_buffer_9490 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_30446) ) ;
    buf_clk new_AGEMA_reg_buffer_9493 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T27), .Q (new_AGEMA_signal_30449) ) ;
    buf_clk new_AGEMA_reg_buffer_9496 ( .C (clk), .D (new_AGEMA_signal_6658), .Q (new_AGEMA_signal_30452) ) ;
    buf_clk new_AGEMA_reg_buffer_9499 ( .C (clk), .D (new_AGEMA_signal_6659), .Q (new_AGEMA_signal_30455) ) ;
    buf_clk new_AGEMA_reg_buffer_9502 ( .C (clk), .D (new_AGEMA_signal_6660), .Q (new_AGEMA_signal_30458) ) ;
    buf_clk new_AGEMA_reg_buffer_9505 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T10), .Q (new_AGEMA_signal_30461) ) ;
    buf_clk new_AGEMA_reg_buffer_9508 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_30464) ) ;
    buf_clk new_AGEMA_reg_buffer_9511 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_30467) ) ;
    buf_clk new_AGEMA_reg_buffer_9514 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_30470) ) ;
    buf_clk new_AGEMA_reg_buffer_9517 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T13), .Q (new_AGEMA_signal_30473) ) ;
    buf_clk new_AGEMA_reg_buffer_9520 ( .C (clk), .D (new_AGEMA_signal_6643), .Q (new_AGEMA_signal_30476) ) ;
    buf_clk new_AGEMA_reg_buffer_9523 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_30479) ) ;
    buf_clk new_AGEMA_reg_buffer_9526 ( .C (clk), .D (new_AGEMA_signal_6645), .Q (new_AGEMA_signal_30482) ) ;
    buf_clk new_AGEMA_reg_buffer_9529 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T23), .Q (new_AGEMA_signal_30485) ) ;
    buf_clk new_AGEMA_reg_buffer_9532 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_30488) ) ;
    buf_clk new_AGEMA_reg_buffer_9535 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_30491) ) ;
    buf_clk new_AGEMA_reg_buffer_9538 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_30494) ) ;
    buf_clk new_AGEMA_reg_buffer_9541 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T19), .Q (new_AGEMA_signal_30497) ) ;
    buf_clk new_AGEMA_reg_buffer_9544 ( .C (clk), .D (new_AGEMA_signal_6652), .Q (new_AGEMA_signal_30500) ) ;
    buf_clk new_AGEMA_reg_buffer_9547 ( .C (clk), .D (new_AGEMA_signal_6653), .Q (new_AGEMA_signal_30503) ) ;
    buf_clk new_AGEMA_reg_buffer_9550 ( .C (clk), .D (new_AGEMA_signal_6654), .Q (new_AGEMA_signal_30506) ) ;
    buf_clk new_AGEMA_reg_buffer_9553 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T3), .Q (new_AGEMA_signal_30509) ) ;
    buf_clk new_AGEMA_reg_buffer_9556 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_30512) ) ;
    buf_clk new_AGEMA_reg_buffer_9559 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_30515) ) ;
    buf_clk new_AGEMA_reg_buffer_9562 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_30518) ) ;
    buf_clk new_AGEMA_reg_buffer_9565 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T22), .Q (new_AGEMA_signal_30521) ) ;
    buf_clk new_AGEMA_reg_buffer_9568 ( .C (clk), .D (new_AGEMA_signal_6655), .Q (new_AGEMA_signal_30524) ) ;
    buf_clk new_AGEMA_reg_buffer_9571 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_30527) ) ;
    buf_clk new_AGEMA_reg_buffer_9574 ( .C (clk), .D (new_AGEMA_signal_6657), .Q (new_AGEMA_signal_30530) ) ;
    buf_clk new_AGEMA_reg_buffer_9577 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T20), .Q (new_AGEMA_signal_30533) ) ;
    buf_clk new_AGEMA_reg_buffer_9580 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_30536) ) ;
    buf_clk new_AGEMA_reg_buffer_9583 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_30539) ) ;
    buf_clk new_AGEMA_reg_buffer_9586 ( .C (clk), .D (new_AGEMA_signal_7341), .Q (new_AGEMA_signal_30542) ) ;
    buf_clk new_AGEMA_reg_buffer_9589 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T1), .Q (new_AGEMA_signal_30545) ) ;
    buf_clk new_AGEMA_reg_buffer_9592 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_30548) ) ;
    buf_clk new_AGEMA_reg_buffer_9595 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_30551) ) ;
    buf_clk new_AGEMA_reg_buffer_9598 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_30554) ) ;
    buf_clk new_AGEMA_reg_buffer_9601 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T4), .Q (new_AGEMA_signal_30557) ) ;
    buf_clk new_AGEMA_reg_buffer_9604 ( .C (clk), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_30560) ) ;
    buf_clk new_AGEMA_reg_buffer_9607 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_30563) ) ;
    buf_clk new_AGEMA_reg_buffer_9610 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_30566) ) ;
    buf_clk new_AGEMA_reg_buffer_9613 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T2), .Q (new_AGEMA_signal_30569) ) ;
    buf_clk new_AGEMA_reg_buffer_9616 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_30572) ) ;
    buf_clk new_AGEMA_reg_buffer_9619 ( .C (clk), .D (new_AGEMA_signal_6125), .Q (new_AGEMA_signal_30575) ) ;
    buf_clk new_AGEMA_reg_buffer_9622 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_30578) ) ;
    buf_clk new_AGEMA_reg_buffer_9625 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T6), .Q (new_AGEMA_signal_30581) ) ;
    buf_clk new_AGEMA_reg_buffer_9628 ( .C (clk), .D (new_AGEMA_signal_6661), .Q (new_AGEMA_signal_30584) ) ;
    buf_clk new_AGEMA_reg_buffer_9631 ( .C (clk), .D (new_AGEMA_signal_6662), .Q (new_AGEMA_signal_30587) ) ;
    buf_clk new_AGEMA_reg_buffer_9634 ( .C (clk), .D (new_AGEMA_signal_6663), .Q (new_AGEMA_signal_30590) ) ;
    buf_clk new_AGEMA_reg_buffer_9637 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T8), .Q (new_AGEMA_signal_30593) ) ;
    buf_clk new_AGEMA_reg_buffer_9640 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_30596) ) ;
    buf_clk new_AGEMA_reg_buffer_9643 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_30599) ) ;
    buf_clk new_AGEMA_reg_buffer_9646 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_30602) ) ;
    buf_clk new_AGEMA_reg_buffer_9649 ( .C (clk), .D (ciphertext_s0[88]), .Q (new_AGEMA_signal_30605) ) ;
    buf_clk new_AGEMA_reg_buffer_9652 ( .C (clk), .D (ciphertext_s1[88]), .Q (new_AGEMA_signal_30608) ) ;
    buf_clk new_AGEMA_reg_buffer_9655 ( .C (clk), .D (ciphertext_s2[88]), .Q (new_AGEMA_signal_30611) ) ;
    buf_clk new_AGEMA_reg_buffer_9658 ( .C (clk), .D (ciphertext_s3[88]), .Q (new_AGEMA_signal_30614) ) ;
    buf_clk new_AGEMA_reg_buffer_9661 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T16), .Q (new_AGEMA_signal_30617) ) ;
    buf_clk new_AGEMA_reg_buffer_9664 ( .C (clk), .D (new_AGEMA_signal_6673), .Q (new_AGEMA_signal_30620) ) ;
    buf_clk new_AGEMA_reg_buffer_9667 ( .C (clk), .D (new_AGEMA_signal_6674), .Q (new_AGEMA_signal_30623) ) ;
    buf_clk new_AGEMA_reg_buffer_9670 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_30626) ) ;
    buf_clk new_AGEMA_reg_buffer_9673 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T9), .Q (new_AGEMA_signal_30629) ) ;
    buf_clk new_AGEMA_reg_buffer_9676 ( .C (clk), .D (new_AGEMA_signal_6664), .Q (new_AGEMA_signal_30632) ) ;
    buf_clk new_AGEMA_reg_buffer_9679 ( .C (clk), .D (new_AGEMA_signal_6665), .Q (new_AGEMA_signal_30635) ) ;
    buf_clk new_AGEMA_reg_buffer_9682 ( .C (clk), .D (new_AGEMA_signal_6666), .Q (new_AGEMA_signal_30638) ) ;
    buf_clk new_AGEMA_reg_buffer_9685 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T17), .Q (new_AGEMA_signal_30641) ) ;
    buf_clk new_AGEMA_reg_buffer_9688 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_30644) ) ;
    buf_clk new_AGEMA_reg_buffer_9691 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_30647) ) ;
    buf_clk new_AGEMA_reg_buffer_9694 ( .C (clk), .D (new_AGEMA_signal_7377), .Q (new_AGEMA_signal_30650) ) ;
    buf_clk new_AGEMA_reg_buffer_9697 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T15), .Q (new_AGEMA_signal_30653) ) ;
    buf_clk new_AGEMA_reg_buffer_9700 ( .C (clk), .D (new_AGEMA_signal_6670), .Q (new_AGEMA_signal_30656) ) ;
    buf_clk new_AGEMA_reg_buffer_9703 ( .C (clk), .D (new_AGEMA_signal_6671), .Q (new_AGEMA_signal_30659) ) ;
    buf_clk new_AGEMA_reg_buffer_9706 ( .C (clk), .D (new_AGEMA_signal_6672), .Q (new_AGEMA_signal_30662) ) ;
    buf_clk new_AGEMA_reg_buffer_9709 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T27), .Q (new_AGEMA_signal_30665) ) ;
    buf_clk new_AGEMA_reg_buffer_9712 ( .C (clk), .D (new_AGEMA_signal_6682), .Q (new_AGEMA_signal_30668) ) ;
    buf_clk new_AGEMA_reg_buffer_9715 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_30671) ) ;
    buf_clk new_AGEMA_reg_buffer_9718 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_30674) ) ;
    buf_clk new_AGEMA_reg_buffer_9721 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T10), .Q (new_AGEMA_signal_30677) ) ;
    buf_clk new_AGEMA_reg_buffer_9724 ( .C (clk), .D (new_AGEMA_signal_7369), .Q (new_AGEMA_signal_30680) ) ;
    buf_clk new_AGEMA_reg_buffer_9727 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_30683) ) ;
    buf_clk new_AGEMA_reg_buffer_9730 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_30686) ) ;
    buf_clk new_AGEMA_reg_buffer_9733 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T13), .Q (new_AGEMA_signal_30689) ) ;
    buf_clk new_AGEMA_reg_buffer_9736 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_30692) ) ;
    buf_clk new_AGEMA_reg_buffer_9739 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_30695) ) ;
    buf_clk new_AGEMA_reg_buffer_9742 ( .C (clk), .D (new_AGEMA_signal_6669), .Q (new_AGEMA_signal_30698) ) ;
    buf_clk new_AGEMA_reg_buffer_9745 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T23), .Q (new_AGEMA_signal_30701) ) ;
    buf_clk new_AGEMA_reg_buffer_9748 ( .C (clk), .D (new_AGEMA_signal_7381), .Q (new_AGEMA_signal_30704) ) ;
    buf_clk new_AGEMA_reg_buffer_9751 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_30707) ) ;
    buf_clk new_AGEMA_reg_buffer_9754 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_30710) ) ;
    buf_clk new_AGEMA_reg_buffer_9757 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T19), .Q (new_AGEMA_signal_30713) ) ;
    buf_clk new_AGEMA_reg_buffer_9760 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_30716) ) ;
    buf_clk new_AGEMA_reg_buffer_9763 ( .C (clk), .D (new_AGEMA_signal_6677), .Q (new_AGEMA_signal_30719) ) ;
    buf_clk new_AGEMA_reg_buffer_9766 ( .C (clk), .D (new_AGEMA_signal_6678), .Q (new_AGEMA_signal_30722) ) ;
    buf_clk new_AGEMA_reg_buffer_9769 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T3), .Q (new_AGEMA_signal_30725) ) ;
    buf_clk new_AGEMA_reg_buffer_9772 ( .C (clk), .D (new_AGEMA_signal_6157), .Q (new_AGEMA_signal_30728) ) ;
    buf_clk new_AGEMA_reg_buffer_9775 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_30731) ) ;
    buf_clk new_AGEMA_reg_buffer_9778 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_30734) ) ;
    buf_clk new_AGEMA_reg_buffer_9781 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T22), .Q (new_AGEMA_signal_30737) ) ;
    buf_clk new_AGEMA_reg_buffer_9784 ( .C (clk), .D (new_AGEMA_signal_6679), .Q (new_AGEMA_signal_30740) ) ;
    buf_clk new_AGEMA_reg_buffer_9787 ( .C (clk), .D (new_AGEMA_signal_6680), .Q (new_AGEMA_signal_30743) ) ;
    buf_clk new_AGEMA_reg_buffer_9790 ( .C (clk), .D (new_AGEMA_signal_6681), .Q (new_AGEMA_signal_30746) ) ;
    buf_clk new_AGEMA_reg_buffer_9793 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T20), .Q (new_AGEMA_signal_30749) ) ;
    buf_clk new_AGEMA_reg_buffer_9796 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_30752) ) ;
    buf_clk new_AGEMA_reg_buffer_9799 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_30755) ) ;
    buf_clk new_AGEMA_reg_buffer_9802 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_30758) ) ;
    buf_clk new_AGEMA_reg_buffer_9805 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T1), .Q (new_AGEMA_signal_30761) ) ;
    buf_clk new_AGEMA_reg_buffer_9808 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_30764) ) ;
    buf_clk new_AGEMA_reg_buffer_9811 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_30767) ) ;
    buf_clk new_AGEMA_reg_buffer_9814 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_30770) ) ;
    buf_clk new_AGEMA_reg_buffer_9817 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T4), .Q (new_AGEMA_signal_30773) ) ;
    buf_clk new_AGEMA_reg_buffer_9820 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_30776) ) ;
    buf_clk new_AGEMA_reg_buffer_9823 ( .C (clk), .D (new_AGEMA_signal_6161), .Q (new_AGEMA_signal_30779) ) ;
    buf_clk new_AGEMA_reg_buffer_9826 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_30782) ) ;
    buf_clk new_AGEMA_reg_buffer_9829 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T2), .Q (new_AGEMA_signal_30785) ) ;
    buf_clk new_AGEMA_reg_buffer_9832 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_30788) ) ;
    buf_clk new_AGEMA_reg_buffer_9835 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_30791) ) ;
    buf_clk new_AGEMA_reg_buffer_9838 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_30794) ) ;
    buf_clk new_AGEMA_reg_buffer_9841 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T6), .Q (new_AGEMA_signal_30797) ) ;
    buf_clk new_AGEMA_reg_buffer_9844 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_30800) ) ;
    buf_clk new_AGEMA_reg_buffer_9847 ( .C (clk), .D (new_AGEMA_signal_6686), .Q (new_AGEMA_signal_30803) ) ;
    buf_clk new_AGEMA_reg_buffer_9850 ( .C (clk), .D (new_AGEMA_signal_6687), .Q (new_AGEMA_signal_30806) ) ;
    buf_clk new_AGEMA_reg_buffer_9853 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T8), .Q (new_AGEMA_signal_30809) ) ;
    buf_clk new_AGEMA_reg_buffer_9856 ( .C (clk), .D (new_AGEMA_signal_7405), .Q (new_AGEMA_signal_30812) ) ;
    buf_clk new_AGEMA_reg_buffer_9859 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_30815) ) ;
    buf_clk new_AGEMA_reg_buffer_9862 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_30818) ) ;
    buf_clk new_AGEMA_reg_buffer_9865 ( .C (clk), .D (ciphertext_s0[96]), .Q (new_AGEMA_signal_30821) ) ;
    buf_clk new_AGEMA_reg_buffer_9868 ( .C (clk), .D (ciphertext_s1[96]), .Q (new_AGEMA_signal_30824) ) ;
    buf_clk new_AGEMA_reg_buffer_9871 ( .C (clk), .D (ciphertext_s2[96]), .Q (new_AGEMA_signal_30827) ) ;
    buf_clk new_AGEMA_reg_buffer_9874 ( .C (clk), .D (ciphertext_s3[96]), .Q (new_AGEMA_signal_30830) ) ;
    buf_clk new_AGEMA_reg_buffer_9877 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T16), .Q (new_AGEMA_signal_30833) ) ;
    buf_clk new_AGEMA_reg_buffer_9880 ( .C (clk), .D (new_AGEMA_signal_6697), .Q (new_AGEMA_signal_30836) ) ;
    buf_clk new_AGEMA_reg_buffer_9883 ( .C (clk), .D (new_AGEMA_signal_6698), .Q (new_AGEMA_signal_30839) ) ;
    buf_clk new_AGEMA_reg_buffer_9886 ( .C (clk), .D (new_AGEMA_signal_6699), .Q (new_AGEMA_signal_30842) ) ;
    buf_clk new_AGEMA_reg_buffer_9889 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T9), .Q (new_AGEMA_signal_30845) ) ;
    buf_clk new_AGEMA_reg_buffer_9892 ( .C (clk), .D (new_AGEMA_signal_6688), .Q (new_AGEMA_signal_30848) ) ;
    buf_clk new_AGEMA_reg_buffer_9895 ( .C (clk), .D (new_AGEMA_signal_6689), .Q (new_AGEMA_signal_30851) ) ;
    buf_clk new_AGEMA_reg_buffer_9898 ( .C (clk), .D (new_AGEMA_signal_6690), .Q (new_AGEMA_signal_30854) ) ;
    buf_clk new_AGEMA_reg_buffer_9901 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T17), .Q (new_AGEMA_signal_30857) ) ;
    buf_clk new_AGEMA_reg_buffer_9904 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_30860) ) ;
    buf_clk new_AGEMA_reg_buffer_9907 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_30863) ) ;
    buf_clk new_AGEMA_reg_buffer_9910 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_30866) ) ;
    buf_clk new_AGEMA_reg_buffer_9913 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T15), .Q (new_AGEMA_signal_30869) ) ;
    buf_clk new_AGEMA_reg_buffer_9916 ( .C (clk), .D (new_AGEMA_signal_6694), .Q (new_AGEMA_signal_30872) ) ;
    buf_clk new_AGEMA_reg_buffer_9919 ( .C (clk), .D (new_AGEMA_signal_6695), .Q (new_AGEMA_signal_30875) ) ;
    buf_clk new_AGEMA_reg_buffer_9922 ( .C (clk), .D (new_AGEMA_signal_6696), .Q (new_AGEMA_signal_30878) ) ;
    buf_clk new_AGEMA_reg_buffer_9925 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T27), .Q (new_AGEMA_signal_30881) ) ;
    buf_clk new_AGEMA_reg_buffer_9928 ( .C (clk), .D (new_AGEMA_signal_6706), .Q (new_AGEMA_signal_30884) ) ;
    buf_clk new_AGEMA_reg_buffer_9931 ( .C (clk), .D (new_AGEMA_signal_6707), .Q (new_AGEMA_signal_30887) ) ;
    buf_clk new_AGEMA_reg_buffer_9934 ( .C (clk), .D (new_AGEMA_signal_6708), .Q (new_AGEMA_signal_30890) ) ;
    buf_clk new_AGEMA_reg_buffer_9937 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T10), .Q (new_AGEMA_signal_30893) ) ;
    buf_clk new_AGEMA_reg_buffer_9940 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_30896) ) ;
    buf_clk new_AGEMA_reg_buffer_9943 ( .C (clk), .D (new_AGEMA_signal_7409), .Q (new_AGEMA_signal_30899) ) ;
    buf_clk new_AGEMA_reg_buffer_9946 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_30902) ) ;
    buf_clk new_AGEMA_reg_buffer_9949 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T13), .Q (new_AGEMA_signal_30905) ) ;
    buf_clk new_AGEMA_reg_buffer_9952 ( .C (clk), .D (new_AGEMA_signal_6691), .Q (new_AGEMA_signal_30908) ) ;
    buf_clk new_AGEMA_reg_buffer_9955 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_30911) ) ;
    buf_clk new_AGEMA_reg_buffer_9958 ( .C (clk), .D (new_AGEMA_signal_6693), .Q (new_AGEMA_signal_30914) ) ;
    buf_clk new_AGEMA_reg_buffer_9961 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T23), .Q (new_AGEMA_signal_30917) ) ;
    buf_clk new_AGEMA_reg_buffer_9964 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_30920) ) ;
    buf_clk new_AGEMA_reg_buffer_9967 ( .C (clk), .D (new_AGEMA_signal_7421), .Q (new_AGEMA_signal_30923) ) ;
    buf_clk new_AGEMA_reg_buffer_9970 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_30926) ) ;
    buf_clk new_AGEMA_reg_buffer_9973 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T19), .Q (new_AGEMA_signal_30929) ) ;
    buf_clk new_AGEMA_reg_buffer_9976 ( .C (clk), .D (new_AGEMA_signal_6700), .Q (new_AGEMA_signal_30932) ) ;
    buf_clk new_AGEMA_reg_buffer_9979 ( .C (clk), .D (new_AGEMA_signal_6701), .Q (new_AGEMA_signal_30935) ) ;
    buf_clk new_AGEMA_reg_buffer_9982 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_30938) ) ;
    buf_clk new_AGEMA_reg_buffer_9985 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T3), .Q (new_AGEMA_signal_30941) ) ;
    buf_clk new_AGEMA_reg_buffer_9988 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_30944) ) ;
    buf_clk new_AGEMA_reg_buffer_9991 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_30947) ) ;
    buf_clk new_AGEMA_reg_buffer_9994 ( .C (clk), .D (new_AGEMA_signal_6189), .Q (new_AGEMA_signal_30950) ) ;
    buf_clk new_AGEMA_reg_buffer_9997 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T22), .Q (new_AGEMA_signal_30953) ) ;
    buf_clk new_AGEMA_reg_buffer_10000 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_30956) ) ;
    buf_clk new_AGEMA_reg_buffer_10003 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_30959) ) ;
    buf_clk new_AGEMA_reg_buffer_10006 ( .C (clk), .D (new_AGEMA_signal_6705), .Q (new_AGEMA_signal_30962) ) ;
    buf_clk new_AGEMA_reg_buffer_10009 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T20), .Q (new_AGEMA_signal_30965) ) ;
    buf_clk new_AGEMA_reg_buffer_10012 ( .C (clk), .D (new_AGEMA_signal_7417), .Q (new_AGEMA_signal_30968) ) ;
    buf_clk new_AGEMA_reg_buffer_10015 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_30971) ) ;
    buf_clk new_AGEMA_reg_buffer_10018 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_30974) ) ;
    buf_clk new_AGEMA_reg_buffer_10021 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T1), .Q (new_AGEMA_signal_30977) ) ;
    buf_clk new_AGEMA_reg_buffer_10024 ( .C (clk), .D (new_AGEMA_signal_6181), .Q (new_AGEMA_signal_30980) ) ;
    buf_clk new_AGEMA_reg_buffer_10027 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_30983) ) ;
    buf_clk new_AGEMA_reg_buffer_10030 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_30986) ) ;
    buf_clk new_AGEMA_reg_buffer_10033 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T4), .Q (new_AGEMA_signal_30989) ) ;
    buf_clk new_AGEMA_reg_buffer_10036 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_30992) ) ;
    buf_clk new_AGEMA_reg_buffer_10039 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_30995) ) ;
    buf_clk new_AGEMA_reg_buffer_10042 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_30998) ) ;
    buf_clk new_AGEMA_reg_buffer_10045 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T2), .Q (new_AGEMA_signal_31001) ) ;
    buf_clk new_AGEMA_reg_buffer_10048 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_31004) ) ;
    buf_clk new_AGEMA_reg_buffer_10051 ( .C (clk), .D (new_AGEMA_signal_6185), .Q (new_AGEMA_signal_31007) ) ;
    buf_clk new_AGEMA_reg_buffer_10054 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_31010) ) ;
    buf_clk new_AGEMA_reg_buffer_10057 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T6), .Q (new_AGEMA_signal_31013) ) ;
    buf_clk new_AGEMA_reg_buffer_10060 ( .C (clk), .D (new_AGEMA_signal_6709), .Q (new_AGEMA_signal_31016) ) ;
    buf_clk new_AGEMA_reg_buffer_10063 ( .C (clk), .D (new_AGEMA_signal_6710), .Q (new_AGEMA_signal_31019) ) ;
    buf_clk new_AGEMA_reg_buffer_10066 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_31022) ) ;
    buf_clk new_AGEMA_reg_buffer_10069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T8), .Q (new_AGEMA_signal_31025) ) ;
    buf_clk new_AGEMA_reg_buffer_10072 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_31028) ) ;
    buf_clk new_AGEMA_reg_buffer_10075 ( .C (clk), .D (new_AGEMA_signal_7445), .Q (new_AGEMA_signal_31031) ) ;
    buf_clk new_AGEMA_reg_buffer_10078 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_31034) ) ;
    buf_clk new_AGEMA_reg_buffer_10081 ( .C (clk), .D (ciphertext_s0[104]), .Q (new_AGEMA_signal_31037) ) ;
    buf_clk new_AGEMA_reg_buffer_10084 ( .C (clk), .D (ciphertext_s1[104]), .Q (new_AGEMA_signal_31040) ) ;
    buf_clk new_AGEMA_reg_buffer_10087 ( .C (clk), .D (ciphertext_s2[104]), .Q (new_AGEMA_signal_31043) ) ;
    buf_clk new_AGEMA_reg_buffer_10090 ( .C (clk), .D (ciphertext_s3[104]), .Q (new_AGEMA_signal_31046) ) ;
    buf_clk new_AGEMA_reg_buffer_10093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T16), .Q (new_AGEMA_signal_31049) ) ;
    buf_clk new_AGEMA_reg_buffer_10096 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_31052) ) ;
    buf_clk new_AGEMA_reg_buffer_10099 ( .C (clk), .D (new_AGEMA_signal_6722), .Q (new_AGEMA_signal_31055) ) ;
    buf_clk new_AGEMA_reg_buffer_10102 ( .C (clk), .D (new_AGEMA_signal_6723), .Q (new_AGEMA_signal_31058) ) ;
    buf_clk new_AGEMA_reg_buffer_10105 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T9), .Q (new_AGEMA_signal_31061) ) ;
    buf_clk new_AGEMA_reg_buffer_10108 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_31064) ) ;
    buf_clk new_AGEMA_reg_buffer_10111 ( .C (clk), .D (new_AGEMA_signal_6713), .Q (new_AGEMA_signal_31067) ) ;
    buf_clk new_AGEMA_reg_buffer_10114 ( .C (clk), .D (new_AGEMA_signal_6714), .Q (new_AGEMA_signal_31070) ) ;
    buf_clk new_AGEMA_reg_buffer_10117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T17), .Q (new_AGEMA_signal_31073) ) ;
    buf_clk new_AGEMA_reg_buffer_10120 ( .C (clk), .D (new_AGEMA_signal_7453), .Q (new_AGEMA_signal_31076) ) ;
    buf_clk new_AGEMA_reg_buffer_10123 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_31079) ) ;
    buf_clk new_AGEMA_reg_buffer_10126 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_31082) ) ;
    buf_clk new_AGEMA_reg_buffer_10129 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T15), .Q (new_AGEMA_signal_31085) ) ;
    buf_clk new_AGEMA_reg_buffer_10132 ( .C (clk), .D (new_AGEMA_signal_6718), .Q (new_AGEMA_signal_31088) ) ;
    buf_clk new_AGEMA_reg_buffer_10135 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_31091) ) ;
    buf_clk new_AGEMA_reg_buffer_10138 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_31094) ) ;
    buf_clk new_AGEMA_reg_buffer_10141 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T27), .Q (new_AGEMA_signal_31097) ) ;
    buf_clk new_AGEMA_reg_buffer_10144 ( .C (clk), .D (new_AGEMA_signal_6730), .Q (new_AGEMA_signal_31100) ) ;
    buf_clk new_AGEMA_reg_buffer_10147 ( .C (clk), .D (new_AGEMA_signal_6731), .Q (new_AGEMA_signal_31103) ) ;
    buf_clk new_AGEMA_reg_buffer_10150 ( .C (clk), .D (new_AGEMA_signal_6732), .Q (new_AGEMA_signal_31106) ) ;
    buf_clk new_AGEMA_reg_buffer_10153 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T10), .Q (new_AGEMA_signal_31109) ) ;
    buf_clk new_AGEMA_reg_buffer_10156 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_31112) ) ;
    buf_clk new_AGEMA_reg_buffer_10159 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_31115) ) ;
    buf_clk new_AGEMA_reg_buffer_10162 ( .C (clk), .D (new_AGEMA_signal_7449), .Q (new_AGEMA_signal_31118) ) ;
    buf_clk new_AGEMA_reg_buffer_10165 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T13), .Q (new_AGEMA_signal_31121) ) ;
    buf_clk new_AGEMA_reg_buffer_10168 ( .C (clk), .D (new_AGEMA_signal_6715), .Q (new_AGEMA_signal_31124) ) ;
    buf_clk new_AGEMA_reg_buffer_10171 ( .C (clk), .D (new_AGEMA_signal_6716), .Q (new_AGEMA_signal_31127) ) ;
    buf_clk new_AGEMA_reg_buffer_10174 ( .C (clk), .D (new_AGEMA_signal_6717), .Q (new_AGEMA_signal_31130) ) ;
    buf_clk new_AGEMA_reg_buffer_10177 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T23), .Q (new_AGEMA_signal_31133) ) ;
    buf_clk new_AGEMA_reg_buffer_10180 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_31136) ) ;
    buf_clk new_AGEMA_reg_buffer_10183 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_31139) ) ;
    buf_clk new_AGEMA_reg_buffer_10186 ( .C (clk), .D (new_AGEMA_signal_7461), .Q (new_AGEMA_signal_31142) ) ;
    buf_clk new_AGEMA_reg_buffer_10189 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T19), .Q (new_AGEMA_signal_31145) ) ;
    buf_clk new_AGEMA_reg_buffer_10192 ( .C (clk), .D (new_AGEMA_signal_6724), .Q (new_AGEMA_signal_31148) ) ;
    buf_clk new_AGEMA_reg_buffer_10195 ( .C (clk), .D (new_AGEMA_signal_6725), .Q (new_AGEMA_signal_31151) ) ;
    buf_clk new_AGEMA_reg_buffer_10198 ( .C (clk), .D (new_AGEMA_signal_6726), .Q (new_AGEMA_signal_31154) ) ;
    buf_clk new_AGEMA_reg_buffer_10201 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T3), .Q (new_AGEMA_signal_31157) ) ;
    buf_clk new_AGEMA_reg_buffer_10204 ( .C (clk), .D (new_AGEMA_signal_6217), .Q (new_AGEMA_signal_31160) ) ;
    buf_clk new_AGEMA_reg_buffer_10207 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_31163) ) ;
    buf_clk new_AGEMA_reg_buffer_10210 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_31166) ) ;
    buf_clk new_AGEMA_reg_buffer_10213 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T22), .Q (new_AGEMA_signal_31169) ) ;
    buf_clk new_AGEMA_reg_buffer_10216 ( .C (clk), .D (new_AGEMA_signal_6727), .Q (new_AGEMA_signal_31172) ) ;
    buf_clk new_AGEMA_reg_buffer_10219 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_31175) ) ;
    buf_clk new_AGEMA_reg_buffer_10222 ( .C (clk), .D (new_AGEMA_signal_6729), .Q (new_AGEMA_signal_31178) ) ;
    buf_clk new_AGEMA_reg_buffer_10225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T20), .Q (new_AGEMA_signal_31181) ) ;
    buf_clk new_AGEMA_reg_buffer_10228 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_31184) ) ;
    buf_clk new_AGEMA_reg_buffer_10231 ( .C (clk), .D (new_AGEMA_signal_7457), .Q (new_AGEMA_signal_31187) ) ;
    buf_clk new_AGEMA_reg_buffer_10234 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_31190) ) ;
    buf_clk new_AGEMA_reg_buffer_10237 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T1), .Q (new_AGEMA_signal_31193) ) ;
    buf_clk new_AGEMA_reg_buffer_10240 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_31196) ) ;
    buf_clk new_AGEMA_reg_buffer_10243 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_31199) ) ;
    buf_clk new_AGEMA_reg_buffer_10246 ( .C (clk), .D (new_AGEMA_signal_6213), .Q (new_AGEMA_signal_31202) ) ;
    buf_clk new_AGEMA_reg_buffer_10249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T4), .Q (new_AGEMA_signal_31205) ) ;
    buf_clk new_AGEMA_reg_buffer_10252 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_31208) ) ;
    buf_clk new_AGEMA_reg_buffer_10255 ( .C (clk), .D (new_AGEMA_signal_6221), .Q (new_AGEMA_signal_31211) ) ;
    buf_clk new_AGEMA_reg_buffer_10258 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_31214) ) ;
    buf_clk new_AGEMA_reg_buffer_10261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T2), .Q (new_AGEMA_signal_31217) ) ;
    buf_clk new_AGEMA_reg_buffer_10264 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_31220) ) ;
    buf_clk new_AGEMA_reg_buffer_10267 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_31223) ) ;
    buf_clk new_AGEMA_reg_buffer_10270 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_31226) ) ;
    buf_clk new_AGEMA_reg_buffer_10273 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T6), .Q (new_AGEMA_signal_31229) ) ;
    buf_clk new_AGEMA_reg_buffer_10276 ( .C (clk), .D (new_AGEMA_signal_6733), .Q (new_AGEMA_signal_31232) ) ;
    buf_clk new_AGEMA_reg_buffer_10279 ( .C (clk), .D (new_AGEMA_signal_6734), .Q (new_AGEMA_signal_31235) ) ;
    buf_clk new_AGEMA_reg_buffer_10282 ( .C (clk), .D (new_AGEMA_signal_6735), .Q (new_AGEMA_signal_31238) ) ;
    buf_clk new_AGEMA_reg_buffer_10285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T8), .Q (new_AGEMA_signal_31241) ) ;
    buf_clk new_AGEMA_reg_buffer_10288 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_31244) ) ;
    buf_clk new_AGEMA_reg_buffer_10291 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_31247) ) ;
    buf_clk new_AGEMA_reg_buffer_10294 ( .C (clk), .D (new_AGEMA_signal_7485), .Q (new_AGEMA_signal_31250) ) ;
    buf_clk new_AGEMA_reg_buffer_10297 ( .C (clk), .D (ciphertext_s0[112]), .Q (new_AGEMA_signal_31253) ) ;
    buf_clk new_AGEMA_reg_buffer_10300 ( .C (clk), .D (ciphertext_s1[112]), .Q (new_AGEMA_signal_31256) ) ;
    buf_clk new_AGEMA_reg_buffer_10303 ( .C (clk), .D (ciphertext_s2[112]), .Q (new_AGEMA_signal_31259) ) ;
    buf_clk new_AGEMA_reg_buffer_10306 ( .C (clk), .D (ciphertext_s3[112]), .Q (new_AGEMA_signal_31262) ) ;
    buf_clk new_AGEMA_reg_buffer_10309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T16), .Q (new_AGEMA_signal_31265) ) ;
    buf_clk new_AGEMA_reg_buffer_10312 ( .C (clk), .D (new_AGEMA_signal_6745), .Q (new_AGEMA_signal_31268) ) ;
    buf_clk new_AGEMA_reg_buffer_10315 ( .C (clk), .D (new_AGEMA_signal_6746), .Q (new_AGEMA_signal_31271) ) ;
    buf_clk new_AGEMA_reg_buffer_10318 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_31274) ) ;
    buf_clk new_AGEMA_reg_buffer_10321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T9), .Q (new_AGEMA_signal_31277) ) ;
    buf_clk new_AGEMA_reg_buffer_10324 ( .C (clk), .D (new_AGEMA_signal_6736), .Q (new_AGEMA_signal_31280) ) ;
    buf_clk new_AGEMA_reg_buffer_10327 ( .C (clk), .D (new_AGEMA_signal_6737), .Q (new_AGEMA_signal_31283) ) ;
    buf_clk new_AGEMA_reg_buffer_10330 ( .C (clk), .D (new_AGEMA_signal_6738), .Q (new_AGEMA_signal_31286) ) ;
    buf_clk new_AGEMA_reg_buffer_10333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T17), .Q (new_AGEMA_signal_31289) ) ;
    buf_clk new_AGEMA_reg_buffer_10336 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_31292) ) ;
    buf_clk new_AGEMA_reg_buffer_10339 ( .C (clk), .D (new_AGEMA_signal_7493), .Q (new_AGEMA_signal_31295) ) ;
    buf_clk new_AGEMA_reg_buffer_10342 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_31298) ) ;
    buf_clk new_AGEMA_reg_buffer_10345 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T15), .Q (new_AGEMA_signal_31301) ) ;
    buf_clk new_AGEMA_reg_buffer_10348 ( .C (clk), .D (new_AGEMA_signal_6742), .Q (new_AGEMA_signal_31304) ) ;
    buf_clk new_AGEMA_reg_buffer_10351 ( .C (clk), .D (new_AGEMA_signal_6743), .Q (new_AGEMA_signal_31307) ) ;
    buf_clk new_AGEMA_reg_buffer_10354 ( .C (clk), .D (new_AGEMA_signal_6744), .Q (new_AGEMA_signal_31310) ) ;
    buf_clk new_AGEMA_reg_buffer_10357 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T27), .Q (new_AGEMA_signal_31313) ) ;
    buf_clk new_AGEMA_reg_buffer_10360 ( .C (clk), .D (new_AGEMA_signal_6754), .Q (new_AGEMA_signal_31316) ) ;
    buf_clk new_AGEMA_reg_buffer_10363 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_31319) ) ;
    buf_clk new_AGEMA_reg_buffer_10366 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_31322) ) ;
    buf_clk new_AGEMA_reg_buffer_10369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T10), .Q (new_AGEMA_signal_31325) ) ;
    buf_clk new_AGEMA_reg_buffer_10372 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_31328) ) ;
    buf_clk new_AGEMA_reg_buffer_10375 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_31331) ) ;
    buf_clk new_AGEMA_reg_buffer_10378 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_31334) ) ;
    buf_clk new_AGEMA_reg_buffer_10381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T13), .Q (new_AGEMA_signal_31337) ) ;
    buf_clk new_AGEMA_reg_buffer_10384 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_31340) ) ;
    buf_clk new_AGEMA_reg_buffer_10387 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_31343) ) ;
    buf_clk new_AGEMA_reg_buffer_10390 ( .C (clk), .D (new_AGEMA_signal_6741), .Q (new_AGEMA_signal_31346) ) ;
    buf_clk new_AGEMA_reg_buffer_10393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T23), .Q (new_AGEMA_signal_31349) ) ;
    buf_clk new_AGEMA_reg_buffer_10396 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_31352) ) ;
    buf_clk new_AGEMA_reg_buffer_10399 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_31355) ) ;
    buf_clk new_AGEMA_reg_buffer_10402 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_31358) ) ;
    buf_clk new_AGEMA_reg_buffer_10405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T19), .Q (new_AGEMA_signal_31361) ) ;
    buf_clk new_AGEMA_reg_buffer_10408 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_31364) ) ;
    buf_clk new_AGEMA_reg_buffer_10411 ( .C (clk), .D (new_AGEMA_signal_6749), .Q (new_AGEMA_signal_31367) ) ;
    buf_clk new_AGEMA_reg_buffer_10414 ( .C (clk), .D (new_AGEMA_signal_6750), .Q (new_AGEMA_signal_31370) ) ;
    buf_clk new_AGEMA_reg_buffer_10417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T3), .Q (new_AGEMA_signal_31373) ) ;
    buf_clk new_AGEMA_reg_buffer_10420 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_31376) ) ;
    buf_clk new_AGEMA_reg_buffer_10423 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_31379) ) ;
    buf_clk new_AGEMA_reg_buffer_10426 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_31382) ) ;
    buf_clk new_AGEMA_reg_buffer_10429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T22), .Q (new_AGEMA_signal_31385) ) ;
    buf_clk new_AGEMA_reg_buffer_10432 ( .C (clk), .D (new_AGEMA_signal_6751), .Q (new_AGEMA_signal_31388) ) ;
    buf_clk new_AGEMA_reg_buffer_10435 ( .C (clk), .D (new_AGEMA_signal_6752), .Q (new_AGEMA_signal_31391) ) ;
    buf_clk new_AGEMA_reg_buffer_10438 ( .C (clk), .D (new_AGEMA_signal_6753), .Q (new_AGEMA_signal_31394) ) ;
    buf_clk new_AGEMA_reg_buffer_10441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T20), .Q (new_AGEMA_signal_31397) ) ;
    buf_clk new_AGEMA_reg_buffer_10444 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_31400) ) ;
    buf_clk new_AGEMA_reg_buffer_10447 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_31403) ) ;
    buf_clk new_AGEMA_reg_buffer_10450 ( .C (clk), .D (new_AGEMA_signal_7497), .Q (new_AGEMA_signal_31406) ) ;
    buf_clk new_AGEMA_reg_buffer_10453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T1), .Q (new_AGEMA_signal_31409) ) ;
    buf_clk new_AGEMA_reg_buffer_10456 ( .C (clk), .D (new_AGEMA_signal_6241), .Q (new_AGEMA_signal_31412) ) ;
    buf_clk new_AGEMA_reg_buffer_10459 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_31415) ) ;
    buf_clk new_AGEMA_reg_buffer_10462 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_31418) ) ;
    buf_clk new_AGEMA_reg_buffer_10465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T4), .Q (new_AGEMA_signal_31421) ) ;
    buf_clk new_AGEMA_reg_buffer_10468 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_31424) ) ;
    buf_clk new_AGEMA_reg_buffer_10471 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_31427) ) ;
    buf_clk new_AGEMA_reg_buffer_10474 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_31430) ) ;
    buf_clk new_AGEMA_reg_buffer_10477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T2), .Q (new_AGEMA_signal_31433) ) ;
    buf_clk new_AGEMA_reg_buffer_10480 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_31436) ) ;
    buf_clk new_AGEMA_reg_buffer_10483 ( .C (clk), .D (new_AGEMA_signal_6245), .Q (new_AGEMA_signal_31439) ) ;
    buf_clk new_AGEMA_reg_buffer_10486 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_31442) ) ;
    buf_clk new_AGEMA_reg_buffer_10489 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T6), .Q (new_AGEMA_signal_31445) ) ;
    buf_clk new_AGEMA_reg_buffer_10492 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_31448) ) ;
    buf_clk new_AGEMA_reg_buffer_10495 ( .C (clk), .D (new_AGEMA_signal_6758), .Q (new_AGEMA_signal_31451) ) ;
    buf_clk new_AGEMA_reg_buffer_10498 ( .C (clk), .D (new_AGEMA_signal_6759), .Q (new_AGEMA_signal_31454) ) ;
    buf_clk new_AGEMA_reg_buffer_10501 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T8), .Q (new_AGEMA_signal_31457) ) ;
    buf_clk new_AGEMA_reg_buffer_10504 ( .C (clk), .D (new_AGEMA_signal_7522), .Q (new_AGEMA_signal_31460) ) ;
    buf_clk new_AGEMA_reg_buffer_10507 ( .C (clk), .D (new_AGEMA_signal_7523), .Q (new_AGEMA_signal_31463) ) ;
    buf_clk new_AGEMA_reg_buffer_10510 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_31466) ) ;
    buf_clk new_AGEMA_reg_buffer_10513 ( .C (clk), .D (ciphertext_s0[120]), .Q (new_AGEMA_signal_31469) ) ;
    buf_clk new_AGEMA_reg_buffer_10516 ( .C (clk), .D (ciphertext_s1[120]), .Q (new_AGEMA_signal_31472) ) ;
    buf_clk new_AGEMA_reg_buffer_10519 ( .C (clk), .D (ciphertext_s2[120]), .Q (new_AGEMA_signal_31475) ) ;
    buf_clk new_AGEMA_reg_buffer_10522 ( .C (clk), .D (ciphertext_s3[120]), .Q (new_AGEMA_signal_31478) ) ;
    buf_clk new_AGEMA_reg_buffer_10525 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T16), .Q (new_AGEMA_signal_31481) ) ;
    buf_clk new_AGEMA_reg_buffer_10528 ( .C (clk), .D (new_AGEMA_signal_6769), .Q (new_AGEMA_signal_31484) ) ;
    buf_clk new_AGEMA_reg_buffer_10531 ( .C (clk), .D (new_AGEMA_signal_6770), .Q (new_AGEMA_signal_31487) ) ;
    buf_clk new_AGEMA_reg_buffer_10534 ( .C (clk), .D (new_AGEMA_signal_6771), .Q (new_AGEMA_signal_31490) ) ;
    buf_clk new_AGEMA_reg_buffer_10537 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T9), .Q (new_AGEMA_signal_31493) ) ;
    buf_clk new_AGEMA_reg_buffer_10540 ( .C (clk), .D (new_AGEMA_signal_6760), .Q (new_AGEMA_signal_31496) ) ;
    buf_clk new_AGEMA_reg_buffer_10543 ( .C (clk), .D (new_AGEMA_signal_6761), .Q (new_AGEMA_signal_31499) ) ;
    buf_clk new_AGEMA_reg_buffer_10546 ( .C (clk), .D (new_AGEMA_signal_6762), .Q (new_AGEMA_signal_31502) ) ;
    buf_clk new_AGEMA_reg_buffer_10549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T17), .Q (new_AGEMA_signal_31505) ) ;
    buf_clk new_AGEMA_reg_buffer_10552 ( .C (clk), .D (new_AGEMA_signal_7531), .Q (new_AGEMA_signal_31508) ) ;
    buf_clk new_AGEMA_reg_buffer_10555 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_31511) ) ;
    buf_clk new_AGEMA_reg_buffer_10558 ( .C (clk), .D (new_AGEMA_signal_7533), .Q (new_AGEMA_signal_31514) ) ;
    buf_clk new_AGEMA_reg_buffer_10561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T15), .Q (new_AGEMA_signal_31517) ) ;
    buf_clk new_AGEMA_reg_buffer_10564 ( .C (clk), .D (new_AGEMA_signal_6766), .Q (new_AGEMA_signal_31520) ) ;
    buf_clk new_AGEMA_reg_buffer_10567 ( .C (clk), .D (new_AGEMA_signal_6767), .Q (new_AGEMA_signal_31523) ) ;
    buf_clk new_AGEMA_reg_buffer_10570 ( .C (clk), .D (new_AGEMA_signal_6768), .Q (new_AGEMA_signal_31526) ) ;
    buf_clk new_AGEMA_reg_buffer_10573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T27), .Q (new_AGEMA_signal_31529) ) ;
    buf_clk new_AGEMA_reg_buffer_10576 ( .C (clk), .D (new_AGEMA_signal_6778), .Q (new_AGEMA_signal_31532) ) ;
    buf_clk new_AGEMA_reg_buffer_10579 ( .C (clk), .D (new_AGEMA_signal_6779), .Q (new_AGEMA_signal_31535) ) ;
    buf_clk new_AGEMA_reg_buffer_10582 ( .C (clk), .D (new_AGEMA_signal_6780), .Q (new_AGEMA_signal_31538) ) ;
    buf_clk new_AGEMA_reg_buffer_10585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T10), .Q (new_AGEMA_signal_31541) ) ;
    buf_clk new_AGEMA_reg_buffer_10588 ( .C (clk), .D (new_AGEMA_signal_7525), .Q (new_AGEMA_signal_31544) ) ;
    buf_clk new_AGEMA_reg_buffer_10591 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_31547) ) ;
    buf_clk new_AGEMA_reg_buffer_10594 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_31550) ) ;
    buf_clk new_AGEMA_reg_buffer_10597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T13), .Q (new_AGEMA_signal_31553) ) ;
    buf_clk new_AGEMA_reg_buffer_10600 ( .C (clk), .D (new_AGEMA_signal_6763), .Q (new_AGEMA_signal_31556) ) ;
    buf_clk new_AGEMA_reg_buffer_10603 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_31559) ) ;
    buf_clk new_AGEMA_reg_buffer_10606 ( .C (clk), .D (new_AGEMA_signal_6765), .Q (new_AGEMA_signal_31562) ) ;
    buf_clk new_AGEMA_reg_buffer_10609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T23), .Q (new_AGEMA_signal_31565) ) ;
    buf_clk new_AGEMA_reg_buffer_10612 ( .C (clk), .D (new_AGEMA_signal_7537), .Q (new_AGEMA_signal_31568) ) ;
    buf_clk new_AGEMA_reg_buffer_10615 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_31571) ) ;
    buf_clk new_AGEMA_reg_buffer_10618 ( .C (clk), .D (new_AGEMA_signal_7539), .Q (new_AGEMA_signal_31574) ) ;
    buf_clk new_AGEMA_reg_buffer_10621 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T19), .Q (new_AGEMA_signal_31577) ) ;
    buf_clk new_AGEMA_reg_buffer_10624 ( .C (clk), .D (new_AGEMA_signal_6772), .Q (new_AGEMA_signal_31580) ) ;
    buf_clk new_AGEMA_reg_buffer_10627 ( .C (clk), .D (new_AGEMA_signal_6773), .Q (new_AGEMA_signal_31583) ) ;
    buf_clk new_AGEMA_reg_buffer_10630 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_31586) ) ;
    buf_clk new_AGEMA_reg_buffer_10633 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T3), .Q (new_AGEMA_signal_31589) ) ;
    buf_clk new_AGEMA_reg_buffer_10636 ( .C (clk), .D (new_AGEMA_signal_6277), .Q (new_AGEMA_signal_31592) ) ;
    buf_clk new_AGEMA_reg_buffer_10639 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_31595) ) ;
    buf_clk new_AGEMA_reg_buffer_10642 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_31598) ) ;
    buf_clk new_AGEMA_reg_buffer_10645 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T22), .Q (new_AGEMA_signal_31601) ) ;
    buf_clk new_AGEMA_reg_buffer_10648 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_31604) ) ;
    buf_clk new_AGEMA_reg_buffer_10651 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_31607) ) ;
    buf_clk new_AGEMA_reg_buffer_10654 ( .C (clk), .D (new_AGEMA_signal_6777), .Q (new_AGEMA_signal_31610) ) ;
    buf_clk new_AGEMA_reg_buffer_10657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T20), .Q (new_AGEMA_signal_31613) ) ;
    buf_clk new_AGEMA_reg_buffer_10660 ( .C (clk), .D (new_AGEMA_signal_7534), .Q (new_AGEMA_signal_31616) ) ;
    buf_clk new_AGEMA_reg_buffer_10663 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_31619) ) ;
    buf_clk new_AGEMA_reg_buffer_10666 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_31622) ) ;
    buf_clk new_AGEMA_reg_buffer_10669 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T1), .Q (new_AGEMA_signal_31625) ) ;
    buf_clk new_AGEMA_reg_buffer_10672 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_31628) ) ;
    buf_clk new_AGEMA_reg_buffer_10675 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_31631) ) ;
    buf_clk new_AGEMA_reg_buffer_10678 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_31634) ) ;
    buf_clk new_AGEMA_reg_buffer_10681 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T4), .Q (new_AGEMA_signal_31637) ) ;
    buf_clk new_AGEMA_reg_buffer_10684 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_31640) ) ;
    buf_clk new_AGEMA_reg_buffer_10687 ( .C (clk), .D (new_AGEMA_signal_6281), .Q (new_AGEMA_signal_31643) ) ;
    buf_clk new_AGEMA_reg_buffer_10690 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_31646) ) ;
    buf_clk new_AGEMA_reg_buffer_10693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T2), .Q (new_AGEMA_signal_31649) ) ;
    buf_clk new_AGEMA_reg_buffer_10696 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_31652) ) ;
    buf_clk new_AGEMA_reg_buffer_10699 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_31655) ) ;
    buf_clk new_AGEMA_reg_buffer_10702 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_31658) ) ;
    buf_clk new_AGEMA_reg_buffer_10705 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_31661) ) ;
    buf_clk new_AGEMA_reg_buffer_10709 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_31665) ) ;
    buf_clk new_AGEMA_reg_buffer_10713 ( .C (clk), .D (key_s2[0]), .Q (new_AGEMA_signal_31669) ) ;
    buf_clk new_AGEMA_reg_buffer_10717 ( .C (clk), .D (key_s3[0]), .Q (new_AGEMA_signal_31673) ) ;
    buf_clk new_AGEMA_reg_buffer_10721 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_31677) ) ;
    buf_clk new_AGEMA_reg_buffer_10725 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_31681) ) ;
    buf_clk new_AGEMA_reg_buffer_10729 ( .C (clk), .D (key_s2[1]), .Q (new_AGEMA_signal_31685) ) ;
    buf_clk new_AGEMA_reg_buffer_10733 ( .C (clk), .D (key_s3[1]), .Q (new_AGEMA_signal_31689) ) ;
    buf_clk new_AGEMA_reg_buffer_10737 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_31693) ) ;
    buf_clk new_AGEMA_reg_buffer_10741 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_31697) ) ;
    buf_clk new_AGEMA_reg_buffer_10745 ( .C (clk), .D (key_s2[2]), .Q (new_AGEMA_signal_31701) ) ;
    buf_clk new_AGEMA_reg_buffer_10749 ( .C (clk), .D (key_s3[2]), .Q (new_AGEMA_signal_31705) ) ;
    buf_clk new_AGEMA_reg_buffer_10753 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_31709) ) ;
    buf_clk new_AGEMA_reg_buffer_10757 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_31713) ) ;
    buf_clk new_AGEMA_reg_buffer_10761 ( .C (clk), .D (key_s2[3]), .Q (new_AGEMA_signal_31717) ) ;
    buf_clk new_AGEMA_reg_buffer_10765 ( .C (clk), .D (key_s3[3]), .Q (new_AGEMA_signal_31721) ) ;
    buf_clk new_AGEMA_reg_buffer_10769 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_31725) ) ;
    buf_clk new_AGEMA_reg_buffer_10773 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_31729) ) ;
    buf_clk new_AGEMA_reg_buffer_10777 ( .C (clk), .D (key_s2[4]), .Q (new_AGEMA_signal_31733) ) ;
    buf_clk new_AGEMA_reg_buffer_10781 ( .C (clk), .D (key_s3[4]), .Q (new_AGEMA_signal_31737) ) ;
    buf_clk new_AGEMA_reg_buffer_10785 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_31741) ) ;
    buf_clk new_AGEMA_reg_buffer_10789 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_31745) ) ;
    buf_clk new_AGEMA_reg_buffer_10793 ( .C (clk), .D (key_s2[5]), .Q (new_AGEMA_signal_31749) ) ;
    buf_clk new_AGEMA_reg_buffer_10797 ( .C (clk), .D (key_s3[5]), .Q (new_AGEMA_signal_31753) ) ;
    buf_clk new_AGEMA_reg_buffer_10801 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_31757) ) ;
    buf_clk new_AGEMA_reg_buffer_10805 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_31761) ) ;
    buf_clk new_AGEMA_reg_buffer_10809 ( .C (clk), .D (key_s2[6]), .Q (new_AGEMA_signal_31765) ) ;
    buf_clk new_AGEMA_reg_buffer_10813 ( .C (clk), .D (key_s3[6]), .Q (new_AGEMA_signal_31769) ) ;
    buf_clk new_AGEMA_reg_buffer_10817 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_31773) ) ;
    buf_clk new_AGEMA_reg_buffer_10821 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_31777) ) ;
    buf_clk new_AGEMA_reg_buffer_10825 ( .C (clk), .D (key_s2[7]), .Q (new_AGEMA_signal_31781) ) ;
    buf_clk new_AGEMA_reg_buffer_10829 ( .C (clk), .D (key_s3[7]), .Q (new_AGEMA_signal_31785) ) ;
    buf_clk new_AGEMA_reg_buffer_10833 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_31789) ) ;
    buf_clk new_AGEMA_reg_buffer_10837 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_31793) ) ;
    buf_clk new_AGEMA_reg_buffer_10841 ( .C (clk), .D (key_s2[8]), .Q (new_AGEMA_signal_31797) ) ;
    buf_clk new_AGEMA_reg_buffer_10845 ( .C (clk), .D (key_s3[8]), .Q (new_AGEMA_signal_31801) ) ;
    buf_clk new_AGEMA_reg_buffer_10849 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_31805) ) ;
    buf_clk new_AGEMA_reg_buffer_10853 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_31809) ) ;
    buf_clk new_AGEMA_reg_buffer_10857 ( .C (clk), .D (key_s2[9]), .Q (new_AGEMA_signal_31813) ) ;
    buf_clk new_AGEMA_reg_buffer_10861 ( .C (clk), .D (key_s3[9]), .Q (new_AGEMA_signal_31817) ) ;
    buf_clk new_AGEMA_reg_buffer_10865 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_31821) ) ;
    buf_clk new_AGEMA_reg_buffer_10869 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_31825) ) ;
    buf_clk new_AGEMA_reg_buffer_10873 ( .C (clk), .D (key_s2[10]), .Q (new_AGEMA_signal_31829) ) ;
    buf_clk new_AGEMA_reg_buffer_10877 ( .C (clk), .D (key_s3[10]), .Q (new_AGEMA_signal_31833) ) ;
    buf_clk new_AGEMA_reg_buffer_10881 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_31837) ) ;
    buf_clk new_AGEMA_reg_buffer_10885 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_31841) ) ;
    buf_clk new_AGEMA_reg_buffer_10889 ( .C (clk), .D (key_s2[11]), .Q (new_AGEMA_signal_31845) ) ;
    buf_clk new_AGEMA_reg_buffer_10893 ( .C (clk), .D (key_s3[11]), .Q (new_AGEMA_signal_31849) ) ;
    buf_clk new_AGEMA_reg_buffer_10897 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_31853) ) ;
    buf_clk new_AGEMA_reg_buffer_10901 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_31857) ) ;
    buf_clk new_AGEMA_reg_buffer_10905 ( .C (clk), .D (key_s2[12]), .Q (new_AGEMA_signal_31861) ) ;
    buf_clk new_AGEMA_reg_buffer_10909 ( .C (clk), .D (key_s3[12]), .Q (new_AGEMA_signal_31865) ) ;
    buf_clk new_AGEMA_reg_buffer_10913 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_31869) ) ;
    buf_clk new_AGEMA_reg_buffer_10917 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_31873) ) ;
    buf_clk new_AGEMA_reg_buffer_10921 ( .C (clk), .D (key_s2[13]), .Q (new_AGEMA_signal_31877) ) ;
    buf_clk new_AGEMA_reg_buffer_10925 ( .C (clk), .D (key_s3[13]), .Q (new_AGEMA_signal_31881) ) ;
    buf_clk new_AGEMA_reg_buffer_10929 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_31885) ) ;
    buf_clk new_AGEMA_reg_buffer_10933 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_31889) ) ;
    buf_clk new_AGEMA_reg_buffer_10937 ( .C (clk), .D (key_s2[14]), .Q (new_AGEMA_signal_31893) ) ;
    buf_clk new_AGEMA_reg_buffer_10941 ( .C (clk), .D (key_s3[14]), .Q (new_AGEMA_signal_31897) ) ;
    buf_clk new_AGEMA_reg_buffer_10945 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_31901) ) ;
    buf_clk new_AGEMA_reg_buffer_10949 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_31905) ) ;
    buf_clk new_AGEMA_reg_buffer_10953 ( .C (clk), .D (key_s2[15]), .Q (new_AGEMA_signal_31909) ) ;
    buf_clk new_AGEMA_reg_buffer_10957 ( .C (clk), .D (key_s3[15]), .Q (new_AGEMA_signal_31913) ) ;
    buf_clk new_AGEMA_reg_buffer_10961 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_31917) ) ;
    buf_clk new_AGEMA_reg_buffer_10965 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_31921) ) ;
    buf_clk new_AGEMA_reg_buffer_10969 ( .C (clk), .D (key_s2[16]), .Q (new_AGEMA_signal_31925) ) ;
    buf_clk new_AGEMA_reg_buffer_10973 ( .C (clk), .D (key_s3[16]), .Q (new_AGEMA_signal_31929) ) ;
    buf_clk new_AGEMA_reg_buffer_10977 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_31933) ) ;
    buf_clk new_AGEMA_reg_buffer_10981 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_31937) ) ;
    buf_clk new_AGEMA_reg_buffer_10985 ( .C (clk), .D (key_s2[17]), .Q (new_AGEMA_signal_31941) ) ;
    buf_clk new_AGEMA_reg_buffer_10989 ( .C (clk), .D (key_s3[17]), .Q (new_AGEMA_signal_31945) ) ;
    buf_clk new_AGEMA_reg_buffer_10993 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_31949) ) ;
    buf_clk new_AGEMA_reg_buffer_10997 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_31953) ) ;
    buf_clk new_AGEMA_reg_buffer_11001 ( .C (clk), .D (key_s2[18]), .Q (new_AGEMA_signal_31957) ) ;
    buf_clk new_AGEMA_reg_buffer_11005 ( .C (clk), .D (key_s3[18]), .Q (new_AGEMA_signal_31961) ) ;
    buf_clk new_AGEMA_reg_buffer_11009 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_31965) ) ;
    buf_clk new_AGEMA_reg_buffer_11013 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_31969) ) ;
    buf_clk new_AGEMA_reg_buffer_11017 ( .C (clk), .D (key_s2[19]), .Q (new_AGEMA_signal_31973) ) ;
    buf_clk new_AGEMA_reg_buffer_11021 ( .C (clk), .D (key_s3[19]), .Q (new_AGEMA_signal_31977) ) ;
    buf_clk new_AGEMA_reg_buffer_11025 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_31981) ) ;
    buf_clk new_AGEMA_reg_buffer_11029 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_31985) ) ;
    buf_clk new_AGEMA_reg_buffer_11033 ( .C (clk), .D (key_s2[20]), .Q (new_AGEMA_signal_31989) ) ;
    buf_clk new_AGEMA_reg_buffer_11037 ( .C (clk), .D (key_s3[20]), .Q (new_AGEMA_signal_31993) ) ;
    buf_clk new_AGEMA_reg_buffer_11041 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_31997) ) ;
    buf_clk new_AGEMA_reg_buffer_11045 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_32001) ) ;
    buf_clk new_AGEMA_reg_buffer_11049 ( .C (clk), .D (key_s2[21]), .Q (new_AGEMA_signal_32005) ) ;
    buf_clk new_AGEMA_reg_buffer_11053 ( .C (clk), .D (key_s3[21]), .Q (new_AGEMA_signal_32009) ) ;
    buf_clk new_AGEMA_reg_buffer_11057 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_32013) ) ;
    buf_clk new_AGEMA_reg_buffer_11061 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_32017) ) ;
    buf_clk new_AGEMA_reg_buffer_11065 ( .C (clk), .D (key_s2[22]), .Q (new_AGEMA_signal_32021) ) ;
    buf_clk new_AGEMA_reg_buffer_11069 ( .C (clk), .D (key_s3[22]), .Q (new_AGEMA_signal_32025) ) ;
    buf_clk new_AGEMA_reg_buffer_11073 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_32029) ) ;
    buf_clk new_AGEMA_reg_buffer_11077 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_32033) ) ;
    buf_clk new_AGEMA_reg_buffer_11081 ( .C (clk), .D (key_s2[23]), .Q (new_AGEMA_signal_32037) ) ;
    buf_clk new_AGEMA_reg_buffer_11085 ( .C (clk), .D (key_s3[23]), .Q (new_AGEMA_signal_32041) ) ;
    buf_clk new_AGEMA_reg_buffer_11089 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_32045) ) ;
    buf_clk new_AGEMA_reg_buffer_11093 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_32049) ) ;
    buf_clk new_AGEMA_reg_buffer_11097 ( .C (clk), .D (key_s2[24]), .Q (new_AGEMA_signal_32053) ) ;
    buf_clk new_AGEMA_reg_buffer_11101 ( .C (clk), .D (key_s3[24]), .Q (new_AGEMA_signal_32057) ) ;
    buf_clk new_AGEMA_reg_buffer_11105 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_32061) ) ;
    buf_clk new_AGEMA_reg_buffer_11109 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_32065) ) ;
    buf_clk new_AGEMA_reg_buffer_11113 ( .C (clk), .D (key_s2[25]), .Q (new_AGEMA_signal_32069) ) ;
    buf_clk new_AGEMA_reg_buffer_11117 ( .C (clk), .D (key_s3[25]), .Q (new_AGEMA_signal_32073) ) ;
    buf_clk new_AGEMA_reg_buffer_11121 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_32077) ) ;
    buf_clk new_AGEMA_reg_buffer_11125 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_32081) ) ;
    buf_clk new_AGEMA_reg_buffer_11129 ( .C (clk), .D (key_s2[26]), .Q (new_AGEMA_signal_32085) ) ;
    buf_clk new_AGEMA_reg_buffer_11133 ( .C (clk), .D (key_s3[26]), .Q (new_AGEMA_signal_32089) ) ;
    buf_clk new_AGEMA_reg_buffer_11137 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_32093) ) ;
    buf_clk new_AGEMA_reg_buffer_11141 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_32097) ) ;
    buf_clk new_AGEMA_reg_buffer_11145 ( .C (clk), .D (key_s2[27]), .Q (new_AGEMA_signal_32101) ) ;
    buf_clk new_AGEMA_reg_buffer_11149 ( .C (clk), .D (key_s3[27]), .Q (new_AGEMA_signal_32105) ) ;
    buf_clk new_AGEMA_reg_buffer_11153 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_32109) ) ;
    buf_clk new_AGEMA_reg_buffer_11157 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_32113) ) ;
    buf_clk new_AGEMA_reg_buffer_11161 ( .C (clk), .D (key_s2[28]), .Q (new_AGEMA_signal_32117) ) ;
    buf_clk new_AGEMA_reg_buffer_11165 ( .C (clk), .D (key_s3[28]), .Q (new_AGEMA_signal_32121) ) ;
    buf_clk new_AGEMA_reg_buffer_11169 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_32125) ) ;
    buf_clk new_AGEMA_reg_buffer_11173 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_32129) ) ;
    buf_clk new_AGEMA_reg_buffer_11177 ( .C (clk), .D (key_s2[29]), .Q (new_AGEMA_signal_32133) ) ;
    buf_clk new_AGEMA_reg_buffer_11181 ( .C (clk), .D (key_s3[29]), .Q (new_AGEMA_signal_32137) ) ;
    buf_clk new_AGEMA_reg_buffer_11185 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_32141) ) ;
    buf_clk new_AGEMA_reg_buffer_11189 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_32145) ) ;
    buf_clk new_AGEMA_reg_buffer_11193 ( .C (clk), .D (key_s2[30]), .Q (new_AGEMA_signal_32149) ) ;
    buf_clk new_AGEMA_reg_buffer_11197 ( .C (clk), .D (key_s3[30]), .Q (new_AGEMA_signal_32153) ) ;
    buf_clk new_AGEMA_reg_buffer_11201 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_32157) ) ;
    buf_clk new_AGEMA_reg_buffer_11205 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_32161) ) ;
    buf_clk new_AGEMA_reg_buffer_11209 ( .C (clk), .D (key_s2[31]), .Q (new_AGEMA_signal_32165) ) ;
    buf_clk new_AGEMA_reg_buffer_11213 ( .C (clk), .D (key_s3[31]), .Q (new_AGEMA_signal_32169) ) ;
    buf_clk new_AGEMA_reg_buffer_11217 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_32173) ) ;
    buf_clk new_AGEMA_reg_buffer_11221 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_32177) ) ;
    buf_clk new_AGEMA_reg_buffer_11225 ( .C (clk), .D (key_s2[32]), .Q (new_AGEMA_signal_32181) ) ;
    buf_clk new_AGEMA_reg_buffer_11229 ( .C (clk), .D (key_s3[32]), .Q (new_AGEMA_signal_32185) ) ;
    buf_clk new_AGEMA_reg_buffer_11233 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_32189) ) ;
    buf_clk new_AGEMA_reg_buffer_11237 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_32193) ) ;
    buf_clk new_AGEMA_reg_buffer_11241 ( .C (clk), .D (key_s2[33]), .Q (new_AGEMA_signal_32197) ) ;
    buf_clk new_AGEMA_reg_buffer_11245 ( .C (clk), .D (key_s3[33]), .Q (new_AGEMA_signal_32201) ) ;
    buf_clk new_AGEMA_reg_buffer_11249 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_32205) ) ;
    buf_clk new_AGEMA_reg_buffer_11253 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_32209) ) ;
    buf_clk new_AGEMA_reg_buffer_11257 ( .C (clk), .D (key_s2[34]), .Q (new_AGEMA_signal_32213) ) ;
    buf_clk new_AGEMA_reg_buffer_11261 ( .C (clk), .D (key_s3[34]), .Q (new_AGEMA_signal_32217) ) ;
    buf_clk new_AGEMA_reg_buffer_11265 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_32221) ) ;
    buf_clk new_AGEMA_reg_buffer_11269 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_32225) ) ;
    buf_clk new_AGEMA_reg_buffer_11273 ( .C (clk), .D (key_s2[35]), .Q (new_AGEMA_signal_32229) ) ;
    buf_clk new_AGEMA_reg_buffer_11277 ( .C (clk), .D (key_s3[35]), .Q (new_AGEMA_signal_32233) ) ;
    buf_clk new_AGEMA_reg_buffer_11281 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_32237) ) ;
    buf_clk new_AGEMA_reg_buffer_11285 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_32241) ) ;
    buf_clk new_AGEMA_reg_buffer_11289 ( .C (clk), .D (key_s2[36]), .Q (new_AGEMA_signal_32245) ) ;
    buf_clk new_AGEMA_reg_buffer_11293 ( .C (clk), .D (key_s3[36]), .Q (new_AGEMA_signal_32249) ) ;
    buf_clk new_AGEMA_reg_buffer_11297 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_32253) ) ;
    buf_clk new_AGEMA_reg_buffer_11301 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_32257) ) ;
    buf_clk new_AGEMA_reg_buffer_11305 ( .C (clk), .D (key_s2[37]), .Q (new_AGEMA_signal_32261) ) ;
    buf_clk new_AGEMA_reg_buffer_11309 ( .C (clk), .D (key_s3[37]), .Q (new_AGEMA_signal_32265) ) ;
    buf_clk new_AGEMA_reg_buffer_11313 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_32269) ) ;
    buf_clk new_AGEMA_reg_buffer_11317 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_32273) ) ;
    buf_clk new_AGEMA_reg_buffer_11321 ( .C (clk), .D (key_s2[38]), .Q (new_AGEMA_signal_32277) ) ;
    buf_clk new_AGEMA_reg_buffer_11325 ( .C (clk), .D (key_s3[38]), .Q (new_AGEMA_signal_32281) ) ;
    buf_clk new_AGEMA_reg_buffer_11329 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_32285) ) ;
    buf_clk new_AGEMA_reg_buffer_11333 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_32289) ) ;
    buf_clk new_AGEMA_reg_buffer_11337 ( .C (clk), .D (key_s2[39]), .Q (new_AGEMA_signal_32293) ) ;
    buf_clk new_AGEMA_reg_buffer_11341 ( .C (clk), .D (key_s3[39]), .Q (new_AGEMA_signal_32297) ) ;
    buf_clk new_AGEMA_reg_buffer_11345 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_32301) ) ;
    buf_clk new_AGEMA_reg_buffer_11349 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_32305) ) ;
    buf_clk new_AGEMA_reg_buffer_11353 ( .C (clk), .D (key_s2[40]), .Q (new_AGEMA_signal_32309) ) ;
    buf_clk new_AGEMA_reg_buffer_11357 ( .C (clk), .D (key_s3[40]), .Q (new_AGEMA_signal_32313) ) ;
    buf_clk new_AGEMA_reg_buffer_11361 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_32317) ) ;
    buf_clk new_AGEMA_reg_buffer_11365 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_32321) ) ;
    buf_clk new_AGEMA_reg_buffer_11369 ( .C (clk), .D (key_s2[41]), .Q (new_AGEMA_signal_32325) ) ;
    buf_clk new_AGEMA_reg_buffer_11373 ( .C (clk), .D (key_s3[41]), .Q (new_AGEMA_signal_32329) ) ;
    buf_clk new_AGEMA_reg_buffer_11377 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_32333) ) ;
    buf_clk new_AGEMA_reg_buffer_11381 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_32337) ) ;
    buf_clk new_AGEMA_reg_buffer_11385 ( .C (clk), .D (key_s2[42]), .Q (new_AGEMA_signal_32341) ) ;
    buf_clk new_AGEMA_reg_buffer_11389 ( .C (clk), .D (key_s3[42]), .Q (new_AGEMA_signal_32345) ) ;
    buf_clk new_AGEMA_reg_buffer_11393 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_32349) ) ;
    buf_clk new_AGEMA_reg_buffer_11397 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_32353) ) ;
    buf_clk new_AGEMA_reg_buffer_11401 ( .C (clk), .D (key_s2[43]), .Q (new_AGEMA_signal_32357) ) ;
    buf_clk new_AGEMA_reg_buffer_11405 ( .C (clk), .D (key_s3[43]), .Q (new_AGEMA_signal_32361) ) ;
    buf_clk new_AGEMA_reg_buffer_11409 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_32365) ) ;
    buf_clk new_AGEMA_reg_buffer_11413 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_32369) ) ;
    buf_clk new_AGEMA_reg_buffer_11417 ( .C (clk), .D (key_s2[44]), .Q (new_AGEMA_signal_32373) ) ;
    buf_clk new_AGEMA_reg_buffer_11421 ( .C (clk), .D (key_s3[44]), .Q (new_AGEMA_signal_32377) ) ;
    buf_clk new_AGEMA_reg_buffer_11425 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_32381) ) ;
    buf_clk new_AGEMA_reg_buffer_11429 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_32385) ) ;
    buf_clk new_AGEMA_reg_buffer_11433 ( .C (clk), .D (key_s2[45]), .Q (new_AGEMA_signal_32389) ) ;
    buf_clk new_AGEMA_reg_buffer_11437 ( .C (clk), .D (key_s3[45]), .Q (new_AGEMA_signal_32393) ) ;
    buf_clk new_AGEMA_reg_buffer_11441 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_32397) ) ;
    buf_clk new_AGEMA_reg_buffer_11445 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_32401) ) ;
    buf_clk new_AGEMA_reg_buffer_11449 ( .C (clk), .D (key_s2[46]), .Q (new_AGEMA_signal_32405) ) ;
    buf_clk new_AGEMA_reg_buffer_11453 ( .C (clk), .D (key_s3[46]), .Q (new_AGEMA_signal_32409) ) ;
    buf_clk new_AGEMA_reg_buffer_11457 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_32413) ) ;
    buf_clk new_AGEMA_reg_buffer_11461 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_32417) ) ;
    buf_clk new_AGEMA_reg_buffer_11465 ( .C (clk), .D (key_s2[47]), .Q (new_AGEMA_signal_32421) ) ;
    buf_clk new_AGEMA_reg_buffer_11469 ( .C (clk), .D (key_s3[47]), .Q (new_AGEMA_signal_32425) ) ;
    buf_clk new_AGEMA_reg_buffer_11473 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_32429) ) ;
    buf_clk new_AGEMA_reg_buffer_11477 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_32433) ) ;
    buf_clk new_AGEMA_reg_buffer_11481 ( .C (clk), .D (key_s2[48]), .Q (new_AGEMA_signal_32437) ) ;
    buf_clk new_AGEMA_reg_buffer_11485 ( .C (clk), .D (key_s3[48]), .Q (new_AGEMA_signal_32441) ) ;
    buf_clk new_AGEMA_reg_buffer_11489 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_32445) ) ;
    buf_clk new_AGEMA_reg_buffer_11493 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_32449) ) ;
    buf_clk new_AGEMA_reg_buffer_11497 ( .C (clk), .D (key_s2[49]), .Q (new_AGEMA_signal_32453) ) ;
    buf_clk new_AGEMA_reg_buffer_11501 ( .C (clk), .D (key_s3[49]), .Q (new_AGEMA_signal_32457) ) ;
    buf_clk new_AGEMA_reg_buffer_11505 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_32461) ) ;
    buf_clk new_AGEMA_reg_buffer_11509 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_32465) ) ;
    buf_clk new_AGEMA_reg_buffer_11513 ( .C (clk), .D (key_s2[50]), .Q (new_AGEMA_signal_32469) ) ;
    buf_clk new_AGEMA_reg_buffer_11517 ( .C (clk), .D (key_s3[50]), .Q (new_AGEMA_signal_32473) ) ;
    buf_clk new_AGEMA_reg_buffer_11521 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_32477) ) ;
    buf_clk new_AGEMA_reg_buffer_11525 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_32481) ) ;
    buf_clk new_AGEMA_reg_buffer_11529 ( .C (clk), .D (key_s2[51]), .Q (new_AGEMA_signal_32485) ) ;
    buf_clk new_AGEMA_reg_buffer_11533 ( .C (clk), .D (key_s3[51]), .Q (new_AGEMA_signal_32489) ) ;
    buf_clk new_AGEMA_reg_buffer_11537 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_32493) ) ;
    buf_clk new_AGEMA_reg_buffer_11541 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_32497) ) ;
    buf_clk new_AGEMA_reg_buffer_11545 ( .C (clk), .D (key_s2[52]), .Q (new_AGEMA_signal_32501) ) ;
    buf_clk new_AGEMA_reg_buffer_11549 ( .C (clk), .D (key_s3[52]), .Q (new_AGEMA_signal_32505) ) ;
    buf_clk new_AGEMA_reg_buffer_11553 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_32509) ) ;
    buf_clk new_AGEMA_reg_buffer_11557 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_32513) ) ;
    buf_clk new_AGEMA_reg_buffer_11561 ( .C (clk), .D (key_s2[53]), .Q (new_AGEMA_signal_32517) ) ;
    buf_clk new_AGEMA_reg_buffer_11565 ( .C (clk), .D (key_s3[53]), .Q (new_AGEMA_signal_32521) ) ;
    buf_clk new_AGEMA_reg_buffer_11569 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_32525) ) ;
    buf_clk new_AGEMA_reg_buffer_11573 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_32529) ) ;
    buf_clk new_AGEMA_reg_buffer_11577 ( .C (clk), .D (key_s2[54]), .Q (new_AGEMA_signal_32533) ) ;
    buf_clk new_AGEMA_reg_buffer_11581 ( .C (clk), .D (key_s3[54]), .Q (new_AGEMA_signal_32537) ) ;
    buf_clk new_AGEMA_reg_buffer_11585 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_32541) ) ;
    buf_clk new_AGEMA_reg_buffer_11589 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_32545) ) ;
    buf_clk new_AGEMA_reg_buffer_11593 ( .C (clk), .D (key_s2[55]), .Q (new_AGEMA_signal_32549) ) ;
    buf_clk new_AGEMA_reg_buffer_11597 ( .C (clk), .D (key_s3[55]), .Q (new_AGEMA_signal_32553) ) ;
    buf_clk new_AGEMA_reg_buffer_11601 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_32557) ) ;
    buf_clk new_AGEMA_reg_buffer_11605 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_32561) ) ;
    buf_clk new_AGEMA_reg_buffer_11609 ( .C (clk), .D (key_s2[56]), .Q (new_AGEMA_signal_32565) ) ;
    buf_clk new_AGEMA_reg_buffer_11613 ( .C (clk), .D (key_s3[56]), .Q (new_AGEMA_signal_32569) ) ;
    buf_clk new_AGEMA_reg_buffer_11617 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_32573) ) ;
    buf_clk new_AGEMA_reg_buffer_11621 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_32577) ) ;
    buf_clk new_AGEMA_reg_buffer_11625 ( .C (clk), .D (key_s2[57]), .Q (new_AGEMA_signal_32581) ) ;
    buf_clk new_AGEMA_reg_buffer_11629 ( .C (clk), .D (key_s3[57]), .Q (new_AGEMA_signal_32585) ) ;
    buf_clk new_AGEMA_reg_buffer_11633 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_32589) ) ;
    buf_clk new_AGEMA_reg_buffer_11637 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_32593) ) ;
    buf_clk new_AGEMA_reg_buffer_11641 ( .C (clk), .D (key_s2[58]), .Q (new_AGEMA_signal_32597) ) ;
    buf_clk new_AGEMA_reg_buffer_11645 ( .C (clk), .D (key_s3[58]), .Q (new_AGEMA_signal_32601) ) ;
    buf_clk new_AGEMA_reg_buffer_11649 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_32605) ) ;
    buf_clk new_AGEMA_reg_buffer_11653 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_32609) ) ;
    buf_clk new_AGEMA_reg_buffer_11657 ( .C (clk), .D (key_s2[59]), .Q (new_AGEMA_signal_32613) ) ;
    buf_clk new_AGEMA_reg_buffer_11661 ( .C (clk), .D (key_s3[59]), .Q (new_AGEMA_signal_32617) ) ;
    buf_clk new_AGEMA_reg_buffer_11665 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_32621) ) ;
    buf_clk new_AGEMA_reg_buffer_11669 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_32625) ) ;
    buf_clk new_AGEMA_reg_buffer_11673 ( .C (clk), .D (key_s2[60]), .Q (new_AGEMA_signal_32629) ) ;
    buf_clk new_AGEMA_reg_buffer_11677 ( .C (clk), .D (key_s3[60]), .Q (new_AGEMA_signal_32633) ) ;
    buf_clk new_AGEMA_reg_buffer_11681 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_32637) ) ;
    buf_clk new_AGEMA_reg_buffer_11685 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_32641) ) ;
    buf_clk new_AGEMA_reg_buffer_11689 ( .C (clk), .D (key_s2[61]), .Q (new_AGEMA_signal_32645) ) ;
    buf_clk new_AGEMA_reg_buffer_11693 ( .C (clk), .D (key_s3[61]), .Q (new_AGEMA_signal_32649) ) ;
    buf_clk new_AGEMA_reg_buffer_11697 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_32653) ) ;
    buf_clk new_AGEMA_reg_buffer_11701 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_32657) ) ;
    buf_clk new_AGEMA_reg_buffer_11705 ( .C (clk), .D (key_s2[62]), .Q (new_AGEMA_signal_32661) ) ;
    buf_clk new_AGEMA_reg_buffer_11709 ( .C (clk), .D (key_s3[62]), .Q (new_AGEMA_signal_32665) ) ;
    buf_clk new_AGEMA_reg_buffer_11713 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_32669) ) ;
    buf_clk new_AGEMA_reg_buffer_11717 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_32673) ) ;
    buf_clk new_AGEMA_reg_buffer_11721 ( .C (clk), .D (key_s2[63]), .Q (new_AGEMA_signal_32677) ) ;
    buf_clk new_AGEMA_reg_buffer_11725 ( .C (clk), .D (key_s3[63]), .Q (new_AGEMA_signal_32681) ) ;
    buf_clk new_AGEMA_reg_buffer_11729 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_32685) ) ;
    buf_clk new_AGEMA_reg_buffer_11733 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_32689) ) ;
    buf_clk new_AGEMA_reg_buffer_11737 ( .C (clk), .D (key_s2[64]), .Q (new_AGEMA_signal_32693) ) ;
    buf_clk new_AGEMA_reg_buffer_11741 ( .C (clk), .D (key_s3[64]), .Q (new_AGEMA_signal_32697) ) ;
    buf_clk new_AGEMA_reg_buffer_11745 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_32701) ) ;
    buf_clk new_AGEMA_reg_buffer_11749 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_32705) ) ;
    buf_clk new_AGEMA_reg_buffer_11753 ( .C (clk), .D (key_s2[65]), .Q (new_AGEMA_signal_32709) ) ;
    buf_clk new_AGEMA_reg_buffer_11757 ( .C (clk), .D (key_s3[65]), .Q (new_AGEMA_signal_32713) ) ;
    buf_clk new_AGEMA_reg_buffer_11761 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_32717) ) ;
    buf_clk new_AGEMA_reg_buffer_11765 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_32721) ) ;
    buf_clk new_AGEMA_reg_buffer_11769 ( .C (clk), .D (key_s2[66]), .Q (new_AGEMA_signal_32725) ) ;
    buf_clk new_AGEMA_reg_buffer_11773 ( .C (clk), .D (key_s3[66]), .Q (new_AGEMA_signal_32729) ) ;
    buf_clk new_AGEMA_reg_buffer_11777 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_32733) ) ;
    buf_clk new_AGEMA_reg_buffer_11781 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_32737) ) ;
    buf_clk new_AGEMA_reg_buffer_11785 ( .C (clk), .D (key_s2[67]), .Q (new_AGEMA_signal_32741) ) ;
    buf_clk new_AGEMA_reg_buffer_11789 ( .C (clk), .D (key_s3[67]), .Q (new_AGEMA_signal_32745) ) ;
    buf_clk new_AGEMA_reg_buffer_11793 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_32749) ) ;
    buf_clk new_AGEMA_reg_buffer_11797 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_32753) ) ;
    buf_clk new_AGEMA_reg_buffer_11801 ( .C (clk), .D (key_s2[68]), .Q (new_AGEMA_signal_32757) ) ;
    buf_clk new_AGEMA_reg_buffer_11805 ( .C (clk), .D (key_s3[68]), .Q (new_AGEMA_signal_32761) ) ;
    buf_clk new_AGEMA_reg_buffer_11809 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_32765) ) ;
    buf_clk new_AGEMA_reg_buffer_11813 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_32769) ) ;
    buf_clk new_AGEMA_reg_buffer_11817 ( .C (clk), .D (key_s2[69]), .Q (new_AGEMA_signal_32773) ) ;
    buf_clk new_AGEMA_reg_buffer_11821 ( .C (clk), .D (key_s3[69]), .Q (new_AGEMA_signal_32777) ) ;
    buf_clk new_AGEMA_reg_buffer_11825 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_32781) ) ;
    buf_clk new_AGEMA_reg_buffer_11829 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_32785) ) ;
    buf_clk new_AGEMA_reg_buffer_11833 ( .C (clk), .D (key_s2[70]), .Q (new_AGEMA_signal_32789) ) ;
    buf_clk new_AGEMA_reg_buffer_11837 ( .C (clk), .D (key_s3[70]), .Q (new_AGEMA_signal_32793) ) ;
    buf_clk new_AGEMA_reg_buffer_11841 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_32797) ) ;
    buf_clk new_AGEMA_reg_buffer_11845 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_32801) ) ;
    buf_clk new_AGEMA_reg_buffer_11849 ( .C (clk), .D (key_s2[71]), .Q (new_AGEMA_signal_32805) ) ;
    buf_clk new_AGEMA_reg_buffer_11853 ( .C (clk), .D (key_s3[71]), .Q (new_AGEMA_signal_32809) ) ;
    buf_clk new_AGEMA_reg_buffer_11857 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_32813) ) ;
    buf_clk new_AGEMA_reg_buffer_11861 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_32817) ) ;
    buf_clk new_AGEMA_reg_buffer_11865 ( .C (clk), .D (key_s2[72]), .Q (new_AGEMA_signal_32821) ) ;
    buf_clk new_AGEMA_reg_buffer_11869 ( .C (clk), .D (key_s3[72]), .Q (new_AGEMA_signal_32825) ) ;
    buf_clk new_AGEMA_reg_buffer_11873 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_32829) ) ;
    buf_clk new_AGEMA_reg_buffer_11877 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_32833) ) ;
    buf_clk new_AGEMA_reg_buffer_11881 ( .C (clk), .D (key_s2[73]), .Q (new_AGEMA_signal_32837) ) ;
    buf_clk new_AGEMA_reg_buffer_11885 ( .C (clk), .D (key_s3[73]), .Q (new_AGEMA_signal_32841) ) ;
    buf_clk new_AGEMA_reg_buffer_11889 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_32845) ) ;
    buf_clk new_AGEMA_reg_buffer_11893 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_32849) ) ;
    buf_clk new_AGEMA_reg_buffer_11897 ( .C (clk), .D (key_s2[74]), .Q (new_AGEMA_signal_32853) ) ;
    buf_clk new_AGEMA_reg_buffer_11901 ( .C (clk), .D (key_s3[74]), .Q (new_AGEMA_signal_32857) ) ;
    buf_clk new_AGEMA_reg_buffer_11905 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_32861) ) ;
    buf_clk new_AGEMA_reg_buffer_11909 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_32865) ) ;
    buf_clk new_AGEMA_reg_buffer_11913 ( .C (clk), .D (key_s2[75]), .Q (new_AGEMA_signal_32869) ) ;
    buf_clk new_AGEMA_reg_buffer_11917 ( .C (clk), .D (key_s3[75]), .Q (new_AGEMA_signal_32873) ) ;
    buf_clk new_AGEMA_reg_buffer_11921 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_32877) ) ;
    buf_clk new_AGEMA_reg_buffer_11925 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_32881) ) ;
    buf_clk new_AGEMA_reg_buffer_11929 ( .C (clk), .D (key_s2[76]), .Q (new_AGEMA_signal_32885) ) ;
    buf_clk new_AGEMA_reg_buffer_11933 ( .C (clk), .D (key_s3[76]), .Q (new_AGEMA_signal_32889) ) ;
    buf_clk new_AGEMA_reg_buffer_11937 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_32893) ) ;
    buf_clk new_AGEMA_reg_buffer_11941 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_32897) ) ;
    buf_clk new_AGEMA_reg_buffer_11945 ( .C (clk), .D (key_s2[77]), .Q (new_AGEMA_signal_32901) ) ;
    buf_clk new_AGEMA_reg_buffer_11949 ( .C (clk), .D (key_s3[77]), .Q (new_AGEMA_signal_32905) ) ;
    buf_clk new_AGEMA_reg_buffer_11953 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_32909) ) ;
    buf_clk new_AGEMA_reg_buffer_11957 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_32913) ) ;
    buf_clk new_AGEMA_reg_buffer_11961 ( .C (clk), .D (key_s2[78]), .Q (new_AGEMA_signal_32917) ) ;
    buf_clk new_AGEMA_reg_buffer_11965 ( .C (clk), .D (key_s3[78]), .Q (new_AGEMA_signal_32921) ) ;
    buf_clk new_AGEMA_reg_buffer_11969 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_32925) ) ;
    buf_clk new_AGEMA_reg_buffer_11973 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_32929) ) ;
    buf_clk new_AGEMA_reg_buffer_11977 ( .C (clk), .D (key_s2[79]), .Q (new_AGEMA_signal_32933) ) ;
    buf_clk new_AGEMA_reg_buffer_11981 ( .C (clk), .D (key_s3[79]), .Q (new_AGEMA_signal_32937) ) ;
    buf_clk new_AGEMA_reg_buffer_11985 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_32941) ) ;
    buf_clk new_AGEMA_reg_buffer_11989 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_32945) ) ;
    buf_clk new_AGEMA_reg_buffer_11993 ( .C (clk), .D (key_s2[80]), .Q (new_AGEMA_signal_32949) ) ;
    buf_clk new_AGEMA_reg_buffer_11997 ( .C (clk), .D (key_s3[80]), .Q (new_AGEMA_signal_32953) ) ;
    buf_clk new_AGEMA_reg_buffer_12001 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_32957) ) ;
    buf_clk new_AGEMA_reg_buffer_12005 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_32961) ) ;
    buf_clk new_AGEMA_reg_buffer_12009 ( .C (clk), .D (key_s2[81]), .Q (new_AGEMA_signal_32965) ) ;
    buf_clk new_AGEMA_reg_buffer_12013 ( .C (clk), .D (key_s3[81]), .Q (new_AGEMA_signal_32969) ) ;
    buf_clk new_AGEMA_reg_buffer_12017 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_32973) ) ;
    buf_clk new_AGEMA_reg_buffer_12021 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_32977) ) ;
    buf_clk new_AGEMA_reg_buffer_12025 ( .C (clk), .D (key_s2[82]), .Q (new_AGEMA_signal_32981) ) ;
    buf_clk new_AGEMA_reg_buffer_12029 ( .C (clk), .D (key_s3[82]), .Q (new_AGEMA_signal_32985) ) ;
    buf_clk new_AGEMA_reg_buffer_12033 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_32989) ) ;
    buf_clk new_AGEMA_reg_buffer_12037 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_32993) ) ;
    buf_clk new_AGEMA_reg_buffer_12041 ( .C (clk), .D (key_s2[83]), .Q (new_AGEMA_signal_32997) ) ;
    buf_clk new_AGEMA_reg_buffer_12045 ( .C (clk), .D (key_s3[83]), .Q (new_AGEMA_signal_33001) ) ;
    buf_clk new_AGEMA_reg_buffer_12049 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_33005) ) ;
    buf_clk new_AGEMA_reg_buffer_12053 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_33009) ) ;
    buf_clk new_AGEMA_reg_buffer_12057 ( .C (clk), .D (key_s2[84]), .Q (new_AGEMA_signal_33013) ) ;
    buf_clk new_AGEMA_reg_buffer_12061 ( .C (clk), .D (key_s3[84]), .Q (new_AGEMA_signal_33017) ) ;
    buf_clk new_AGEMA_reg_buffer_12065 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_33021) ) ;
    buf_clk new_AGEMA_reg_buffer_12069 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_33025) ) ;
    buf_clk new_AGEMA_reg_buffer_12073 ( .C (clk), .D (key_s2[85]), .Q (new_AGEMA_signal_33029) ) ;
    buf_clk new_AGEMA_reg_buffer_12077 ( .C (clk), .D (key_s3[85]), .Q (new_AGEMA_signal_33033) ) ;
    buf_clk new_AGEMA_reg_buffer_12081 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_33037) ) ;
    buf_clk new_AGEMA_reg_buffer_12085 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_33041) ) ;
    buf_clk new_AGEMA_reg_buffer_12089 ( .C (clk), .D (key_s2[86]), .Q (new_AGEMA_signal_33045) ) ;
    buf_clk new_AGEMA_reg_buffer_12093 ( .C (clk), .D (key_s3[86]), .Q (new_AGEMA_signal_33049) ) ;
    buf_clk new_AGEMA_reg_buffer_12097 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_33053) ) ;
    buf_clk new_AGEMA_reg_buffer_12101 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_33057) ) ;
    buf_clk new_AGEMA_reg_buffer_12105 ( .C (clk), .D (key_s2[87]), .Q (new_AGEMA_signal_33061) ) ;
    buf_clk new_AGEMA_reg_buffer_12109 ( .C (clk), .D (key_s3[87]), .Q (new_AGEMA_signal_33065) ) ;
    buf_clk new_AGEMA_reg_buffer_12113 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_33069) ) ;
    buf_clk new_AGEMA_reg_buffer_12117 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_33073) ) ;
    buf_clk new_AGEMA_reg_buffer_12121 ( .C (clk), .D (key_s2[88]), .Q (new_AGEMA_signal_33077) ) ;
    buf_clk new_AGEMA_reg_buffer_12125 ( .C (clk), .D (key_s3[88]), .Q (new_AGEMA_signal_33081) ) ;
    buf_clk new_AGEMA_reg_buffer_12129 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_33085) ) ;
    buf_clk new_AGEMA_reg_buffer_12133 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_33089) ) ;
    buf_clk new_AGEMA_reg_buffer_12137 ( .C (clk), .D (key_s2[89]), .Q (new_AGEMA_signal_33093) ) ;
    buf_clk new_AGEMA_reg_buffer_12141 ( .C (clk), .D (key_s3[89]), .Q (new_AGEMA_signal_33097) ) ;
    buf_clk new_AGEMA_reg_buffer_12145 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_33101) ) ;
    buf_clk new_AGEMA_reg_buffer_12149 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_33105) ) ;
    buf_clk new_AGEMA_reg_buffer_12153 ( .C (clk), .D (key_s2[90]), .Q (new_AGEMA_signal_33109) ) ;
    buf_clk new_AGEMA_reg_buffer_12157 ( .C (clk), .D (key_s3[90]), .Q (new_AGEMA_signal_33113) ) ;
    buf_clk new_AGEMA_reg_buffer_12161 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_33117) ) ;
    buf_clk new_AGEMA_reg_buffer_12165 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_33121) ) ;
    buf_clk new_AGEMA_reg_buffer_12169 ( .C (clk), .D (key_s2[91]), .Q (new_AGEMA_signal_33125) ) ;
    buf_clk new_AGEMA_reg_buffer_12173 ( .C (clk), .D (key_s3[91]), .Q (new_AGEMA_signal_33129) ) ;
    buf_clk new_AGEMA_reg_buffer_12177 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_33133) ) ;
    buf_clk new_AGEMA_reg_buffer_12181 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_33137) ) ;
    buf_clk new_AGEMA_reg_buffer_12185 ( .C (clk), .D (key_s2[92]), .Q (new_AGEMA_signal_33141) ) ;
    buf_clk new_AGEMA_reg_buffer_12189 ( .C (clk), .D (key_s3[92]), .Q (new_AGEMA_signal_33145) ) ;
    buf_clk new_AGEMA_reg_buffer_12193 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_33149) ) ;
    buf_clk new_AGEMA_reg_buffer_12197 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_33153) ) ;
    buf_clk new_AGEMA_reg_buffer_12201 ( .C (clk), .D (key_s2[93]), .Q (new_AGEMA_signal_33157) ) ;
    buf_clk new_AGEMA_reg_buffer_12205 ( .C (clk), .D (key_s3[93]), .Q (new_AGEMA_signal_33161) ) ;
    buf_clk new_AGEMA_reg_buffer_12209 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_33165) ) ;
    buf_clk new_AGEMA_reg_buffer_12213 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_33169) ) ;
    buf_clk new_AGEMA_reg_buffer_12217 ( .C (clk), .D (key_s2[94]), .Q (new_AGEMA_signal_33173) ) ;
    buf_clk new_AGEMA_reg_buffer_12221 ( .C (clk), .D (key_s3[94]), .Q (new_AGEMA_signal_33177) ) ;
    buf_clk new_AGEMA_reg_buffer_12225 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_33181) ) ;
    buf_clk new_AGEMA_reg_buffer_12229 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_33185) ) ;
    buf_clk new_AGEMA_reg_buffer_12233 ( .C (clk), .D (key_s2[95]), .Q (new_AGEMA_signal_33189) ) ;
    buf_clk new_AGEMA_reg_buffer_12237 ( .C (clk), .D (key_s3[95]), .Q (new_AGEMA_signal_33193) ) ;
    buf_clk new_AGEMA_reg_buffer_12241 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_33197) ) ;
    buf_clk new_AGEMA_reg_buffer_12245 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_33201) ) ;
    buf_clk new_AGEMA_reg_buffer_12249 ( .C (clk), .D (key_s2[96]), .Q (new_AGEMA_signal_33205) ) ;
    buf_clk new_AGEMA_reg_buffer_12253 ( .C (clk), .D (key_s3[96]), .Q (new_AGEMA_signal_33209) ) ;
    buf_clk new_AGEMA_reg_buffer_12257 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_33213) ) ;
    buf_clk new_AGEMA_reg_buffer_12261 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_33217) ) ;
    buf_clk new_AGEMA_reg_buffer_12265 ( .C (clk), .D (key_s2[97]), .Q (new_AGEMA_signal_33221) ) ;
    buf_clk new_AGEMA_reg_buffer_12269 ( .C (clk), .D (key_s3[97]), .Q (new_AGEMA_signal_33225) ) ;
    buf_clk new_AGEMA_reg_buffer_12273 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_33229) ) ;
    buf_clk new_AGEMA_reg_buffer_12277 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_33233) ) ;
    buf_clk new_AGEMA_reg_buffer_12281 ( .C (clk), .D (key_s2[98]), .Q (new_AGEMA_signal_33237) ) ;
    buf_clk new_AGEMA_reg_buffer_12285 ( .C (clk), .D (key_s3[98]), .Q (new_AGEMA_signal_33241) ) ;
    buf_clk new_AGEMA_reg_buffer_12289 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_33245) ) ;
    buf_clk new_AGEMA_reg_buffer_12293 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_33249) ) ;
    buf_clk new_AGEMA_reg_buffer_12297 ( .C (clk), .D (key_s2[99]), .Q (new_AGEMA_signal_33253) ) ;
    buf_clk new_AGEMA_reg_buffer_12301 ( .C (clk), .D (key_s3[99]), .Q (new_AGEMA_signal_33257) ) ;
    buf_clk new_AGEMA_reg_buffer_12305 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_33261) ) ;
    buf_clk new_AGEMA_reg_buffer_12309 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_33265) ) ;
    buf_clk new_AGEMA_reg_buffer_12313 ( .C (clk), .D (key_s2[100]), .Q (new_AGEMA_signal_33269) ) ;
    buf_clk new_AGEMA_reg_buffer_12317 ( .C (clk), .D (key_s3[100]), .Q (new_AGEMA_signal_33273) ) ;
    buf_clk new_AGEMA_reg_buffer_12321 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_33277) ) ;
    buf_clk new_AGEMA_reg_buffer_12325 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_33281) ) ;
    buf_clk new_AGEMA_reg_buffer_12329 ( .C (clk), .D (key_s2[101]), .Q (new_AGEMA_signal_33285) ) ;
    buf_clk new_AGEMA_reg_buffer_12333 ( .C (clk), .D (key_s3[101]), .Q (new_AGEMA_signal_33289) ) ;
    buf_clk new_AGEMA_reg_buffer_12337 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_33293) ) ;
    buf_clk new_AGEMA_reg_buffer_12341 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_33297) ) ;
    buf_clk new_AGEMA_reg_buffer_12345 ( .C (clk), .D (key_s2[102]), .Q (new_AGEMA_signal_33301) ) ;
    buf_clk new_AGEMA_reg_buffer_12349 ( .C (clk), .D (key_s3[102]), .Q (new_AGEMA_signal_33305) ) ;
    buf_clk new_AGEMA_reg_buffer_12353 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_33309) ) ;
    buf_clk new_AGEMA_reg_buffer_12357 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_33313) ) ;
    buf_clk new_AGEMA_reg_buffer_12361 ( .C (clk), .D (key_s2[103]), .Q (new_AGEMA_signal_33317) ) ;
    buf_clk new_AGEMA_reg_buffer_12365 ( .C (clk), .D (key_s3[103]), .Q (new_AGEMA_signal_33321) ) ;
    buf_clk new_AGEMA_reg_buffer_12369 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_33325) ) ;
    buf_clk new_AGEMA_reg_buffer_12373 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_33329) ) ;
    buf_clk new_AGEMA_reg_buffer_12377 ( .C (clk), .D (key_s2[104]), .Q (new_AGEMA_signal_33333) ) ;
    buf_clk new_AGEMA_reg_buffer_12381 ( .C (clk), .D (key_s3[104]), .Q (new_AGEMA_signal_33337) ) ;
    buf_clk new_AGEMA_reg_buffer_12385 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_33341) ) ;
    buf_clk new_AGEMA_reg_buffer_12389 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_33345) ) ;
    buf_clk new_AGEMA_reg_buffer_12393 ( .C (clk), .D (key_s2[105]), .Q (new_AGEMA_signal_33349) ) ;
    buf_clk new_AGEMA_reg_buffer_12397 ( .C (clk), .D (key_s3[105]), .Q (new_AGEMA_signal_33353) ) ;
    buf_clk new_AGEMA_reg_buffer_12401 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_33357) ) ;
    buf_clk new_AGEMA_reg_buffer_12405 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_33361) ) ;
    buf_clk new_AGEMA_reg_buffer_12409 ( .C (clk), .D (key_s2[106]), .Q (new_AGEMA_signal_33365) ) ;
    buf_clk new_AGEMA_reg_buffer_12413 ( .C (clk), .D (key_s3[106]), .Q (new_AGEMA_signal_33369) ) ;
    buf_clk new_AGEMA_reg_buffer_12417 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_33373) ) ;
    buf_clk new_AGEMA_reg_buffer_12421 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_33377) ) ;
    buf_clk new_AGEMA_reg_buffer_12425 ( .C (clk), .D (key_s2[107]), .Q (new_AGEMA_signal_33381) ) ;
    buf_clk new_AGEMA_reg_buffer_12429 ( .C (clk), .D (key_s3[107]), .Q (new_AGEMA_signal_33385) ) ;
    buf_clk new_AGEMA_reg_buffer_12433 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_33389) ) ;
    buf_clk new_AGEMA_reg_buffer_12437 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_33393) ) ;
    buf_clk new_AGEMA_reg_buffer_12441 ( .C (clk), .D (key_s2[108]), .Q (new_AGEMA_signal_33397) ) ;
    buf_clk new_AGEMA_reg_buffer_12445 ( .C (clk), .D (key_s3[108]), .Q (new_AGEMA_signal_33401) ) ;
    buf_clk new_AGEMA_reg_buffer_12449 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_33405) ) ;
    buf_clk new_AGEMA_reg_buffer_12453 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_33409) ) ;
    buf_clk new_AGEMA_reg_buffer_12457 ( .C (clk), .D (key_s2[109]), .Q (new_AGEMA_signal_33413) ) ;
    buf_clk new_AGEMA_reg_buffer_12461 ( .C (clk), .D (key_s3[109]), .Q (new_AGEMA_signal_33417) ) ;
    buf_clk new_AGEMA_reg_buffer_12465 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_33421) ) ;
    buf_clk new_AGEMA_reg_buffer_12469 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_33425) ) ;
    buf_clk new_AGEMA_reg_buffer_12473 ( .C (clk), .D (key_s2[110]), .Q (new_AGEMA_signal_33429) ) ;
    buf_clk new_AGEMA_reg_buffer_12477 ( .C (clk), .D (key_s3[110]), .Q (new_AGEMA_signal_33433) ) ;
    buf_clk new_AGEMA_reg_buffer_12481 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_33437) ) ;
    buf_clk new_AGEMA_reg_buffer_12485 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_33441) ) ;
    buf_clk new_AGEMA_reg_buffer_12489 ( .C (clk), .D (key_s2[111]), .Q (new_AGEMA_signal_33445) ) ;
    buf_clk new_AGEMA_reg_buffer_12493 ( .C (clk), .D (key_s3[111]), .Q (new_AGEMA_signal_33449) ) ;
    buf_clk new_AGEMA_reg_buffer_12497 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_33453) ) ;
    buf_clk new_AGEMA_reg_buffer_12501 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_33457) ) ;
    buf_clk new_AGEMA_reg_buffer_12505 ( .C (clk), .D (key_s2[112]), .Q (new_AGEMA_signal_33461) ) ;
    buf_clk new_AGEMA_reg_buffer_12509 ( .C (clk), .D (key_s3[112]), .Q (new_AGEMA_signal_33465) ) ;
    buf_clk new_AGEMA_reg_buffer_12513 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_33469) ) ;
    buf_clk new_AGEMA_reg_buffer_12517 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_33473) ) ;
    buf_clk new_AGEMA_reg_buffer_12521 ( .C (clk), .D (key_s2[113]), .Q (new_AGEMA_signal_33477) ) ;
    buf_clk new_AGEMA_reg_buffer_12525 ( .C (clk), .D (key_s3[113]), .Q (new_AGEMA_signal_33481) ) ;
    buf_clk new_AGEMA_reg_buffer_12529 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_33485) ) ;
    buf_clk new_AGEMA_reg_buffer_12533 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_33489) ) ;
    buf_clk new_AGEMA_reg_buffer_12537 ( .C (clk), .D (key_s2[114]), .Q (new_AGEMA_signal_33493) ) ;
    buf_clk new_AGEMA_reg_buffer_12541 ( .C (clk), .D (key_s3[114]), .Q (new_AGEMA_signal_33497) ) ;
    buf_clk new_AGEMA_reg_buffer_12545 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_33501) ) ;
    buf_clk new_AGEMA_reg_buffer_12549 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_33505) ) ;
    buf_clk new_AGEMA_reg_buffer_12553 ( .C (clk), .D (key_s2[115]), .Q (new_AGEMA_signal_33509) ) ;
    buf_clk new_AGEMA_reg_buffer_12557 ( .C (clk), .D (key_s3[115]), .Q (new_AGEMA_signal_33513) ) ;
    buf_clk new_AGEMA_reg_buffer_12561 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_33517) ) ;
    buf_clk new_AGEMA_reg_buffer_12565 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_33521) ) ;
    buf_clk new_AGEMA_reg_buffer_12569 ( .C (clk), .D (key_s2[116]), .Q (new_AGEMA_signal_33525) ) ;
    buf_clk new_AGEMA_reg_buffer_12573 ( .C (clk), .D (key_s3[116]), .Q (new_AGEMA_signal_33529) ) ;
    buf_clk new_AGEMA_reg_buffer_12577 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_33533) ) ;
    buf_clk new_AGEMA_reg_buffer_12581 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_33537) ) ;
    buf_clk new_AGEMA_reg_buffer_12585 ( .C (clk), .D (key_s2[117]), .Q (new_AGEMA_signal_33541) ) ;
    buf_clk new_AGEMA_reg_buffer_12589 ( .C (clk), .D (key_s3[117]), .Q (new_AGEMA_signal_33545) ) ;
    buf_clk new_AGEMA_reg_buffer_12593 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_33549) ) ;
    buf_clk new_AGEMA_reg_buffer_12597 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_33553) ) ;
    buf_clk new_AGEMA_reg_buffer_12601 ( .C (clk), .D (key_s2[118]), .Q (new_AGEMA_signal_33557) ) ;
    buf_clk new_AGEMA_reg_buffer_12605 ( .C (clk), .D (key_s3[118]), .Q (new_AGEMA_signal_33561) ) ;
    buf_clk new_AGEMA_reg_buffer_12609 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_33565) ) ;
    buf_clk new_AGEMA_reg_buffer_12613 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_33569) ) ;
    buf_clk new_AGEMA_reg_buffer_12617 ( .C (clk), .D (key_s2[119]), .Q (new_AGEMA_signal_33573) ) ;
    buf_clk new_AGEMA_reg_buffer_12621 ( .C (clk), .D (key_s3[119]), .Q (new_AGEMA_signal_33577) ) ;
    buf_clk new_AGEMA_reg_buffer_12625 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_33581) ) ;
    buf_clk new_AGEMA_reg_buffer_12629 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_33585) ) ;
    buf_clk new_AGEMA_reg_buffer_12633 ( .C (clk), .D (key_s2[120]), .Q (new_AGEMA_signal_33589) ) ;
    buf_clk new_AGEMA_reg_buffer_12637 ( .C (clk), .D (key_s3[120]), .Q (new_AGEMA_signal_33593) ) ;
    buf_clk new_AGEMA_reg_buffer_12641 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_33597) ) ;
    buf_clk new_AGEMA_reg_buffer_12645 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_33601) ) ;
    buf_clk new_AGEMA_reg_buffer_12649 ( .C (clk), .D (key_s2[121]), .Q (new_AGEMA_signal_33605) ) ;
    buf_clk new_AGEMA_reg_buffer_12653 ( .C (clk), .D (key_s3[121]), .Q (new_AGEMA_signal_33609) ) ;
    buf_clk new_AGEMA_reg_buffer_12657 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_33613) ) ;
    buf_clk new_AGEMA_reg_buffer_12661 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_33617) ) ;
    buf_clk new_AGEMA_reg_buffer_12665 ( .C (clk), .D (key_s2[122]), .Q (new_AGEMA_signal_33621) ) ;
    buf_clk new_AGEMA_reg_buffer_12669 ( .C (clk), .D (key_s3[122]), .Q (new_AGEMA_signal_33625) ) ;
    buf_clk new_AGEMA_reg_buffer_12673 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_33629) ) ;
    buf_clk new_AGEMA_reg_buffer_12677 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_33633) ) ;
    buf_clk new_AGEMA_reg_buffer_12681 ( .C (clk), .D (key_s2[123]), .Q (new_AGEMA_signal_33637) ) ;
    buf_clk new_AGEMA_reg_buffer_12685 ( .C (clk), .D (key_s3[123]), .Q (new_AGEMA_signal_33641) ) ;
    buf_clk new_AGEMA_reg_buffer_12689 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_33645) ) ;
    buf_clk new_AGEMA_reg_buffer_12693 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_33649) ) ;
    buf_clk new_AGEMA_reg_buffer_12697 ( .C (clk), .D (key_s2[124]), .Q (new_AGEMA_signal_33653) ) ;
    buf_clk new_AGEMA_reg_buffer_12701 ( .C (clk), .D (key_s3[124]), .Q (new_AGEMA_signal_33657) ) ;
    buf_clk new_AGEMA_reg_buffer_12705 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_33661) ) ;
    buf_clk new_AGEMA_reg_buffer_12709 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_33665) ) ;
    buf_clk new_AGEMA_reg_buffer_12713 ( .C (clk), .D (key_s2[125]), .Q (new_AGEMA_signal_33669) ) ;
    buf_clk new_AGEMA_reg_buffer_12717 ( .C (clk), .D (key_s3[125]), .Q (new_AGEMA_signal_33673) ) ;
    buf_clk new_AGEMA_reg_buffer_12721 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_33677) ) ;
    buf_clk new_AGEMA_reg_buffer_12725 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_33681) ) ;
    buf_clk new_AGEMA_reg_buffer_12729 ( .C (clk), .D (key_s2[126]), .Q (new_AGEMA_signal_33685) ) ;
    buf_clk new_AGEMA_reg_buffer_12733 ( .C (clk), .D (key_s3[126]), .Q (new_AGEMA_signal_33689) ) ;
    buf_clk new_AGEMA_reg_buffer_12737 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_33693) ) ;
    buf_clk new_AGEMA_reg_buffer_12741 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_33697) ) ;
    buf_clk new_AGEMA_reg_buffer_12745 ( .C (clk), .D (key_s2[127]), .Q (new_AGEMA_signal_33701) ) ;
    buf_clk new_AGEMA_reg_buffer_12749 ( .C (clk), .D (key_s3[127]), .Q (new_AGEMA_signal_33705) ) ;
    buf_clk new_AGEMA_reg_buffer_12753 ( .C (clk), .D (RoundKey[9]), .Q (new_AGEMA_signal_33709) ) ;
    buf_clk new_AGEMA_reg_buffer_12757 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_33713) ) ;
    buf_clk new_AGEMA_reg_buffer_12761 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_33717) ) ;
    buf_clk new_AGEMA_reg_buffer_12765 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_33721) ) ;
    buf_clk new_AGEMA_reg_buffer_12769 ( .C (clk), .D (RoundKey[8]), .Q (new_AGEMA_signal_33725) ) ;
    buf_clk new_AGEMA_reg_buffer_12773 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_33729) ) ;
    buf_clk new_AGEMA_reg_buffer_12777 ( .C (clk), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_33733) ) ;
    buf_clk new_AGEMA_reg_buffer_12781 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_33737) ) ;
    buf_clk new_AGEMA_reg_buffer_12785 ( .C (clk), .D (RoundKey[7]), .Q (new_AGEMA_signal_33741) ) ;
    buf_clk new_AGEMA_reg_buffer_12789 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_33745) ) ;
    buf_clk new_AGEMA_reg_buffer_12793 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_33749) ) ;
    buf_clk new_AGEMA_reg_buffer_12797 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_33753) ) ;
    buf_clk new_AGEMA_reg_buffer_12801 ( .C (clk), .D (RoundKey[6]), .Q (new_AGEMA_signal_33757) ) ;
    buf_clk new_AGEMA_reg_buffer_12805 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_33761) ) ;
    buf_clk new_AGEMA_reg_buffer_12809 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_33765) ) ;
    buf_clk new_AGEMA_reg_buffer_12813 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_33769) ) ;
    buf_clk new_AGEMA_reg_buffer_12817 ( .C (clk), .D (RoundKey[5]), .Q (new_AGEMA_signal_33773) ) ;
    buf_clk new_AGEMA_reg_buffer_12821 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_33777) ) ;
    buf_clk new_AGEMA_reg_buffer_12825 ( .C (clk), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_33781) ) ;
    buf_clk new_AGEMA_reg_buffer_12829 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_33785) ) ;
    buf_clk new_AGEMA_reg_buffer_12833 ( .C (clk), .D (RoundKey[4]), .Q (new_AGEMA_signal_33789) ) ;
    buf_clk new_AGEMA_reg_buffer_12837 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_33793) ) ;
    buf_clk new_AGEMA_reg_buffer_12841 ( .C (clk), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_33797) ) ;
    buf_clk new_AGEMA_reg_buffer_12845 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_33801) ) ;
    buf_clk new_AGEMA_reg_buffer_12849 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_33805) ) ;
    buf_clk new_AGEMA_reg_buffer_12853 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_33809) ) ;
    buf_clk new_AGEMA_reg_buffer_12857 ( .C (clk), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_33813) ) ;
    buf_clk new_AGEMA_reg_buffer_12861 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_33817) ) ;
    buf_clk new_AGEMA_reg_buffer_12865 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_33821) ) ;
    buf_clk new_AGEMA_reg_buffer_12869 ( .C (clk), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_33825) ) ;
    buf_clk new_AGEMA_reg_buffer_12873 ( .C (clk), .D (new_AGEMA_signal_5435), .Q (new_AGEMA_signal_33829) ) ;
    buf_clk new_AGEMA_reg_buffer_12877 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_33833) ) ;
    buf_clk new_AGEMA_reg_buffer_12881 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_33837) ) ;
    buf_clk new_AGEMA_reg_buffer_12885 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_33841) ) ;
    buf_clk new_AGEMA_reg_buffer_12889 ( .C (clk), .D (new_AGEMA_signal_5111), .Q (new_AGEMA_signal_33845) ) ;
    buf_clk new_AGEMA_reg_buffer_12893 ( .C (clk), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_33849) ) ;
    buf_clk new_AGEMA_reg_buffer_12897 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_33853) ) ;
    buf_clk new_AGEMA_reg_buffer_12901 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_33857) ) ;
    buf_clk new_AGEMA_reg_buffer_12905 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_33861) ) ;
    buf_clk new_AGEMA_reg_buffer_12909 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_33865) ) ;
    buf_clk new_AGEMA_reg_buffer_12913 ( .C (clk), .D (RoundKey[3]), .Q (new_AGEMA_signal_33869) ) ;
    buf_clk new_AGEMA_reg_buffer_12917 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_33873) ) ;
    buf_clk new_AGEMA_reg_buffer_12921 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_33877) ) ;
    buf_clk new_AGEMA_reg_buffer_12925 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_33881) ) ;
    buf_clk new_AGEMA_reg_buffer_12929 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_33885) ) ;
    buf_clk new_AGEMA_reg_buffer_12933 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_33889) ) ;
    buf_clk new_AGEMA_reg_buffer_12937 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_33893) ) ;
    buf_clk new_AGEMA_reg_buffer_12941 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_33897) ) ;
    buf_clk new_AGEMA_reg_buffer_12945 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_33901) ) ;
    buf_clk new_AGEMA_reg_buffer_12949 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_33905) ) ;
    buf_clk new_AGEMA_reg_buffer_12953 ( .C (clk), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_33909) ) ;
    buf_clk new_AGEMA_reg_buffer_12957 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_33913) ) ;
    buf_clk new_AGEMA_reg_buffer_12961 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_33917) ) ;
    buf_clk new_AGEMA_reg_buffer_12965 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_33921) ) ;
    buf_clk new_AGEMA_reg_buffer_12969 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_33925) ) ;
    buf_clk new_AGEMA_reg_buffer_12973 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_33929) ) ;
    buf_clk new_AGEMA_reg_buffer_12977 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_33933) ) ;
    buf_clk new_AGEMA_reg_buffer_12981 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_33937) ) ;
    buf_clk new_AGEMA_reg_buffer_12985 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_33941) ) ;
    buf_clk new_AGEMA_reg_buffer_12989 ( .C (clk), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_33945) ) ;
    buf_clk new_AGEMA_reg_buffer_12993 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_33949) ) ;
    buf_clk new_AGEMA_reg_buffer_12997 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_33953) ) ;
    buf_clk new_AGEMA_reg_buffer_13001 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_33957) ) ;
    buf_clk new_AGEMA_reg_buffer_13005 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_33961) ) ;
    buf_clk new_AGEMA_reg_buffer_13009 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_33965) ) ;
    buf_clk new_AGEMA_reg_buffer_13013 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_33969) ) ;
    buf_clk new_AGEMA_reg_buffer_13017 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_33973) ) ;
    buf_clk new_AGEMA_reg_buffer_13021 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_33977) ) ;
    buf_clk new_AGEMA_reg_buffer_13025 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_33981) ) ;
    buf_clk new_AGEMA_reg_buffer_13029 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_33985) ) ;
    buf_clk new_AGEMA_reg_buffer_13033 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_33989) ) ;
    buf_clk new_AGEMA_reg_buffer_13037 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_33993) ) ;
    buf_clk new_AGEMA_reg_buffer_13041 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_33997) ) ;
    buf_clk new_AGEMA_reg_buffer_13045 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_34001) ) ;
    buf_clk new_AGEMA_reg_buffer_13049 ( .C (clk), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_34005) ) ;
    buf_clk new_AGEMA_reg_buffer_13053 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_34009) ) ;
    buf_clk new_AGEMA_reg_buffer_13057 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_34013) ) ;
    buf_clk new_AGEMA_reg_buffer_13061 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_34017) ) ;
    buf_clk new_AGEMA_reg_buffer_13065 ( .C (clk), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_34021) ) ;
    buf_clk new_AGEMA_reg_buffer_13069 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_34025) ) ;
    buf_clk new_AGEMA_reg_buffer_13073 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_34029) ) ;
    buf_clk new_AGEMA_reg_buffer_13077 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_34033) ) ;
    buf_clk new_AGEMA_reg_buffer_13081 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_34037) ) ;
    buf_clk new_AGEMA_reg_buffer_13085 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_34041) ) ;
    buf_clk new_AGEMA_reg_buffer_13089 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_34045) ) ;
    buf_clk new_AGEMA_reg_buffer_13093 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_34049) ) ;
    buf_clk new_AGEMA_reg_buffer_13097 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_34053) ) ;
    buf_clk new_AGEMA_reg_buffer_13101 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_34057) ) ;
    buf_clk new_AGEMA_reg_buffer_13105 ( .C (clk), .D (RoundKey[31]), .Q (new_AGEMA_signal_34061) ) ;
    buf_clk new_AGEMA_reg_buffer_13109 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_34065) ) ;
    buf_clk new_AGEMA_reg_buffer_13113 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_34069) ) ;
    buf_clk new_AGEMA_reg_buffer_13117 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_34073) ) ;
    buf_clk new_AGEMA_reg_buffer_13121 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_34077) ) ;
    buf_clk new_AGEMA_reg_buffer_13125 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_34081) ) ;
    buf_clk new_AGEMA_reg_buffer_13129 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_34085) ) ;
    buf_clk new_AGEMA_reg_buffer_13133 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_34089) ) ;
    buf_clk new_AGEMA_reg_buffer_13137 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_34093) ) ;
    buf_clk new_AGEMA_reg_buffer_13141 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_34097) ) ;
    buf_clk new_AGEMA_reg_buffer_13145 ( .C (clk), .D (new_AGEMA_signal_5651), .Q (new_AGEMA_signal_34101) ) ;
    buf_clk new_AGEMA_reg_buffer_13149 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_34105) ) ;
    buf_clk new_AGEMA_reg_buffer_13153 ( .C (clk), .D (RoundKey[30]), .Q (new_AGEMA_signal_34109) ) ;
    buf_clk new_AGEMA_reg_buffer_13157 ( .C (clk), .D (new_AGEMA_signal_5011), .Q (new_AGEMA_signal_34113) ) ;
    buf_clk new_AGEMA_reg_buffer_13161 ( .C (clk), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_34117) ) ;
    buf_clk new_AGEMA_reg_buffer_13165 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_34121) ) ;
    buf_clk new_AGEMA_reg_buffer_13169 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_34125) ) ;
    buf_clk new_AGEMA_reg_buffer_13173 ( .C (clk), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_34129) ) ;
    buf_clk new_AGEMA_reg_buffer_13177 ( .C (clk), .D (new_AGEMA_signal_5327), .Q (new_AGEMA_signal_34133) ) ;
    buf_clk new_AGEMA_reg_buffer_13181 ( .C (clk), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_34137) ) ;
    buf_clk new_AGEMA_reg_buffer_13185 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_34141) ) ;
    buf_clk new_AGEMA_reg_buffer_13189 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_34145) ) ;
    buf_clk new_AGEMA_reg_buffer_13193 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_34149) ) ;
    buf_clk new_AGEMA_reg_buffer_13197 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_34153) ) ;
    buf_clk new_AGEMA_reg_buffer_13201 ( .C (clk), .D (RoundKey[2]), .Q (new_AGEMA_signal_34157) ) ;
    buf_clk new_AGEMA_reg_buffer_13205 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_34161) ) ;
    buf_clk new_AGEMA_reg_buffer_13209 ( .C (clk), .D (new_AGEMA_signal_5003), .Q (new_AGEMA_signal_34165) ) ;
    buf_clk new_AGEMA_reg_buffer_13213 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_34169) ) ;
    buf_clk new_AGEMA_reg_buffer_13217 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_34173) ) ;
    buf_clk new_AGEMA_reg_buffer_13221 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_34177) ) ;
    buf_clk new_AGEMA_reg_buffer_13225 ( .C (clk), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_34181) ) ;
    buf_clk new_AGEMA_reg_buffer_13229 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_34185) ) ;
    buf_clk new_AGEMA_reg_buffer_13233 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_34189) ) ;
    buf_clk new_AGEMA_reg_buffer_13237 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_34193) ) ;
    buf_clk new_AGEMA_reg_buffer_13241 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_34197) ) ;
    buf_clk new_AGEMA_reg_buffer_13245 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_34201) ) ;
    buf_clk new_AGEMA_reg_buffer_13249 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_34205) ) ;
    buf_clk new_AGEMA_reg_buffer_13253 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_34209) ) ;
    buf_clk new_AGEMA_reg_buffer_13257 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_34213) ) ;
    buf_clk new_AGEMA_reg_buffer_13261 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_34217) ) ;
    buf_clk new_AGEMA_reg_buffer_13265 ( .C (clk), .D (RoundKey[29]), .Q (new_AGEMA_signal_34221) ) ;
    buf_clk new_AGEMA_reg_buffer_13269 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_34225) ) ;
    buf_clk new_AGEMA_reg_buffer_13273 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_34229) ) ;
    buf_clk new_AGEMA_reg_buffer_13277 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_34233) ) ;
    buf_clk new_AGEMA_reg_buffer_13281 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_34237) ) ;
    buf_clk new_AGEMA_reg_buffer_13285 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_34241) ) ;
    buf_clk new_AGEMA_reg_buffer_13289 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_34245) ) ;
    buf_clk new_AGEMA_reg_buffer_13293 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_34249) ) ;
    buf_clk new_AGEMA_reg_buffer_13297 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_34253) ) ;
    buf_clk new_AGEMA_reg_buffer_13301 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_34257) ) ;
    buf_clk new_AGEMA_reg_buffer_13305 ( .C (clk), .D (new_AGEMA_signal_5633), .Q (new_AGEMA_signal_34261) ) ;
    buf_clk new_AGEMA_reg_buffer_13309 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_34265) ) ;
    buf_clk new_AGEMA_reg_buffer_13313 ( .C (clk), .D (RoundKey[28]), .Q (new_AGEMA_signal_34269) ) ;
    buf_clk new_AGEMA_reg_buffer_13317 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_34273) ) ;
    buf_clk new_AGEMA_reg_buffer_13321 ( .C (clk), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_34277) ) ;
    buf_clk new_AGEMA_reg_buffer_13325 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_34281) ) ;
    buf_clk new_AGEMA_reg_buffer_13329 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_34285) ) ;
    buf_clk new_AGEMA_reg_buffer_13333 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_34289) ) ;
    buf_clk new_AGEMA_reg_buffer_13337 ( .C (clk), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_34293) ) ;
    buf_clk new_AGEMA_reg_buffer_13341 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_34297) ) ;
    buf_clk new_AGEMA_reg_buffer_13345 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_34301) ) ;
    buf_clk new_AGEMA_reg_buffer_13349 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_34305) ) ;
    buf_clk new_AGEMA_reg_buffer_13353 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_34309) ) ;
    buf_clk new_AGEMA_reg_buffer_13357 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_34313) ) ;
    buf_clk new_AGEMA_reg_buffer_13361 ( .C (clk), .D (RoundKey[27]), .Q (new_AGEMA_signal_34317) ) ;
    buf_clk new_AGEMA_reg_buffer_13365 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_34321) ) ;
    buf_clk new_AGEMA_reg_buffer_13369 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_34325) ) ;
    buf_clk new_AGEMA_reg_buffer_13373 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_34329) ) ;
    buf_clk new_AGEMA_reg_buffer_13377 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_34333) ) ;
    buf_clk new_AGEMA_reg_buffer_13381 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_34337) ) ;
    buf_clk new_AGEMA_reg_buffer_13385 ( .C (clk), .D (new_AGEMA_signal_5291), .Q (new_AGEMA_signal_34341) ) ;
    buf_clk new_AGEMA_reg_buffer_13389 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_34345) ) ;
    buf_clk new_AGEMA_reg_buffer_13393 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_34349) ) ;
    buf_clk new_AGEMA_reg_buffer_13397 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_34353) ) ;
    buf_clk new_AGEMA_reg_buffer_13401 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_34357) ) ;
    buf_clk new_AGEMA_reg_buffer_13405 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_34361) ) ;
    buf_clk new_AGEMA_reg_buffer_13409 ( .C (clk), .D (RoundKey[26]), .Q (new_AGEMA_signal_34365) ) ;
    buf_clk new_AGEMA_reg_buffer_13413 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_34369) ) ;
    buf_clk new_AGEMA_reg_buffer_13417 ( .C (clk), .D (new_AGEMA_signal_4967), .Q (new_AGEMA_signal_34373) ) ;
    buf_clk new_AGEMA_reg_buffer_13421 ( .C (clk), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_34377) ) ;
    buf_clk new_AGEMA_reg_buffer_13425 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_34381) ) ;
    buf_clk new_AGEMA_reg_buffer_13429 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_34385) ) ;
    buf_clk new_AGEMA_reg_buffer_13433 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_34389) ) ;
    buf_clk new_AGEMA_reg_buffer_13437 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_34393) ) ;
    buf_clk new_AGEMA_reg_buffer_13441 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_34397) ) ;
    buf_clk new_AGEMA_reg_buffer_13445 ( .C (clk), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_34401) ) ;
    buf_clk new_AGEMA_reg_buffer_13449 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_34405) ) ;
    buf_clk new_AGEMA_reg_buffer_13453 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_34409) ) ;
    buf_clk new_AGEMA_reg_buffer_13457 ( .C (clk), .D (RoundKey[25]), .Q (new_AGEMA_signal_34413) ) ;
    buf_clk new_AGEMA_reg_buffer_13461 ( .C (clk), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_34417) ) ;
    buf_clk new_AGEMA_reg_buffer_13465 ( .C (clk), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_34421) ) ;
    buf_clk new_AGEMA_reg_buffer_13469 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_34425) ) ;
    buf_clk new_AGEMA_reg_buffer_13473 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_34429) ) ;
    buf_clk new_AGEMA_reg_buffer_13477 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_34433) ) ;
    buf_clk new_AGEMA_reg_buffer_13481 ( .C (clk), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_34437) ) ;
    buf_clk new_AGEMA_reg_buffer_13485 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_34441) ) ;
    buf_clk new_AGEMA_reg_buffer_13489 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_34445) ) ;
    buf_clk new_AGEMA_reg_buffer_13493 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_34449) ) ;
    buf_clk new_AGEMA_reg_buffer_13497 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_34453) ) ;
    buf_clk new_AGEMA_reg_buffer_13501 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_34457) ) ;
    buf_clk new_AGEMA_reg_buffer_13505 ( .C (clk), .D (RoundKey[24]), .Q (new_AGEMA_signal_34461) ) ;
    buf_clk new_AGEMA_reg_buffer_13509 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_34465) ) ;
    buf_clk new_AGEMA_reg_buffer_13513 ( .C (clk), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_34469) ) ;
    buf_clk new_AGEMA_reg_buffer_13517 ( .C (clk), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_34473) ) ;
    buf_clk new_AGEMA_reg_buffer_13521 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_34477) ) ;
    buf_clk new_AGEMA_reg_buffer_13525 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_34481) ) ;
    buf_clk new_AGEMA_reg_buffer_13529 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_34485) ) ;
    buf_clk new_AGEMA_reg_buffer_13533 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_34489) ) ;
    buf_clk new_AGEMA_reg_buffer_13537 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_34493) ) ;
    buf_clk new_AGEMA_reg_buffer_13541 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_34497) ) ;
    buf_clk new_AGEMA_reg_buffer_13545 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_34501) ) ;
    buf_clk new_AGEMA_reg_buffer_13549 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_34505) ) ;
    buf_clk new_AGEMA_reg_buffer_13553 ( .C (clk), .D (RoundKey[23]), .Q (new_AGEMA_signal_34509) ) ;
    buf_clk new_AGEMA_reg_buffer_13557 ( .C (clk), .D (new_AGEMA_signal_4939), .Q (new_AGEMA_signal_34513) ) ;
    buf_clk new_AGEMA_reg_buffer_13561 ( .C (clk), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_34517) ) ;
    buf_clk new_AGEMA_reg_buffer_13565 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_34521) ) ;
    buf_clk new_AGEMA_reg_buffer_13569 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_34525) ) ;
    buf_clk new_AGEMA_reg_buffer_13573 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_34529) ) ;
    buf_clk new_AGEMA_reg_buffer_13577 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_34533) ) ;
    buf_clk new_AGEMA_reg_buffer_13581 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_34537) ) ;
    buf_clk new_AGEMA_reg_buffer_13585 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_34541) ) ;
    buf_clk new_AGEMA_reg_buffer_13589 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_34545) ) ;
    buf_clk new_AGEMA_reg_buffer_13593 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_34549) ) ;
    buf_clk new_AGEMA_reg_buffer_13597 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_34553) ) ;
    buf_clk new_AGEMA_reg_buffer_13601 ( .C (clk), .D (RoundKey[22]), .Q (new_AGEMA_signal_34557) ) ;
    buf_clk new_AGEMA_reg_buffer_13605 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_34561) ) ;
    buf_clk new_AGEMA_reg_buffer_13609 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_34565) ) ;
    buf_clk new_AGEMA_reg_buffer_13613 ( .C (clk), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_34569) ) ;
    buf_clk new_AGEMA_reg_buffer_13617 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_34573) ) ;
    buf_clk new_AGEMA_reg_buffer_13621 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_34577) ) ;
    buf_clk new_AGEMA_reg_buffer_13625 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_34581) ) ;
    buf_clk new_AGEMA_reg_buffer_13629 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_34585) ) ;
    buf_clk new_AGEMA_reg_buffer_13633 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_34589) ) ;
    buf_clk new_AGEMA_reg_buffer_13637 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_34593) ) ;
    buf_clk new_AGEMA_reg_buffer_13641 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_34597) ) ;
    buf_clk new_AGEMA_reg_buffer_13645 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_34601) ) ;
    buf_clk new_AGEMA_reg_buffer_13649 ( .C (clk), .D (RoundKey[21]), .Q (new_AGEMA_signal_34605) ) ;
    buf_clk new_AGEMA_reg_buffer_13653 ( .C (clk), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_34609) ) ;
    buf_clk new_AGEMA_reg_buffer_13657 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_34613) ) ;
    buf_clk new_AGEMA_reg_buffer_13661 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_34617) ) ;
    buf_clk new_AGEMA_reg_buffer_13665 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_34621) ) ;
    buf_clk new_AGEMA_reg_buffer_13669 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_34625) ) ;
    buf_clk new_AGEMA_reg_buffer_13673 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_34629) ) ;
    buf_clk new_AGEMA_reg_buffer_13677 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_34633) ) ;
    buf_clk new_AGEMA_reg_buffer_13681 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_34637) ) ;
    buf_clk new_AGEMA_reg_buffer_13685 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_34641) ) ;
    buf_clk new_AGEMA_reg_buffer_13689 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_34645) ) ;
    buf_clk new_AGEMA_reg_buffer_13693 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_34649) ) ;
    buf_clk new_AGEMA_reg_buffer_13697 ( .C (clk), .D (RoundKey[20]), .Q (new_AGEMA_signal_34653) ) ;
    buf_clk new_AGEMA_reg_buffer_13701 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_34657) ) ;
    buf_clk new_AGEMA_reg_buffer_13705 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_34661) ) ;
    buf_clk new_AGEMA_reg_buffer_13709 ( .C (clk), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_34665) ) ;
    buf_clk new_AGEMA_reg_buffer_13713 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_34669) ) ;
    buf_clk new_AGEMA_reg_buffer_13717 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_34673) ) ;
    buf_clk new_AGEMA_reg_buffer_13721 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_34677) ) ;
    buf_clk new_AGEMA_reg_buffer_13725 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_34681) ) ;
    buf_clk new_AGEMA_reg_buffer_13729 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_34685) ) ;
    buf_clk new_AGEMA_reg_buffer_13733 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_34689) ) ;
    buf_clk new_AGEMA_reg_buffer_13737 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_34693) ) ;
    buf_clk new_AGEMA_reg_buffer_13741 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_34697) ) ;
    buf_clk new_AGEMA_reg_buffer_13745 ( .C (clk), .D (RoundKey[1]), .Q (new_AGEMA_signal_34701) ) ;
    buf_clk new_AGEMA_reg_buffer_13749 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_34705) ) ;
    buf_clk new_AGEMA_reg_buffer_13753 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_34709) ) ;
    buf_clk new_AGEMA_reg_buffer_13757 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_34713) ) ;
    buf_clk new_AGEMA_reg_buffer_13761 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_34717) ) ;
    buf_clk new_AGEMA_reg_buffer_13765 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_34721) ) ;
    buf_clk new_AGEMA_reg_buffer_13769 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_34725) ) ;
    buf_clk new_AGEMA_reg_buffer_13773 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_34729) ) ;
    buf_clk new_AGEMA_reg_buffer_13777 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_34733) ) ;
    buf_clk new_AGEMA_reg_buffer_13781 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_34737) ) ;
    buf_clk new_AGEMA_reg_buffer_13785 ( .C (clk), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_34741) ) ;
    buf_clk new_AGEMA_reg_buffer_13789 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_34745) ) ;
    buf_clk new_AGEMA_reg_buffer_13793 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_34749) ) ;
    buf_clk new_AGEMA_reg_buffer_13797 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_34753) ) ;
    buf_clk new_AGEMA_reg_buffer_13801 ( .C (clk), .D (new_AGEMA_signal_5669), .Q (new_AGEMA_signal_34757) ) ;
    buf_clk new_AGEMA_reg_buffer_13805 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_34761) ) ;
    buf_clk new_AGEMA_reg_buffer_13809 ( .C (clk), .D (RoundKey[19]), .Q (new_AGEMA_signal_34765) ) ;
    buf_clk new_AGEMA_reg_buffer_13813 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_34769) ) ;
    buf_clk new_AGEMA_reg_buffer_13817 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_34773) ) ;
    buf_clk new_AGEMA_reg_buffer_13821 ( .C (clk), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_34777) ) ;
    buf_clk new_AGEMA_reg_buffer_13825 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_34781) ) ;
    buf_clk new_AGEMA_reg_buffer_13829 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_34785) ) ;
    buf_clk new_AGEMA_reg_buffer_13833 ( .C (clk), .D (new_AGEMA_signal_5219), .Q (new_AGEMA_signal_34789) ) ;
    buf_clk new_AGEMA_reg_buffer_13837 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_34793) ) ;
    buf_clk new_AGEMA_reg_buffer_13841 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_34797) ) ;
    buf_clk new_AGEMA_reg_buffer_13845 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_34801) ) ;
    buf_clk new_AGEMA_reg_buffer_13849 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_34805) ) ;
    buf_clk new_AGEMA_reg_buffer_13853 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_34809) ) ;
    buf_clk new_AGEMA_reg_buffer_13857 ( .C (clk), .D (RoundKey[18]), .Q (new_AGEMA_signal_34813) ) ;
    buf_clk new_AGEMA_reg_buffer_13861 ( .C (clk), .D (new_AGEMA_signal_4885), .Q (new_AGEMA_signal_34817) ) ;
    buf_clk new_AGEMA_reg_buffer_13865 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_34821) ) ;
    buf_clk new_AGEMA_reg_buffer_13869 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_34825) ) ;
    buf_clk new_AGEMA_reg_buffer_13873 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_34829) ) ;
    buf_clk new_AGEMA_reg_buffer_13877 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_34833) ) ;
    buf_clk new_AGEMA_reg_buffer_13881 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_34837) ) ;
    buf_clk new_AGEMA_reg_buffer_13885 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_34841) ) ;
    buf_clk new_AGEMA_reg_buffer_13889 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_34845) ) ;
    buf_clk new_AGEMA_reg_buffer_13893 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_34849) ) ;
    buf_clk new_AGEMA_reg_buffer_13897 ( .C (clk), .D (new_AGEMA_signal_5525), .Q (new_AGEMA_signal_34853) ) ;
    buf_clk new_AGEMA_reg_buffer_13901 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_34857) ) ;
    buf_clk new_AGEMA_reg_buffer_13905 ( .C (clk), .D (RoundKey[17]), .Q (new_AGEMA_signal_34861) ) ;
    buf_clk new_AGEMA_reg_buffer_13909 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_34865) ) ;
    buf_clk new_AGEMA_reg_buffer_13913 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_34869) ) ;
    buf_clk new_AGEMA_reg_buffer_13917 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_34873) ) ;
    buf_clk new_AGEMA_reg_buffer_13921 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_34877) ) ;
    buf_clk new_AGEMA_reg_buffer_13925 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_34881) ) ;
    buf_clk new_AGEMA_reg_buffer_13929 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_34885) ) ;
    buf_clk new_AGEMA_reg_buffer_13933 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_34889) ) ;
    buf_clk new_AGEMA_reg_buffer_13937 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_34893) ) ;
    buf_clk new_AGEMA_reg_buffer_13941 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_34897) ) ;
    buf_clk new_AGEMA_reg_buffer_13945 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_34901) ) ;
    buf_clk new_AGEMA_reg_buffer_13949 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_34905) ) ;
    buf_clk new_AGEMA_reg_buffer_13953 ( .C (clk), .D (RoundKey[16]), .Q (new_AGEMA_signal_34909) ) ;
    buf_clk new_AGEMA_reg_buffer_13957 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (new_AGEMA_signal_34913) ) ;
    buf_clk new_AGEMA_reg_buffer_13961 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_34917) ) ;
    buf_clk new_AGEMA_reg_buffer_13965 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_34921) ) ;
    buf_clk new_AGEMA_reg_buffer_13969 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_34925) ) ;
    buf_clk new_AGEMA_reg_buffer_13973 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_34929) ) ;
    buf_clk new_AGEMA_reg_buffer_13977 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_34933) ) ;
    buf_clk new_AGEMA_reg_buffer_13981 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_34937) ) ;
    buf_clk new_AGEMA_reg_buffer_13985 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_34941) ) ;
    buf_clk new_AGEMA_reg_buffer_13989 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_34945) ) ;
    buf_clk new_AGEMA_reg_buffer_13993 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_34949) ) ;
    buf_clk new_AGEMA_reg_buffer_13997 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_34953) ) ;
    buf_clk new_AGEMA_reg_buffer_14001 ( .C (clk), .D (RoundKey[15]), .Q (new_AGEMA_signal_34957) ) ;
    buf_clk new_AGEMA_reg_buffer_14005 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_34961) ) ;
    buf_clk new_AGEMA_reg_buffer_14009 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_34965) ) ;
    buf_clk new_AGEMA_reg_buffer_14013 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_34969) ) ;
    buf_clk new_AGEMA_reg_buffer_14017 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_34973) ) ;
    buf_clk new_AGEMA_reg_buffer_14021 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_34977) ) ;
    buf_clk new_AGEMA_reg_buffer_14025 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_34981) ) ;
    buf_clk new_AGEMA_reg_buffer_14029 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_34985) ) ;
    buf_clk new_AGEMA_reg_buffer_14033 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_34989) ) ;
    buf_clk new_AGEMA_reg_buffer_14037 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_34993) ) ;
    buf_clk new_AGEMA_reg_buffer_14041 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_34997) ) ;
    buf_clk new_AGEMA_reg_buffer_14045 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_35001) ) ;
    buf_clk new_AGEMA_reg_buffer_14049 ( .C (clk), .D (RoundKey[14]), .Q (new_AGEMA_signal_35005) ) ;
    buf_clk new_AGEMA_reg_buffer_14053 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_35009) ) ;
    buf_clk new_AGEMA_reg_buffer_14057 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_35013) ) ;
    buf_clk new_AGEMA_reg_buffer_14061 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_35017) ) ;
    buf_clk new_AGEMA_reg_buffer_14065 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_35021) ) ;
    buf_clk new_AGEMA_reg_buffer_14069 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_35025) ) ;
    buf_clk new_AGEMA_reg_buffer_14073 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_35029) ) ;
    buf_clk new_AGEMA_reg_buffer_14077 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_35033) ) ;
    buf_clk new_AGEMA_reg_buffer_14081 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_35037) ) ;
    buf_clk new_AGEMA_reg_buffer_14085 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_35041) ) ;
    buf_clk new_AGEMA_reg_buffer_14089 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_35045) ) ;
    buf_clk new_AGEMA_reg_buffer_14093 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_35049) ) ;
    buf_clk new_AGEMA_reg_buffer_14097 ( .C (clk), .D (RoundKey[13]), .Q (new_AGEMA_signal_35053) ) ;
    buf_clk new_AGEMA_reg_buffer_14101 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_35057) ) ;
    buf_clk new_AGEMA_reg_buffer_14105 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_35061) ) ;
    buf_clk new_AGEMA_reg_buffer_14109 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_35065) ) ;
    buf_clk new_AGEMA_reg_buffer_14113 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_35069) ) ;
    buf_clk new_AGEMA_reg_buffer_14117 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_35073) ) ;
    buf_clk new_AGEMA_reg_buffer_14121 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_35077) ) ;
    buf_clk new_AGEMA_reg_buffer_14125 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_35081) ) ;
    buf_clk new_AGEMA_reg_buffer_14129 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_35085) ) ;
    buf_clk new_AGEMA_reg_buffer_14133 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_35089) ) ;
    buf_clk new_AGEMA_reg_buffer_14137 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_35093) ) ;
    buf_clk new_AGEMA_reg_buffer_14141 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_35097) ) ;
    buf_clk new_AGEMA_reg_buffer_14145 ( .C (clk), .D (RoundKey[12]), .Q (new_AGEMA_signal_35101) ) ;
    buf_clk new_AGEMA_reg_buffer_14149 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_35105) ) ;
    buf_clk new_AGEMA_reg_buffer_14153 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_35109) ) ;
    buf_clk new_AGEMA_reg_buffer_14157 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_35113) ) ;
    buf_clk new_AGEMA_reg_buffer_14161 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_35117) ) ;
    buf_clk new_AGEMA_reg_buffer_14165 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_35121) ) ;
    buf_clk new_AGEMA_reg_buffer_14169 ( .C (clk), .D (new_AGEMA_signal_5147), .Q (new_AGEMA_signal_35125) ) ;
    buf_clk new_AGEMA_reg_buffer_14173 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_35129) ) ;
    buf_clk new_AGEMA_reg_buffer_14177 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_35133) ) ;
    buf_clk new_AGEMA_reg_buffer_14181 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_35137) ) ;
    buf_clk new_AGEMA_reg_buffer_14185 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_35141) ) ;
    buf_clk new_AGEMA_reg_buffer_14189 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_35145) ) ;
    buf_clk new_AGEMA_reg_buffer_14193 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_35149) ) ;
    buf_clk new_AGEMA_reg_buffer_14197 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_35153) ) ;
    buf_clk new_AGEMA_reg_buffer_14201 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_35157) ) ;
    buf_clk new_AGEMA_reg_buffer_14205 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_35161) ) ;
    buf_clk new_AGEMA_reg_buffer_14209 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_35165) ) ;
    buf_clk new_AGEMA_reg_buffer_14213 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_35169) ) ;
    buf_clk new_AGEMA_reg_buffer_14217 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_35173) ) ;
    buf_clk new_AGEMA_reg_buffer_14221 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_35177) ) ;
    buf_clk new_AGEMA_reg_buffer_14225 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_35181) ) ;
    buf_clk new_AGEMA_reg_buffer_14229 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_35185) ) ;
    buf_clk new_AGEMA_reg_buffer_14233 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_35189) ) ;
    buf_clk new_AGEMA_reg_buffer_14237 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_35193) ) ;
    buf_clk new_AGEMA_reg_buffer_14241 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_35197) ) ;
    buf_clk new_AGEMA_reg_buffer_14245 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_35201) ) ;
    buf_clk new_AGEMA_reg_buffer_14249 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_35205) ) ;
    buf_clk new_AGEMA_reg_buffer_14253 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_35209) ) ;
    buf_clk new_AGEMA_reg_buffer_14257 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_35213) ) ;
    buf_clk new_AGEMA_reg_buffer_14261 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_35217) ) ;
    buf_clk new_AGEMA_reg_buffer_14265 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_35221) ) ;
    buf_clk new_AGEMA_reg_buffer_14269 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_35225) ) ;
    buf_clk new_AGEMA_reg_buffer_14273 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_35229) ) ;
    buf_clk new_AGEMA_reg_buffer_14277 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_35233) ) ;
    buf_clk new_AGEMA_reg_buffer_14281 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_35237) ) ;
    buf_clk new_AGEMA_reg_buffer_14285 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_35241) ) ;
    buf_clk new_AGEMA_reg_buffer_14289 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_35245) ) ;
    buf_clk new_AGEMA_reg_buffer_14293 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_35249) ) ;
    buf_clk new_AGEMA_reg_buffer_14297 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_35253) ) ;
    buf_clk new_AGEMA_reg_buffer_14301 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_35257) ) ;
    buf_clk new_AGEMA_reg_buffer_14305 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_35261) ) ;
    buf_clk new_AGEMA_reg_buffer_14309 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_35265) ) ;
    buf_clk new_AGEMA_reg_buffer_14313 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_35269) ) ;
    buf_clk new_AGEMA_reg_buffer_14317 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_35273) ) ;
    buf_clk new_AGEMA_reg_buffer_14321 ( .C (clk), .D (RoundKey[11]), .Q (new_AGEMA_signal_35277) ) ;
    buf_clk new_AGEMA_reg_buffer_14325 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_35281) ) ;
    buf_clk new_AGEMA_reg_buffer_14329 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_35285) ) ;
    buf_clk new_AGEMA_reg_buffer_14333 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_35289) ) ;
    buf_clk new_AGEMA_reg_buffer_14337 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_35293) ) ;
    buf_clk new_AGEMA_reg_buffer_14341 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_35297) ) ;
    buf_clk new_AGEMA_reg_buffer_14345 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_35301) ) ;
    buf_clk new_AGEMA_reg_buffer_14349 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_35305) ) ;
    buf_clk new_AGEMA_reg_buffer_14353 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_35309) ) ;
    buf_clk new_AGEMA_reg_buffer_14357 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_35313) ) ;
    buf_clk new_AGEMA_reg_buffer_14361 ( .C (clk), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_35317) ) ;
    buf_clk new_AGEMA_reg_buffer_14365 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_35321) ) ;
    buf_clk new_AGEMA_reg_buffer_14369 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_35325) ) ;
    buf_clk new_AGEMA_reg_buffer_14373 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_35329) ) ;
    buf_clk new_AGEMA_reg_buffer_14377 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_35333) ) ;
    buf_clk new_AGEMA_reg_buffer_14381 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_35337) ) ;
    buf_clk new_AGEMA_reg_buffer_14385 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_35341) ) ;
    buf_clk new_AGEMA_reg_buffer_14389 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_35345) ) ;
    buf_clk new_AGEMA_reg_buffer_14393 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_35349) ) ;
    buf_clk new_AGEMA_reg_buffer_14397 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_35353) ) ;
    buf_clk new_AGEMA_reg_buffer_14401 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_35357) ) ;
    buf_clk new_AGEMA_reg_buffer_14405 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_35361) ) ;
    buf_clk new_AGEMA_reg_buffer_14409 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_35365) ) ;
    buf_clk new_AGEMA_reg_buffer_14413 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_35369) ) ;
    buf_clk new_AGEMA_reg_buffer_14417 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_35373) ) ;
    buf_clk new_AGEMA_reg_buffer_14421 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_35377) ) ;
    buf_clk new_AGEMA_reg_buffer_14425 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_35381) ) ;
    buf_clk new_AGEMA_reg_buffer_14429 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_35385) ) ;
    buf_clk new_AGEMA_reg_buffer_14433 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_35389) ) ;
    buf_clk new_AGEMA_reg_buffer_14437 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_35393) ) ;
    buf_clk new_AGEMA_reg_buffer_14441 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_35397) ) ;
    buf_clk new_AGEMA_reg_buffer_14445 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_35401) ) ;
    buf_clk new_AGEMA_reg_buffer_14449 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_35405) ) ;
    buf_clk new_AGEMA_reg_buffer_14453 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_35409) ) ;
    buf_clk new_AGEMA_reg_buffer_14457 ( .C (clk), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_35413) ) ;
    buf_clk new_AGEMA_reg_buffer_14461 ( .C (clk), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_35417) ) ;
    buf_clk new_AGEMA_reg_buffer_14465 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_35421) ) ;
    buf_clk new_AGEMA_reg_buffer_14469 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_35425) ) ;
    buf_clk new_AGEMA_reg_buffer_14473 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_35429) ) ;
    buf_clk new_AGEMA_reg_buffer_14477 ( .C (clk), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_35433) ) ;
    buf_clk new_AGEMA_reg_buffer_14481 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_35437) ) ;
    buf_clk new_AGEMA_reg_buffer_14485 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_35441) ) ;
    buf_clk new_AGEMA_reg_buffer_14489 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_35445) ) ;
    buf_clk new_AGEMA_reg_buffer_14493 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_35449) ) ;
    buf_clk new_AGEMA_reg_buffer_14497 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_35453) ) ;
    buf_clk new_AGEMA_reg_buffer_14501 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_35457) ) ;
    buf_clk new_AGEMA_reg_buffer_14505 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_35461) ) ;
    buf_clk new_AGEMA_reg_buffer_14509 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_35465) ) ;
    buf_clk new_AGEMA_reg_buffer_14513 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_35469) ) ;
    buf_clk new_AGEMA_reg_buffer_14517 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_35473) ) ;
    buf_clk new_AGEMA_reg_buffer_14521 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_35477) ) ;
    buf_clk new_AGEMA_reg_buffer_14525 ( .C (clk), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_35481) ) ;
    buf_clk new_AGEMA_reg_buffer_14529 ( .C (clk), .D (RoundKey[10]), .Q (new_AGEMA_signal_35485) ) ;
    buf_clk new_AGEMA_reg_buffer_14533 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_35489) ) ;
    buf_clk new_AGEMA_reg_buffer_14537 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_35493) ) ;
    buf_clk new_AGEMA_reg_buffer_14541 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_35497) ) ;
    buf_clk new_AGEMA_reg_buffer_14545 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_35501) ) ;
    buf_clk new_AGEMA_reg_buffer_14549 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_35505) ) ;
    buf_clk new_AGEMA_reg_buffer_14553 ( .C (clk), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_35509) ) ;
    buf_clk new_AGEMA_reg_buffer_14557 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_35513) ) ;
    buf_clk new_AGEMA_reg_buffer_14561 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_35517) ) ;
    buf_clk new_AGEMA_reg_buffer_14565 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_35521) ) ;
    buf_clk new_AGEMA_reg_buffer_14569 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_35525) ) ;
    buf_clk new_AGEMA_reg_buffer_14573 ( .C (clk), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_35529) ) ;
    buf_clk new_AGEMA_reg_buffer_14577 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_35533) ) ;
    buf_clk new_AGEMA_reg_buffer_14581 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_35537) ) ;
    buf_clk new_AGEMA_reg_buffer_14585 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_35541) ) ;
    buf_clk new_AGEMA_reg_buffer_14589 ( .C (clk), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_35545) ) ;
    buf_clk new_AGEMA_reg_buffer_14593 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_35549) ) ;
    buf_clk new_AGEMA_reg_buffer_14597 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_35553) ) ;
    buf_clk new_AGEMA_reg_buffer_14601 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_35557) ) ;
    buf_clk new_AGEMA_reg_buffer_14605 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_35561) ) ;
    buf_clk new_AGEMA_reg_buffer_14609 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_35565) ) ;
    buf_clk new_AGEMA_reg_buffer_14613 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_35569) ) ;
    buf_clk new_AGEMA_reg_buffer_14617 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_35573) ) ;
    buf_clk new_AGEMA_reg_buffer_14621 ( .C (clk), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_35577) ) ;
    buf_clk new_AGEMA_reg_buffer_14625 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_35581) ) ;
    buf_clk new_AGEMA_reg_buffer_14629 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_35585) ) ;
    buf_clk new_AGEMA_reg_buffer_14633 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_35589) ) ;
    buf_clk new_AGEMA_reg_buffer_14637 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_35593) ) ;
    buf_clk new_AGEMA_reg_buffer_14641 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_35597) ) ;
    buf_clk new_AGEMA_reg_buffer_14645 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_35601) ) ;
    buf_clk new_AGEMA_reg_buffer_14649 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_35605) ) ;
    buf_clk new_AGEMA_reg_buffer_14653 ( .C (clk), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_35609) ) ;
    buf_clk new_AGEMA_reg_buffer_14657 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_35613) ) ;
    buf_clk new_AGEMA_reg_buffer_14661 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_35617) ) ;
    buf_clk new_AGEMA_reg_buffer_14665 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_35621) ) ;
    buf_clk new_AGEMA_reg_buffer_14669 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_35625) ) ;
    buf_clk new_AGEMA_reg_buffer_14673 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_35629) ) ;
    buf_clk new_AGEMA_reg_buffer_14677 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_35633) ) ;
    buf_clk new_AGEMA_reg_buffer_14681 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_35637) ) ;
    buf_clk new_AGEMA_reg_buffer_14685 ( .C (clk), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_35641) ) ;
    buf_clk new_AGEMA_reg_buffer_14689 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_35645) ) ;
    buf_clk new_AGEMA_reg_buffer_14693 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_35649) ) ;
    buf_clk new_AGEMA_reg_buffer_14697 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_35653) ) ;
    buf_clk new_AGEMA_reg_buffer_14701 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_35657) ) ;
    buf_clk new_AGEMA_reg_buffer_14705 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_35661) ) ;
    buf_clk new_AGEMA_reg_buffer_14709 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_35665) ) ;
    buf_clk new_AGEMA_reg_buffer_14713 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_35669) ) ;
    buf_clk new_AGEMA_reg_buffer_14717 ( .C (clk), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_35673) ) ;
    buf_clk new_AGEMA_reg_buffer_14721 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_35677) ) ;
    buf_clk new_AGEMA_reg_buffer_14725 ( .C (clk), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_35681) ) ;
    buf_clk new_AGEMA_reg_buffer_14729 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_35685) ) ;
    buf_clk new_AGEMA_reg_buffer_14733 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_35689) ) ;
    buf_clk new_AGEMA_reg_buffer_14737 ( .C (clk), .D (RoundKey[0]), .Q (new_AGEMA_signal_35693) ) ;
    buf_clk new_AGEMA_reg_buffer_14741 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_35697) ) ;
    buf_clk new_AGEMA_reg_buffer_14745 ( .C (clk), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_35701) ) ;
    buf_clk new_AGEMA_reg_buffer_14749 ( .C (clk), .D (new_AGEMA_signal_4554), .Q (new_AGEMA_signal_35705) ) ;
    buf_clk new_AGEMA_reg_buffer_14753 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_35709) ) ;
    buf_clk new_AGEMA_reg_buffer_14757 ( .C (clk), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_35713) ) ;
    buf_clk new_AGEMA_reg_buffer_14761 ( .C (clk), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_35717) ) ;
    buf_clk new_AGEMA_reg_buffer_14765 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_35721) ) ;
    buf_clk new_AGEMA_reg_buffer_14769 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_35725) ) ;
    buf_clk new_AGEMA_reg_buffer_14773 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_35729) ) ;
    buf_clk new_AGEMA_reg_buffer_14777 ( .C (clk), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_35733) ) ;
    buf_clk new_AGEMA_reg_buffer_14781 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_35737) ) ;
    buf_clk new_AGEMA_reg_buffer_14785 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_35741) ) ;
    buf_clk new_AGEMA_reg_buffer_14789 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_35745) ) ;
    buf_clk new_AGEMA_reg_buffer_14793 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_35749) ) ;
    buf_clk new_AGEMA_reg_buffer_14797 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_35753) ) ;
    buf_clk new_AGEMA_reg_buffer_14801 ( .C (clk), .D (n283), .Q (new_AGEMA_signal_35757) ) ;
    buf_clk new_AGEMA_reg_buffer_14805 ( .C (clk), .D (n285), .Q (new_AGEMA_signal_35761) ) ;
    buf_clk new_AGEMA_reg_buffer_14809 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_35765) ) ;
    buf_clk new_AGEMA_reg_buffer_14813 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_35769) ) ;
    buf_clk new_AGEMA_reg_buffer_14817 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_35773) ) ;
    buf_clk new_AGEMA_reg_buffer_14821 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_35777) ) ;
    buf_clk new_AGEMA_reg_buffer_14825 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_35781) ) ;
    buf_clk new_AGEMA_reg_buffer_14829 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_35785) ) ;
    buf_clk new_AGEMA_reg_buffer_14833 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_35789) ) ;
    buf_clk new_AGEMA_reg_buffer_14836 ( .C (clk), .D (new_AGEMA_signal_6301), .Q (new_AGEMA_signal_35792) ) ;
    buf_clk new_AGEMA_reg_buffer_14839 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_35795) ) ;
    buf_clk new_AGEMA_reg_buffer_14842 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_35798) ) ;
    buf_clk new_AGEMA_reg_buffer_14845 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_35801) ) ;
    buf_clk new_AGEMA_reg_buffer_14848 ( .C (clk), .D (new_AGEMA_signal_6781), .Q (new_AGEMA_signal_35804) ) ;
    buf_clk new_AGEMA_reg_buffer_14851 ( .C (clk), .D (new_AGEMA_signal_6782), .Q (new_AGEMA_signal_35807) ) ;
    buf_clk new_AGEMA_reg_buffer_14854 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_35810) ) ;
    buf_clk new_AGEMA_reg_buffer_14857 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_35813) ) ;
    buf_clk new_AGEMA_reg_buffer_14860 ( .C (clk), .D (new_AGEMA_signal_6313), .Q (new_AGEMA_signal_35816) ) ;
    buf_clk new_AGEMA_reg_buffer_14863 ( .C (clk), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_35819) ) ;
    buf_clk new_AGEMA_reg_buffer_14866 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_35822) ) ;
    buf_clk new_AGEMA_reg_buffer_14869 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_35825) ) ;
    buf_clk new_AGEMA_reg_buffer_14872 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_35828) ) ;
    buf_clk new_AGEMA_reg_buffer_14875 ( .C (clk), .D (new_AGEMA_signal_6305), .Q (new_AGEMA_signal_35831) ) ;
    buf_clk new_AGEMA_reg_buffer_14878 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_35834) ) ;
    buf_clk new_AGEMA_reg_buffer_14881 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_35837) ) ;
    buf_clk new_AGEMA_reg_buffer_14884 ( .C (clk), .D (new_AGEMA_signal_6790), .Q (new_AGEMA_signal_35840) ) ;
    buf_clk new_AGEMA_reg_buffer_14887 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_35843) ) ;
    buf_clk new_AGEMA_reg_buffer_14890 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_35846) ) ;
    buf_clk new_AGEMA_reg_buffer_14893 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_35849) ) ;
    buf_clk new_AGEMA_reg_buffer_14896 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_35852) ) ;
    buf_clk new_AGEMA_reg_buffer_14899 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_35855) ) ;
    buf_clk new_AGEMA_reg_buffer_14902 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_35858) ) ;
    buf_clk new_AGEMA_reg_buffer_14905 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_35861) ) ;
    buf_clk new_AGEMA_reg_buffer_14908 ( .C (clk), .D (new_AGEMA_signal_6322), .Q (new_AGEMA_signal_35864) ) ;
    buf_clk new_AGEMA_reg_buffer_14911 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_35867) ) ;
    buf_clk new_AGEMA_reg_buffer_14914 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_35870) ) ;
    buf_clk new_AGEMA_reg_buffer_14917 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_35873) ) ;
    buf_clk new_AGEMA_reg_buffer_14920 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_35876) ) ;
    buf_clk new_AGEMA_reg_buffer_14923 ( .C (clk), .D (new_AGEMA_signal_6785), .Q (new_AGEMA_signal_35879) ) ;
    buf_clk new_AGEMA_reg_buffer_14926 ( .C (clk), .D (new_AGEMA_signal_6786), .Q (new_AGEMA_signal_35882) ) ;
    buf_clk new_AGEMA_reg_buffer_14929 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_35885) ) ;
    buf_clk new_AGEMA_reg_buffer_14932 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_35888) ) ;
    buf_clk new_AGEMA_reg_buffer_14935 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_35891) ) ;
    buf_clk new_AGEMA_reg_buffer_14938 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_35894) ) ;
    buf_clk new_AGEMA_reg_buffer_14941 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_35897) ) ;
    buf_clk new_AGEMA_reg_buffer_14944 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_35900) ) ;
    buf_clk new_AGEMA_reg_buffer_14947 ( .C (clk), .D (new_AGEMA_signal_6797), .Q (new_AGEMA_signal_35903) ) ;
    buf_clk new_AGEMA_reg_buffer_14950 ( .C (clk), .D (new_AGEMA_signal_6798), .Q (new_AGEMA_signal_35906) ) ;
    buf_clk new_AGEMA_reg_buffer_14953 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_35909) ) ;
    buf_clk new_AGEMA_reg_buffer_14956 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_35912) ) ;
    buf_clk new_AGEMA_reg_buffer_14959 ( .C (clk), .D (new_AGEMA_signal_6317), .Q (new_AGEMA_signal_35915) ) ;
    buf_clk new_AGEMA_reg_buffer_14962 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_35918) ) ;
    buf_clk new_AGEMA_reg_buffer_14965 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_35921) ) ;
    buf_clk new_AGEMA_reg_buffer_14968 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_35924) ) ;
    buf_clk new_AGEMA_reg_buffer_14971 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_35927) ) ;
    buf_clk new_AGEMA_reg_buffer_14974 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_35930) ) ;
    buf_clk new_AGEMA_reg_buffer_14977 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_35933) ) ;
    buf_clk new_AGEMA_reg_buffer_14980 ( .C (clk), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_35936) ) ;
    buf_clk new_AGEMA_reg_buffer_14983 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_35939) ) ;
    buf_clk new_AGEMA_reg_buffer_14986 ( .C (clk), .D (new_AGEMA_signal_6321), .Q (new_AGEMA_signal_35942) ) ;
    buf_clk new_AGEMA_reg_buffer_14989 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_35945) ) ;
    buf_clk new_AGEMA_reg_buffer_14992 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_35948) ) ;
    buf_clk new_AGEMA_reg_buffer_14995 ( .C (clk), .D (new_AGEMA_signal_6794), .Q (new_AGEMA_signal_35951) ) ;
    buf_clk new_AGEMA_reg_buffer_14998 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_35954) ) ;
    buf_clk new_AGEMA_reg_buffer_15001 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_35957) ) ;
    buf_clk new_AGEMA_reg_buffer_15004 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_35960) ) ;
    buf_clk new_AGEMA_reg_buffer_15007 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_35963) ) ;
    buf_clk new_AGEMA_reg_buffer_15010 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_35966) ) ;
    buf_clk new_AGEMA_reg_buffer_15013 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_35969) ) ;
    buf_clk new_AGEMA_reg_buffer_15016 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_35972) ) ;
    buf_clk new_AGEMA_reg_buffer_15019 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_35975) ) ;
    buf_clk new_AGEMA_reg_buffer_15022 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_35978) ) ;
    buf_clk new_AGEMA_reg_buffer_15025 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_35981) ) ;
    buf_clk new_AGEMA_reg_buffer_15028 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_35984) ) ;
    buf_clk new_AGEMA_reg_buffer_15031 ( .C (clk), .D (new_AGEMA_signal_5705), .Q (new_AGEMA_signal_35987) ) ;
    buf_clk new_AGEMA_reg_buffer_15034 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_35990) ) ;
    buf_clk new_AGEMA_reg_buffer_15037 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_35993) ) ;
    buf_clk new_AGEMA_reg_buffer_15040 ( .C (clk), .D (new_AGEMA_signal_6325), .Q (new_AGEMA_signal_35996) ) ;
    buf_clk new_AGEMA_reg_buffer_15043 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_35999) ) ;
    buf_clk new_AGEMA_reg_buffer_15046 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_36002) ) ;
    buf_clk new_AGEMA_reg_buffer_15049 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_36005) ) ;
    buf_clk new_AGEMA_reg_buffer_15052 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_36008) ) ;
    buf_clk new_AGEMA_reg_buffer_15055 ( .C (clk), .D (new_AGEMA_signal_6821), .Q (new_AGEMA_signal_36011) ) ;
    buf_clk new_AGEMA_reg_buffer_15058 ( .C (clk), .D (new_AGEMA_signal_6822), .Q (new_AGEMA_signal_36014) ) ;
    buf_clk new_AGEMA_reg_buffer_15061 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_36017) ) ;
    buf_clk new_AGEMA_reg_buffer_15064 ( .C (clk), .D (new_AGEMA_signal_6337), .Q (new_AGEMA_signal_36020) ) ;
    buf_clk new_AGEMA_reg_buffer_15067 ( .C (clk), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_36023) ) ;
    buf_clk new_AGEMA_reg_buffer_15070 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_36026) ) ;
    buf_clk new_AGEMA_reg_buffer_15073 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_36029) ) ;
    buf_clk new_AGEMA_reg_buffer_15076 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_36032) ) ;
    buf_clk new_AGEMA_reg_buffer_15079 ( .C (clk), .D (new_AGEMA_signal_6329), .Q (new_AGEMA_signal_36035) ) ;
    buf_clk new_AGEMA_reg_buffer_15082 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_36038) ) ;
    buf_clk new_AGEMA_reg_buffer_15085 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_36041) ) ;
    buf_clk new_AGEMA_reg_buffer_15088 ( .C (clk), .D (new_AGEMA_signal_6829), .Q (new_AGEMA_signal_36044) ) ;
    buf_clk new_AGEMA_reg_buffer_15091 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_36047) ) ;
    buf_clk new_AGEMA_reg_buffer_15094 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_36050) ) ;
    buf_clk new_AGEMA_reg_buffer_15097 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_36053) ) ;
    buf_clk new_AGEMA_reg_buffer_15100 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_36056) ) ;
    buf_clk new_AGEMA_reg_buffer_15103 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_36059) ) ;
    buf_clk new_AGEMA_reg_buffer_15106 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_36062) ) ;
    buf_clk new_AGEMA_reg_buffer_15109 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_36065) ) ;
    buf_clk new_AGEMA_reg_buffer_15112 ( .C (clk), .D (new_AGEMA_signal_6346), .Q (new_AGEMA_signal_36068) ) ;
    buf_clk new_AGEMA_reg_buffer_15115 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_36071) ) ;
    buf_clk new_AGEMA_reg_buffer_15118 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_36074) ) ;
    buf_clk new_AGEMA_reg_buffer_15121 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_36077) ) ;
    buf_clk new_AGEMA_reg_buffer_15124 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_36080) ) ;
    buf_clk new_AGEMA_reg_buffer_15127 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_36083) ) ;
    buf_clk new_AGEMA_reg_buffer_15130 ( .C (clk), .D (new_AGEMA_signal_6825), .Q (new_AGEMA_signal_36086) ) ;
    buf_clk new_AGEMA_reg_buffer_15133 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_36089) ) ;
    buf_clk new_AGEMA_reg_buffer_15136 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_36092) ) ;
    buf_clk new_AGEMA_reg_buffer_15139 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_36095) ) ;
    buf_clk new_AGEMA_reg_buffer_15142 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_36098) ) ;
    buf_clk new_AGEMA_reg_buffer_15145 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_36101) ) ;
    buf_clk new_AGEMA_reg_buffer_15148 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_36104) ) ;
    buf_clk new_AGEMA_reg_buffer_15151 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_36107) ) ;
    buf_clk new_AGEMA_reg_buffer_15154 ( .C (clk), .D (new_AGEMA_signal_6837), .Q (new_AGEMA_signal_36110) ) ;
    buf_clk new_AGEMA_reg_buffer_15157 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_36113) ) ;
    buf_clk new_AGEMA_reg_buffer_15160 ( .C (clk), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_36116) ) ;
    buf_clk new_AGEMA_reg_buffer_15163 ( .C (clk), .D (new_AGEMA_signal_6341), .Q (new_AGEMA_signal_36119) ) ;
    buf_clk new_AGEMA_reg_buffer_15166 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_36122) ) ;
    buf_clk new_AGEMA_reg_buffer_15169 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_36125) ) ;
    buf_clk new_AGEMA_reg_buffer_15172 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_36128) ) ;
    buf_clk new_AGEMA_reg_buffer_15175 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_36131) ) ;
    buf_clk new_AGEMA_reg_buffer_15178 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_36134) ) ;
    buf_clk new_AGEMA_reg_buffer_15181 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_36137) ) ;
    buf_clk new_AGEMA_reg_buffer_15184 ( .C (clk), .D (new_AGEMA_signal_6343), .Q (new_AGEMA_signal_36140) ) ;
    buf_clk new_AGEMA_reg_buffer_15187 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_36143) ) ;
    buf_clk new_AGEMA_reg_buffer_15190 ( .C (clk), .D (new_AGEMA_signal_6345), .Q (new_AGEMA_signal_36146) ) ;
    buf_clk new_AGEMA_reg_buffer_15193 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_36149) ) ;
    buf_clk new_AGEMA_reg_buffer_15196 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_36152) ) ;
    buf_clk new_AGEMA_reg_buffer_15199 ( .C (clk), .D (new_AGEMA_signal_6833), .Q (new_AGEMA_signal_36155) ) ;
    buf_clk new_AGEMA_reg_buffer_15202 ( .C (clk), .D (new_AGEMA_signal_6834), .Q (new_AGEMA_signal_36158) ) ;
    buf_clk new_AGEMA_reg_buffer_15205 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_36161) ) ;
    buf_clk new_AGEMA_reg_buffer_15208 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_36164) ) ;
    buf_clk new_AGEMA_reg_buffer_15211 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_36167) ) ;
    buf_clk new_AGEMA_reg_buffer_15214 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_36170) ) ;
    buf_clk new_AGEMA_reg_buffer_15217 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_36173) ) ;
    buf_clk new_AGEMA_reg_buffer_15220 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_36176) ) ;
    buf_clk new_AGEMA_reg_buffer_15223 ( .C (clk), .D (new_AGEMA_signal_5741), .Q (new_AGEMA_signal_36179) ) ;
    buf_clk new_AGEMA_reg_buffer_15226 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_36182) ) ;
    buf_clk new_AGEMA_reg_buffer_15229 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_36185) ) ;
    buf_clk new_AGEMA_reg_buffer_15232 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_36188) ) ;
    buf_clk new_AGEMA_reg_buffer_15235 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_36191) ) ;
    buf_clk new_AGEMA_reg_buffer_15238 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_36194) ) ;
    buf_clk new_AGEMA_reg_buffer_15241 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_36197) ) ;
    buf_clk new_AGEMA_reg_buffer_15244 ( .C (clk), .D (new_AGEMA_signal_6349), .Q (new_AGEMA_signal_36200) ) ;
    buf_clk new_AGEMA_reg_buffer_15247 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_36203) ) ;
    buf_clk new_AGEMA_reg_buffer_15250 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_36206) ) ;
    buf_clk new_AGEMA_reg_buffer_15253 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_36209) ) ;
    buf_clk new_AGEMA_reg_buffer_15256 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_36212) ) ;
    buf_clk new_AGEMA_reg_buffer_15259 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_36215) ) ;
    buf_clk new_AGEMA_reg_buffer_15262 ( .C (clk), .D (new_AGEMA_signal_6861), .Q (new_AGEMA_signal_36218) ) ;
    buf_clk new_AGEMA_reg_buffer_15265 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_36221) ) ;
    buf_clk new_AGEMA_reg_buffer_15268 ( .C (clk), .D (new_AGEMA_signal_6361), .Q (new_AGEMA_signal_36224) ) ;
    buf_clk new_AGEMA_reg_buffer_15271 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_36227) ) ;
    buf_clk new_AGEMA_reg_buffer_15274 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_36230) ) ;
    buf_clk new_AGEMA_reg_buffer_15277 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_36233) ) ;
    buf_clk new_AGEMA_reg_buffer_15280 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_36236) ) ;
    buf_clk new_AGEMA_reg_buffer_15283 ( .C (clk), .D (new_AGEMA_signal_6353), .Q (new_AGEMA_signal_36239) ) ;
    buf_clk new_AGEMA_reg_buffer_15286 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_36242) ) ;
    buf_clk new_AGEMA_reg_buffer_15289 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_36245) ) ;
    buf_clk new_AGEMA_reg_buffer_15292 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_36248) ) ;
    buf_clk new_AGEMA_reg_buffer_15295 ( .C (clk), .D (new_AGEMA_signal_6869), .Q (new_AGEMA_signal_36251) ) ;
    buf_clk new_AGEMA_reg_buffer_15298 ( .C (clk), .D (new_AGEMA_signal_6870), .Q (new_AGEMA_signal_36254) ) ;
    buf_clk new_AGEMA_reg_buffer_15301 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_36257) ) ;
    buf_clk new_AGEMA_reg_buffer_15304 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_36260) ) ;
    buf_clk new_AGEMA_reg_buffer_15307 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_36263) ) ;
    buf_clk new_AGEMA_reg_buffer_15310 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_36266) ) ;
    buf_clk new_AGEMA_reg_buffer_15313 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_36269) ) ;
    buf_clk new_AGEMA_reg_buffer_15316 ( .C (clk), .D (new_AGEMA_signal_6370), .Q (new_AGEMA_signal_36272) ) ;
    buf_clk new_AGEMA_reg_buffer_15319 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_36275) ) ;
    buf_clk new_AGEMA_reg_buffer_15322 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_36278) ) ;
    buf_clk new_AGEMA_reg_buffer_15325 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_36281) ) ;
    buf_clk new_AGEMA_reg_buffer_15328 ( .C (clk), .D (new_AGEMA_signal_6862), .Q (new_AGEMA_signal_36284) ) ;
    buf_clk new_AGEMA_reg_buffer_15331 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_36287) ) ;
    buf_clk new_AGEMA_reg_buffer_15334 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_36290) ) ;
    buf_clk new_AGEMA_reg_buffer_15337 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_36293) ) ;
    buf_clk new_AGEMA_reg_buffer_15340 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_36296) ) ;
    buf_clk new_AGEMA_reg_buffer_15343 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_36299) ) ;
    buf_clk new_AGEMA_reg_buffer_15346 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_36302) ) ;
    buf_clk new_AGEMA_reg_buffer_15349 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_36305) ) ;
    buf_clk new_AGEMA_reg_buffer_15352 ( .C (clk), .D (new_AGEMA_signal_6874), .Q (new_AGEMA_signal_36308) ) ;
    buf_clk new_AGEMA_reg_buffer_15355 ( .C (clk), .D (new_AGEMA_signal_6875), .Q (new_AGEMA_signal_36311) ) ;
    buf_clk new_AGEMA_reg_buffer_15358 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_36314) ) ;
    buf_clk new_AGEMA_reg_buffer_15361 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_36317) ) ;
    buf_clk new_AGEMA_reg_buffer_15364 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_36320) ) ;
    buf_clk new_AGEMA_reg_buffer_15367 ( .C (clk), .D (new_AGEMA_signal_6365), .Q (new_AGEMA_signal_36323) ) ;
    buf_clk new_AGEMA_reg_buffer_15370 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_36326) ) ;
    buf_clk new_AGEMA_reg_buffer_15373 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_36329) ) ;
    buf_clk new_AGEMA_reg_buffer_15376 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_36332) ) ;
    buf_clk new_AGEMA_reg_buffer_15379 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_36335) ) ;
    buf_clk new_AGEMA_reg_buffer_15382 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_36338) ) ;
    buf_clk new_AGEMA_reg_buffer_15385 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_36341) ) ;
    buf_clk new_AGEMA_reg_buffer_15388 ( .C (clk), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_36344) ) ;
    buf_clk new_AGEMA_reg_buffer_15391 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_36347) ) ;
    buf_clk new_AGEMA_reg_buffer_15394 ( .C (clk), .D (new_AGEMA_signal_6369), .Q (new_AGEMA_signal_36350) ) ;
    buf_clk new_AGEMA_reg_buffer_15397 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_36353) ) ;
    buf_clk new_AGEMA_reg_buffer_15400 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_36356) ) ;
    buf_clk new_AGEMA_reg_buffer_15403 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_36359) ) ;
    buf_clk new_AGEMA_reg_buffer_15406 ( .C (clk), .D (new_AGEMA_signal_6873), .Q (new_AGEMA_signal_36362) ) ;
    buf_clk new_AGEMA_reg_buffer_15409 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_36365) ) ;
    buf_clk new_AGEMA_reg_buffer_15412 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_36368) ) ;
    buf_clk new_AGEMA_reg_buffer_15415 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_36371) ) ;
    buf_clk new_AGEMA_reg_buffer_15418 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_36374) ) ;
    buf_clk new_AGEMA_reg_buffer_15421 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_36377) ) ;
    buf_clk new_AGEMA_reg_buffer_15424 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_36380) ) ;
    buf_clk new_AGEMA_reg_buffer_15427 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_36383) ) ;
    buf_clk new_AGEMA_reg_buffer_15430 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_36386) ) ;
    buf_clk new_AGEMA_reg_buffer_15433 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_36389) ) ;
    buf_clk new_AGEMA_reg_buffer_15436 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_36392) ) ;
    buf_clk new_AGEMA_reg_buffer_15439 ( .C (clk), .D (new_AGEMA_signal_5765), .Q (new_AGEMA_signal_36395) ) ;
    buf_clk new_AGEMA_reg_buffer_15442 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_36398) ) ;
    buf_clk new_AGEMA_reg_buffer_15445 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_36401) ) ;
    buf_clk new_AGEMA_reg_buffer_15448 ( .C (clk), .D (new_AGEMA_signal_6373), .Q (new_AGEMA_signal_36404) ) ;
    buf_clk new_AGEMA_reg_buffer_15451 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_36407) ) ;
    buf_clk new_AGEMA_reg_buffer_15454 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_36410) ) ;
    buf_clk new_AGEMA_reg_buffer_15457 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_36413) ) ;
    buf_clk new_AGEMA_reg_buffer_15460 ( .C (clk), .D (new_AGEMA_signal_6898), .Q (new_AGEMA_signal_36416) ) ;
    buf_clk new_AGEMA_reg_buffer_15463 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_36419) ) ;
    buf_clk new_AGEMA_reg_buffer_15466 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_36422) ) ;
    buf_clk new_AGEMA_reg_buffer_15469 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_36425) ) ;
    buf_clk new_AGEMA_reg_buffer_15472 ( .C (clk), .D (new_AGEMA_signal_6385), .Q (new_AGEMA_signal_36428) ) ;
    buf_clk new_AGEMA_reg_buffer_15475 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_36431) ) ;
    buf_clk new_AGEMA_reg_buffer_15478 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_36434) ) ;
    buf_clk new_AGEMA_reg_buffer_15481 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_36437) ) ;
    buf_clk new_AGEMA_reg_buffer_15484 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_36440) ) ;
    buf_clk new_AGEMA_reg_buffer_15487 ( .C (clk), .D (new_AGEMA_signal_6377), .Q (new_AGEMA_signal_36443) ) ;
    buf_clk new_AGEMA_reg_buffer_15490 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_36446) ) ;
    buf_clk new_AGEMA_reg_buffer_15493 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_36449) ) ;
    buf_clk new_AGEMA_reg_buffer_15496 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_36452) ) ;
    buf_clk new_AGEMA_reg_buffer_15499 ( .C (clk), .D (new_AGEMA_signal_6908), .Q (new_AGEMA_signal_36455) ) ;
    buf_clk new_AGEMA_reg_buffer_15502 ( .C (clk), .D (new_AGEMA_signal_6909), .Q (new_AGEMA_signal_36458) ) ;
    buf_clk new_AGEMA_reg_buffer_15505 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_36461) ) ;
    buf_clk new_AGEMA_reg_buffer_15508 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_36464) ) ;
    buf_clk new_AGEMA_reg_buffer_15511 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_36467) ) ;
    buf_clk new_AGEMA_reg_buffer_15514 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_36470) ) ;
    buf_clk new_AGEMA_reg_buffer_15517 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_36473) ) ;
    buf_clk new_AGEMA_reg_buffer_15520 ( .C (clk), .D (new_AGEMA_signal_6394), .Q (new_AGEMA_signal_36476) ) ;
    buf_clk new_AGEMA_reg_buffer_15523 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_36479) ) ;
    buf_clk new_AGEMA_reg_buffer_15526 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_36482) ) ;
    buf_clk new_AGEMA_reg_buffer_15529 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_36485) ) ;
    buf_clk new_AGEMA_reg_buffer_15532 ( .C (clk), .D (new_AGEMA_signal_6901), .Q (new_AGEMA_signal_36488) ) ;
    buf_clk new_AGEMA_reg_buffer_15535 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_36491) ) ;
    buf_clk new_AGEMA_reg_buffer_15538 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_36494) ) ;
    buf_clk new_AGEMA_reg_buffer_15541 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_36497) ) ;
    buf_clk new_AGEMA_reg_buffer_15544 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_36500) ) ;
    buf_clk new_AGEMA_reg_buffer_15547 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_36503) ) ;
    buf_clk new_AGEMA_reg_buffer_15550 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_36506) ) ;
    buf_clk new_AGEMA_reg_buffer_15553 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_36509) ) ;
    buf_clk new_AGEMA_reg_buffer_15556 ( .C (clk), .D (new_AGEMA_signal_6913), .Q (new_AGEMA_signal_36512) ) ;
    buf_clk new_AGEMA_reg_buffer_15559 ( .C (clk), .D (new_AGEMA_signal_6914), .Q (new_AGEMA_signal_36515) ) ;
    buf_clk new_AGEMA_reg_buffer_15562 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_36518) ) ;
    buf_clk new_AGEMA_reg_buffer_15565 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_36521) ) ;
    buf_clk new_AGEMA_reg_buffer_15568 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_36524) ) ;
    buf_clk new_AGEMA_reg_buffer_15571 ( .C (clk), .D (new_AGEMA_signal_6389), .Q (new_AGEMA_signal_36527) ) ;
    buf_clk new_AGEMA_reg_buffer_15574 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_36530) ) ;
    buf_clk new_AGEMA_reg_buffer_15577 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_36533) ) ;
    buf_clk new_AGEMA_reg_buffer_15580 ( .C (clk), .D (new_AGEMA_signal_5797), .Q (new_AGEMA_signal_36536) ) ;
    buf_clk new_AGEMA_reg_buffer_15583 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_36539) ) ;
    buf_clk new_AGEMA_reg_buffer_15586 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_36542) ) ;
    buf_clk new_AGEMA_reg_buffer_15589 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_36545) ) ;
    buf_clk new_AGEMA_reg_buffer_15592 ( .C (clk), .D (new_AGEMA_signal_6391), .Q (new_AGEMA_signal_36548) ) ;
    buf_clk new_AGEMA_reg_buffer_15595 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_36551) ) ;
    buf_clk new_AGEMA_reg_buffer_15598 ( .C (clk), .D (new_AGEMA_signal_6393), .Q (new_AGEMA_signal_36554) ) ;
    buf_clk new_AGEMA_reg_buffer_15601 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_36557) ) ;
    buf_clk new_AGEMA_reg_buffer_15604 ( .C (clk), .D (new_AGEMA_signal_6910), .Q (new_AGEMA_signal_36560) ) ;
    buf_clk new_AGEMA_reg_buffer_15607 ( .C (clk), .D (new_AGEMA_signal_6911), .Q (new_AGEMA_signal_36563) ) ;
    buf_clk new_AGEMA_reg_buffer_15610 ( .C (clk), .D (new_AGEMA_signal_6912), .Q (new_AGEMA_signal_36566) ) ;
    buf_clk new_AGEMA_reg_buffer_15613 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_36569) ) ;
    buf_clk new_AGEMA_reg_buffer_15616 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_36572) ) ;
    buf_clk new_AGEMA_reg_buffer_15619 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_36575) ) ;
    buf_clk new_AGEMA_reg_buffer_15622 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_36578) ) ;
    buf_clk new_AGEMA_reg_buffer_15625 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_36581) ) ;
    buf_clk new_AGEMA_reg_buffer_15628 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_36584) ) ;
    buf_clk new_AGEMA_reg_buffer_15631 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_36587) ) ;
    buf_clk new_AGEMA_reg_buffer_15634 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_36590) ) ;
    buf_clk new_AGEMA_reg_buffer_15637 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_36593) ) ;
    buf_clk new_AGEMA_reg_buffer_15640 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_36596) ) ;
    buf_clk new_AGEMA_reg_buffer_15643 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_36599) ) ;
    buf_clk new_AGEMA_reg_buffer_15646 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_36602) ) ;
    buf_clk new_AGEMA_reg_buffer_15649 ( .C (clk), .D (RoundCounterIns_N7), .Q (new_AGEMA_signal_36605) ) ;
    buf_clk new_AGEMA_reg_buffer_15653 ( .C (clk), .D (RoundCounterIns_N8), .Q (new_AGEMA_signal_36609) ) ;
    buf_clk new_AGEMA_reg_buffer_15657 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_36613) ) ;
    buf_clk new_AGEMA_reg_buffer_15661 ( .C (clk), .D (RoundCounterIns_N10), .Q (new_AGEMA_signal_36617) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_25488, new_AGEMA_signal_25487, new_AGEMA_signal_25486, new_AGEMA_signal_25485}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, new_AGEMA_signal_8944, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_25492, new_AGEMA_signal_25491, new_AGEMA_signal_25490, new_AGEMA_signal_25489}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, new_AGEMA_signal_8950, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_25496, new_AGEMA_signal_25495, new_AGEMA_signal_25494, new_AGEMA_signal_25493}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8955, new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190], Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, new_AGEMA_signal_8698, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_25500, new_AGEMA_signal_25499, new_AGEMA_signal_25498, new_AGEMA_signal_25497}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_9255, new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_25504, new_AGEMA_signal_25503, new_AGEMA_signal_25502, new_AGEMA_signal_25501}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, new_AGEMA_signal_8959, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_25508, new_AGEMA_signal_25507, new_AGEMA_signal_25506, new_AGEMA_signal_25505}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, new_AGEMA_signal_8962, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, new_AGEMA_signal_8965, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_25512, new_AGEMA_signal_25511, new_AGEMA_signal_25510, new_AGEMA_signal_25509}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, new_AGEMA_signal_8968, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, new_AGEMA_signal_8710, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_25516, new_AGEMA_signal_25515, new_AGEMA_signal_25514, new_AGEMA_signal_25513}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, new_AGEMA_signal_9268, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_25520, new_AGEMA_signal_25519, new_AGEMA_signal_25518, new_AGEMA_signal_25517}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, new_AGEMA_signal_8974, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_25524, new_AGEMA_signal_25523, new_AGEMA_signal_25522, new_AGEMA_signal_25521}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, new_AGEMA_signal_8977, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250], Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, new_AGEMA_signal_8980, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_25528, new_AGEMA_signal_25527, new_AGEMA_signal_25526, new_AGEMA_signal_25525}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8985, new_AGEMA_signal_8984, new_AGEMA_signal_8983, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, new_AGEMA_signal_8722, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_25532, new_AGEMA_signal_25531, new_AGEMA_signal_25530, new_AGEMA_signal_25529}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_9285, new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_25536, new_AGEMA_signal_25535, new_AGEMA_signal_25534, new_AGEMA_signal_25533}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, new_AGEMA_signal_8989, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_25540, new_AGEMA_signal_25539, new_AGEMA_signal_25538, new_AGEMA_signal_25537}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, new_AGEMA_signal_8992, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, new_AGEMA_signal_8995, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_25544, new_AGEMA_signal_25543, new_AGEMA_signal_25542, new_AGEMA_signal_25541}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, new_AGEMA_signal_8998, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, new_AGEMA_signal_8734, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_25548, new_AGEMA_signal_25547, new_AGEMA_signal_25546, new_AGEMA_signal_25545}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, new_AGEMA_signal_9298, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310], Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_25552, new_AGEMA_signal_25551, new_AGEMA_signal_25550, new_AGEMA_signal_25549}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, new_AGEMA_signal_9004, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_25556, new_AGEMA_signal_25555, new_AGEMA_signal_25554, new_AGEMA_signal_25553}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, new_AGEMA_signal_9007, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, new_AGEMA_signal_9010, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_25560, new_AGEMA_signal_25559, new_AGEMA_signal_25558, new_AGEMA_signal_25557}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9015, new_AGEMA_signal_9014, new_AGEMA_signal_9013, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, new_AGEMA_signal_8746, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_25564, new_AGEMA_signal_25563, new_AGEMA_signal_25562, new_AGEMA_signal_25561}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_25568, new_AGEMA_signal_25567, new_AGEMA_signal_25566, new_AGEMA_signal_25565}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, new_AGEMA_signal_9019, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_25572, new_AGEMA_signal_25571, new_AGEMA_signal_25570, new_AGEMA_signal_25569}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, new_AGEMA_signal_9022, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, new_AGEMA_signal_9025, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_25576, new_AGEMA_signal_25575, new_AGEMA_signal_25574, new_AGEMA_signal_25573}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, new_AGEMA_signal_9028, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370], Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, new_AGEMA_signal_8758, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_25580, new_AGEMA_signal_25579, new_AGEMA_signal_25578, new_AGEMA_signal_25577}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, new_AGEMA_signal_9328, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_25584, new_AGEMA_signal_25583, new_AGEMA_signal_25582, new_AGEMA_signal_25581}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, new_AGEMA_signal_9034, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_25588, new_AGEMA_signal_25587, new_AGEMA_signal_25586, new_AGEMA_signal_25585}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, new_AGEMA_signal_9040, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_25592, new_AGEMA_signal_25591, new_AGEMA_signal_25590, new_AGEMA_signal_25589}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9045, new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, new_AGEMA_signal_8770, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_25596, new_AGEMA_signal_25595, new_AGEMA_signal_25594, new_AGEMA_signal_25593}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9345, new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_25600, new_AGEMA_signal_25599, new_AGEMA_signal_25598, new_AGEMA_signal_25597}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_25604, new_AGEMA_signal_25603, new_AGEMA_signal_25602, new_AGEMA_signal_25601}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, new_AGEMA_signal_9052, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430], Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_25608, new_AGEMA_signal_25607, new_AGEMA_signal_25606, new_AGEMA_signal_25605}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, new_AGEMA_signal_9058, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, new_AGEMA_signal_8782, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_25612, new_AGEMA_signal_25611, new_AGEMA_signal_25610, new_AGEMA_signal_25609}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, new_AGEMA_signal_9358, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_25616, new_AGEMA_signal_25615, new_AGEMA_signal_25614, new_AGEMA_signal_25613}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, new_AGEMA_signal_9064, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_25620, new_AGEMA_signal_25619, new_AGEMA_signal_25618, new_AGEMA_signal_25617}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, new_AGEMA_signal_9070, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_25624, new_AGEMA_signal_25623, new_AGEMA_signal_25622, new_AGEMA_signal_25621}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, new_AGEMA_signal_8794, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_25628, new_AGEMA_signal_25627, new_AGEMA_signal_25626, new_AGEMA_signal_25625}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9375, new_AGEMA_signal_9374, new_AGEMA_signal_9373, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490], Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_25632, new_AGEMA_signal_25631, new_AGEMA_signal_25630, new_AGEMA_signal_25629}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_25636, new_AGEMA_signal_25635, new_AGEMA_signal_25634, new_AGEMA_signal_25633}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, new_AGEMA_signal_9082, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_25640, new_AGEMA_signal_25639, new_AGEMA_signal_25638, new_AGEMA_signal_25637}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, new_AGEMA_signal_9088, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, new_AGEMA_signal_8806, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_25644, new_AGEMA_signal_25643, new_AGEMA_signal_25642, new_AGEMA_signal_25641}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, new_AGEMA_signal_9388, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_25648, new_AGEMA_signal_25647, new_AGEMA_signal_25646, new_AGEMA_signal_25645}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, new_AGEMA_signal_9094, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_25652, new_AGEMA_signal_25651, new_AGEMA_signal_25650, new_AGEMA_signal_25649}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, new_AGEMA_signal_9100, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_25656, new_AGEMA_signal_25655, new_AGEMA_signal_25654, new_AGEMA_signal_25653}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9105, new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550], Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, new_AGEMA_signal_8818, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_25660, new_AGEMA_signal_25659, new_AGEMA_signal_25658, new_AGEMA_signal_25657}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, new_AGEMA_signal_9403, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_25664, new_AGEMA_signal_25663, new_AGEMA_signal_25662, new_AGEMA_signal_25661}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_25668, new_AGEMA_signal_25667, new_AGEMA_signal_25666, new_AGEMA_signal_25665}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, new_AGEMA_signal_9112, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_25672, new_AGEMA_signal_25671, new_AGEMA_signal_25670, new_AGEMA_signal_25669}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, new_AGEMA_signal_9118, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, new_AGEMA_signal_8830, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_25676, new_AGEMA_signal_25675, new_AGEMA_signal_25674, new_AGEMA_signal_25673}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, new_AGEMA_signal_9418, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_25680, new_AGEMA_signal_25679, new_AGEMA_signal_25678, new_AGEMA_signal_25677}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, new_AGEMA_signal_9124, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_25684, new_AGEMA_signal_25683, new_AGEMA_signal_25682, new_AGEMA_signal_25681}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610], Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, new_AGEMA_signal_9130, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_25688, new_AGEMA_signal_25687, new_AGEMA_signal_25686, new_AGEMA_signal_25685}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9135, new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, new_AGEMA_signal_8842, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_25692, new_AGEMA_signal_25691, new_AGEMA_signal_25690, new_AGEMA_signal_25689}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9435, new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_25696, new_AGEMA_signal_25695, new_AGEMA_signal_25694, new_AGEMA_signal_25693}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_25700, new_AGEMA_signal_25699, new_AGEMA_signal_25698, new_AGEMA_signal_25697}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, new_AGEMA_signal_9142, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_25704, new_AGEMA_signal_25703, new_AGEMA_signal_25702, new_AGEMA_signal_25701}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, new_AGEMA_signal_9148, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, new_AGEMA_signal_8854, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_25708, new_AGEMA_signal_25707, new_AGEMA_signal_25706, new_AGEMA_signal_25705}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, new_AGEMA_signal_9448, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670], Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_25712, new_AGEMA_signal_25711, new_AGEMA_signal_25710, new_AGEMA_signal_25709}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, new_AGEMA_signal_9154, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_25716, new_AGEMA_signal_25715, new_AGEMA_signal_25714, new_AGEMA_signal_25713}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, new_AGEMA_signal_9160, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_25720, new_AGEMA_signal_25719, new_AGEMA_signal_25718, new_AGEMA_signal_25717}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9165, new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, new_AGEMA_signal_8866, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_25724, new_AGEMA_signal_25723, new_AGEMA_signal_25722, new_AGEMA_signal_25721}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_25728, new_AGEMA_signal_25727, new_AGEMA_signal_25726, new_AGEMA_signal_25725}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_25732, new_AGEMA_signal_25731, new_AGEMA_signal_25730, new_AGEMA_signal_25729}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, new_AGEMA_signal_9172, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_25736, new_AGEMA_signal_25735, new_AGEMA_signal_25734, new_AGEMA_signal_25733}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, new_AGEMA_signal_9178, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730], Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, new_AGEMA_signal_8878, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_25740, new_AGEMA_signal_25739, new_AGEMA_signal_25738, new_AGEMA_signal_25737}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, new_AGEMA_signal_9478, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_25744, new_AGEMA_signal_25743, new_AGEMA_signal_25742, new_AGEMA_signal_25741}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, new_AGEMA_signal_8884, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_25748, new_AGEMA_signal_25747, new_AGEMA_signal_25746, new_AGEMA_signal_25745}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, new_AGEMA_signal_8887, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, new_AGEMA_signal_8890, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_25752, new_AGEMA_signal_25751, new_AGEMA_signal_25750, new_AGEMA_signal_25749}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8895, new_AGEMA_signal_8894, new_AGEMA_signal_8893, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, new_AGEMA_signal_8650, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_25756, new_AGEMA_signal_25755, new_AGEMA_signal_25754, new_AGEMA_signal_25753}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, new_AGEMA_signal_9193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_25760, new_AGEMA_signal_25759, new_AGEMA_signal_25758, new_AGEMA_signal_25757}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, new_AGEMA_signal_8899, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_25764, new_AGEMA_signal_25763, new_AGEMA_signal_25762, new_AGEMA_signal_25761}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, new_AGEMA_signal_8902, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790], Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, new_AGEMA_signal_8905, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_25768, new_AGEMA_signal_25767, new_AGEMA_signal_25766, new_AGEMA_signal_25765}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, new_AGEMA_signal_8908, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, new_AGEMA_signal_8662, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_25772, new_AGEMA_signal_25771, new_AGEMA_signal_25770, new_AGEMA_signal_25769}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, new_AGEMA_signal_9208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_25776, new_AGEMA_signal_25775, new_AGEMA_signal_25774, new_AGEMA_signal_25773}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, new_AGEMA_signal_8914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_25780, new_AGEMA_signal_25779, new_AGEMA_signal_25778, new_AGEMA_signal_25777}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, new_AGEMA_signal_8917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, new_AGEMA_signal_8920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_25784, new_AGEMA_signal_25783, new_AGEMA_signal_25782, new_AGEMA_signal_25781}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, new_AGEMA_signal_8923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, new_AGEMA_signal_8674, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_25788, new_AGEMA_signal_25787, new_AGEMA_signal_25786, new_AGEMA_signal_25785}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_9225, new_AGEMA_signal_9224, new_AGEMA_signal_9223, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850], Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_25792, new_AGEMA_signal_25791, new_AGEMA_signal_25790, new_AGEMA_signal_25789}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, new_AGEMA_signal_8929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_25796, new_AGEMA_signal_25795, new_AGEMA_signal_25794, new_AGEMA_signal_25793}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, new_AGEMA_signal_8932, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, new_AGEMA_signal_8935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_25800, new_AGEMA_signal_25799, new_AGEMA_signal_25798, new_AGEMA_signal_25797}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, new_AGEMA_signal_8938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, new_AGEMA_signal_8686, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_25804, new_AGEMA_signal_25803, new_AGEMA_signal_25802, new_AGEMA_signal_25801}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, new_AGEMA_signal_9238, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_25485) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_8455), .Q (new_AGEMA_signal_25486) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_8456), .Q (new_AGEMA_signal_25487) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_8457), .Q (new_AGEMA_signal_25488) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_25489) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_8689), .Q (new_AGEMA_signal_25490) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_8690), .Q (new_AGEMA_signal_25491) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_8691), .Q (new_AGEMA_signal_25492) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_25493) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_8695), .Q (new_AGEMA_signal_25494) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_8696), .Q (new_AGEMA_signal_25495) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_8697), .Q (new_AGEMA_signal_25496) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_25497) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_8941), .Q (new_AGEMA_signal_25498) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_8942), .Q (new_AGEMA_signal_25499) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_8943), .Q (new_AGEMA_signal_25500) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_25501) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_8467), .Q (new_AGEMA_signal_25502) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_8468), .Q (new_AGEMA_signal_25503) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_8469), .Q (new_AGEMA_signal_25504) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_25505) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_8701), .Q (new_AGEMA_signal_25506) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_8702), .Q (new_AGEMA_signal_25507) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_8703), .Q (new_AGEMA_signal_25508) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_25509) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_8707), .Q (new_AGEMA_signal_25510) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_8708), .Q (new_AGEMA_signal_25511) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_8709), .Q (new_AGEMA_signal_25512) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_25513) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_8956), .Q (new_AGEMA_signal_25514) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_8957), .Q (new_AGEMA_signal_25515) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_8958), .Q (new_AGEMA_signal_25516) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_25517) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_8479), .Q (new_AGEMA_signal_25518) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_8480), .Q (new_AGEMA_signal_25519) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_8481), .Q (new_AGEMA_signal_25520) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_25521) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_8713), .Q (new_AGEMA_signal_25522) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_8714), .Q (new_AGEMA_signal_25523) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_8715), .Q (new_AGEMA_signal_25524) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_25525) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_8719), .Q (new_AGEMA_signal_25526) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_8720), .Q (new_AGEMA_signal_25527) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_8721), .Q (new_AGEMA_signal_25528) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_25529) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_8971), .Q (new_AGEMA_signal_25530) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_8972), .Q (new_AGEMA_signal_25531) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_8973), .Q (new_AGEMA_signal_25532) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_25533) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_8491), .Q (new_AGEMA_signal_25534) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_8492), .Q (new_AGEMA_signal_25535) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_8493), .Q (new_AGEMA_signal_25536) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_25537) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_8725), .Q (new_AGEMA_signal_25538) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_8726), .Q (new_AGEMA_signal_25539) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_8727), .Q (new_AGEMA_signal_25540) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_25541) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_8731), .Q (new_AGEMA_signal_25542) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_8732), .Q (new_AGEMA_signal_25543) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_8733), .Q (new_AGEMA_signal_25544) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_25545) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_8986), .Q (new_AGEMA_signal_25546) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_8987), .Q (new_AGEMA_signal_25547) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_8988), .Q (new_AGEMA_signal_25548) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M21), .Q (new_AGEMA_signal_25549) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_8503), .Q (new_AGEMA_signal_25550) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_8504), .Q (new_AGEMA_signal_25551) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_8505), .Q (new_AGEMA_signal_25552) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M23), .Q (new_AGEMA_signal_25553) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_8737), .Q (new_AGEMA_signal_25554) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_8738), .Q (new_AGEMA_signal_25555) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_8739), .Q (new_AGEMA_signal_25556) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M27), .Q (new_AGEMA_signal_25557) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_8743), .Q (new_AGEMA_signal_25558) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_8744), .Q (new_AGEMA_signal_25559) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_8745), .Q (new_AGEMA_signal_25560) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M24), .Q (new_AGEMA_signal_25561) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_9001), .Q (new_AGEMA_signal_25562) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_9002), .Q (new_AGEMA_signal_25563) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_9003), .Q (new_AGEMA_signal_25564) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M21), .Q (new_AGEMA_signal_25565) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_8515), .Q (new_AGEMA_signal_25566) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_8516), .Q (new_AGEMA_signal_25567) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_8517), .Q (new_AGEMA_signal_25568) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M23), .Q (new_AGEMA_signal_25569) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_8749), .Q (new_AGEMA_signal_25570) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_8750), .Q (new_AGEMA_signal_25571) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_8751), .Q (new_AGEMA_signal_25572) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M27), .Q (new_AGEMA_signal_25573) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_8755), .Q (new_AGEMA_signal_25574) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_8756), .Q (new_AGEMA_signal_25575) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_8757), .Q (new_AGEMA_signal_25576) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M24), .Q (new_AGEMA_signal_25577) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_9016), .Q (new_AGEMA_signal_25578) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_9017), .Q (new_AGEMA_signal_25579) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_9018), .Q (new_AGEMA_signal_25580) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M21), .Q (new_AGEMA_signal_25581) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_8527), .Q (new_AGEMA_signal_25582) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_8528), .Q (new_AGEMA_signal_25583) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_8529), .Q (new_AGEMA_signal_25584) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M23), .Q (new_AGEMA_signal_25585) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_8761), .Q (new_AGEMA_signal_25586) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_8762), .Q (new_AGEMA_signal_25587) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_8763), .Q (new_AGEMA_signal_25588) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M27), .Q (new_AGEMA_signal_25589) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_8767), .Q (new_AGEMA_signal_25590) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_8768), .Q (new_AGEMA_signal_25591) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_8769), .Q (new_AGEMA_signal_25592) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M24), .Q (new_AGEMA_signal_25593) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_9031), .Q (new_AGEMA_signal_25594) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_9032), .Q (new_AGEMA_signal_25595) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_9033), .Q (new_AGEMA_signal_25596) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M21), .Q (new_AGEMA_signal_25597) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_8539), .Q (new_AGEMA_signal_25598) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_8540), .Q (new_AGEMA_signal_25599) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_8541), .Q (new_AGEMA_signal_25600) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M23), .Q (new_AGEMA_signal_25601) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_8773), .Q (new_AGEMA_signal_25602) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_8774), .Q (new_AGEMA_signal_25603) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_8775), .Q (new_AGEMA_signal_25604) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M27), .Q (new_AGEMA_signal_25605) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_8779), .Q (new_AGEMA_signal_25606) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_8780), .Q (new_AGEMA_signal_25607) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_8781), .Q (new_AGEMA_signal_25608) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M24), .Q (new_AGEMA_signal_25609) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_9046), .Q (new_AGEMA_signal_25610) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_9047), .Q (new_AGEMA_signal_25611) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_9048), .Q (new_AGEMA_signal_25612) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M21), .Q (new_AGEMA_signal_25613) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_8551), .Q (new_AGEMA_signal_25614) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_8552), .Q (new_AGEMA_signal_25615) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_8553), .Q (new_AGEMA_signal_25616) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M23), .Q (new_AGEMA_signal_25617) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_8785), .Q (new_AGEMA_signal_25618) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_8786), .Q (new_AGEMA_signal_25619) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_8787), .Q (new_AGEMA_signal_25620) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M27), .Q (new_AGEMA_signal_25621) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_8791), .Q (new_AGEMA_signal_25622) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_8792), .Q (new_AGEMA_signal_25623) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_8793), .Q (new_AGEMA_signal_25624) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M24), .Q (new_AGEMA_signal_25625) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_9061), .Q (new_AGEMA_signal_25626) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_9062), .Q (new_AGEMA_signal_25627) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_9063), .Q (new_AGEMA_signal_25628) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M21), .Q (new_AGEMA_signal_25629) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_8563), .Q (new_AGEMA_signal_25630) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_8564), .Q (new_AGEMA_signal_25631) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_8565), .Q (new_AGEMA_signal_25632) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M23), .Q (new_AGEMA_signal_25633) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_8797), .Q (new_AGEMA_signal_25634) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_8798), .Q (new_AGEMA_signal_25635) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_8799), .Q (new_AGEMA_signal_25636) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M27), .Q (new_AGEMA_signal_25637) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_8803), .Q (new_AGEMA_signal_25638) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_8804), .Q (new_AGEMA_signal_25639) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_8805), .Q (new_AGEMA_signal_25640) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M24), .Q (new_AGEMA_signal_25641) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_9076), .Q (new_AGEMA_signal_25642) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_9077), .Q (new_AGEMA_signal_25643) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_9078), .Q (new_AGEMA_signal_25644) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M21), .Q (new_AGEMA_signal_25645) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_8575), .Q (new_AGEMA_signal_25646) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_8576), .Q (new_AGEMA_signal_25647) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_8577), .Q (new_AGEMA_signal_25648) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M23), .Q (new_AGEMA_signal_25649) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_8809), .Q (new_AGEMA_signal_25650) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_8810), .Q (new_AGEMA_signal_25651) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_8811), .Q (new_AGEMA_signal_25652) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M27), .Q (new_AGEMA_signal_25653) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_8815), .Q (new_AGEMA_signal_25654) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_8816), .Q (new_AGEMA_signal_25655) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_8817), .Q (new_AGEMA_signal_25656) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M24), .Q (new_AGEMA_signal_25657) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_9091), .Q (new_AGEMA_signal_25658) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_9092), .Q (new_AGEMA_signal_25659) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_9093), .Q (new_AGEMA_signal_25660) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M21), .Q (new_AGEMA_signal_25661) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_8587), .Q (new_AGEMA_signal_25662) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_8588), .Q (new_AGEMA_signal_25663) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_8589), .Q (new_AGEMA_signal_25664) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M23), .Q (new_AGEMA_signal_25665) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_8821), .Q (new_AGEMA_signal_25666) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_8822), .Q (new_AGEMA_signal_25667) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_8823), .Q (new_AGEMA_signal_25668) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M27), .Q (new_AGEMA_signal_25669) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_8827), .Q (new_AGEMA_signal_25670) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_8828), .Q (new_AGEMA_signal_25671) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_8829), .Q (new_AGEMA_signal_25672) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M24), .Q (new_AGEMA_signal_25673) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_9106), .Q (new_AGEMA_signal_25674) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_9107), .Q (new_AGEMA_signal_25675) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_9108), .Q (new_AGEMA_signal_25676) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M21), .Q (new_AGEMA_signal_25677) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_8599), .Q (new_AGEMA_signal_25678) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_8600), .Q (new_AGEMA_signal_25679) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_8601), .Q (new_AGEMA_signal_25680) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M23), .Q (new_AGEMA_signal_25681) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_8833), .Q (new_AGEMA_signal_25682) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_8834), .Q (new_AGEMA_signal_25683) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_8835), .Q (new_AGEMA_signal_25684) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M27), .Q (new_AGEMA_signal_25685) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_8839), .Q (new_AGEMA_signal_25686) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_8840), .Q (new_AGEMA_signal_25687) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_8841), .Q (new_AGEMA_signal_25688) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M24), .Q (new_AGEMA_signal_25689) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_9121), .Q (new_AGEMA_signal_25690) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_9122), .Q (new_AGEMA_signal_25691) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_9123), .Q (new_AGEMA_signal_25692) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M21), .Q (new_AGEMA_signal_25693) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_8611), .Q (new_AGEMA_signal_25694) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_8612), .Q (new_AGEMA_signal_25695) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_8613), .Q (new_AGEMA_signal_25696) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M23), .Q (new_AGEMA_signal_25697) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_8845), .Q (new_AGEMA_signal_25698) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_8846), .Q (new_AGEMA_signal_25699) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_8847), .Q (new_AGEMA_signal_25700) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M27), .Q (new_AGEMA_signal_25701) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_8851), .Q (new_AGEMA_signal_25702) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_8852), .Q (new_AGEMA_signal_25703) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_8853), .Q (new_AGEMA_signal_25704) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M24), .Q (new_AGEMA_signal_25705) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_9136), .Q (new_AGEMA_signal_25706) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_9137), .Q (new_AGEMA_signal_25707) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_9138), .Q (new_AGEMA_signal_25708) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M21), .Q (new_AGEMA_signal_25709) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_8623), .Q (new_AGEMA_signal_25710) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_8624), .Q (new_AGEMA_signal_25711) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_8625), .Q (new_AGEMA_signal_25712) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M23), .Q (new_AGEMA_signal_25713) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_8857), .Q (new_AGEMA_signal_25714) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_8858), .Q (new_AGEMA_signal_25715) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_8859), .Q (new_AGEMA_signal_25716) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M27), .Q (new_AGEMA_signal_25717) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_8863), .Q (new_AGEMA_signal_25718) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_8864), .Q (new_AGEMA_signal_25719) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_8865), .Q (new_AGEMA_signal_25720) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M24), .Q (new_AGEMA_signal_25721) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_9151), .Q (new_AGEMA_signal_25722) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_9152), .Q (new_AGEMA_signal_25723) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_9153), .Q (new_AGEMA_signal_25724) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M21), .Q (new_AGEMA_signal_25725) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_8635), .Q (new_AGEMA_signal_25726) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_8636), .Q (new_AGEMA_signal_25727) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_8637), .Q (new_AGEMA_signal_25728) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M23), .Q (new_AGEMA_signal_25729) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_8869), .Q (new_AGEMA_signal_25730) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_8870), .Q (new_AGEMA_signal_25731) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_8871), .Q (new_AGEMA_signal_25732) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M27), .Q (new_AGEMA_signal_25733) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_8875), .Q (new_AGEMA_signal_25734) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_8876), .Q (new_AGEMA_signal_25735) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_8877), .Q (new_AGEMA_signal_25736) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M24), .Q (new_AGEMA_signal_25737) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_9166), .Q (new_AGEMA_signal_25738) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_9167), .Q (new_AGEMA_signal_25739) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_9168), .Q (new_AGEMA_signal_25740) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_25741) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_8407), .Q (new_AGEMA_signal_25742) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_8408), .Q (new_AGEMA_signal_25743) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_8409), .Q (new_AGEMA_signal_25744) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_25745) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_8641), .Q (new_AGEMA_signal_25746) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_8642), .Q (new_AGEMA_signal_25747) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_8643), .Q (new_AGEMA_signal_25748) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_25749) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_8647), .Q (new_AGEMA_signal_25750) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_8648), .Q (new_AGEMA_signal_25751) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_8649), .Q (new_AGEMA_signal_25752) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_25753) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_8881), .Q (new_AGEMA_signal_25754) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_8882), .Q (new_AGEMA_signal_25755) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_8883), .Q (new_AGEMA_signal_25756) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_25757) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_8419), .Q (new_AGEMA_signal_25758) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_8420), .Q (new_AGEMA_signal_25759) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_8421), .Q (new_AGEMA_signal_25760) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_25761) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_8653), .Q (new_AGEMA_signal_25762) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_8654), .Q (new_AGEMA_signal_25763) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_8655), .Q (new_AGEMA_signal_25764) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_25765) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_8659), .Q (new_AGEMA_signal_25766) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_8660), .Q (new_AGEMA_signal_25767) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_8661), .Q (new_AGEMA_signal_25768) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_25769) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_8896), .Q (new_AGEMA_signal_25770) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_8897), .Q (new_AGEMA_signal_25771) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_8898), .Q (new_AGEMA_signal_25772) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_25773) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_8431), .Q (new_AGEMA_signal_25774) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_8432), .Q (new_AGEMA_signal_25775) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_8433), .Q (new_AGEMA_signal_25776) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_25777) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_8665), .Q (new_AGEMA_signal_25778) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_8666), .Q (new_AGEMA_signal_25779) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_8667), .Q (new_AGEMA_signal_25780) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_25781) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_8671), .Q (new_AGEMA_signal_25782) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_8672), .Q (new_AGEMA_signal_25783) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_8673), .Q (new_AGEMA_signal_25784) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_25785) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_8911), .Q (new_AGEMA_signal_25786) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_8912), .Q (new_AGEMA_signal_25787) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_8913), .Q (new_AGEMA_signal_25788) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_25789) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_8443), .Q (new_AGEMA_signal_25790) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_8444), .Q (new_AGEMA_signal_25791) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_8445), .Q (new_AGEMA_signal_25792) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_25793) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_8677), .Q (new_AGEMA_signal_25794) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_8678), .Q (new_AGEMA_signal_25795) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_8679), .Q (new_AGEMA_signal_25796) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_25797) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_8683), .Q (new_AGEMA_signal_25798) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_8684), .Q (new_AGEMA_signal_25799) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_8685), .Q (new_AGEMA_signal_25800) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_25801) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_8926), .Q (new_AGEMA_signal_25802) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_8927), .Q (new_AGEMA_signal_25803) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_8928), .Q (new_AGEMA_signal_25804) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_26125), .Q (new_AGEMA_signal_26126) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_26129), .Q (new_AGEMA_signal_26130) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_26133), .Q (new_AGEMA_signal_26134) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_26137), .Q (new_AGEMA_signal_26138) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_26141), .Q (new_AGEMA_signal_26142) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_26145), .Q (new_AGEMA_signal_26146) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_26149), .Q (new_AGEMA_signal_26150) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_26153), .Q (new_AGEMA_signal_26154) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_26157), .Q (new_AGEMA_signal_26158) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_26161), .Q (new_AGEMA_signal_26162) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_26165), .Q (new_AGEMA_signal_26166) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_26169), .Q (new_AGEMA_signal_26170) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_26173), .Q (new_AGEMA_signal_26174) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_26177), .Q (new_AGEMA_signal_26178) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_26181), .Q (new_AGEMA_signal_26182) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_26185), .Q (new_AGEMA_signal_26186) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_26189), .Q (new_AGEMA_signal_26190) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_26193), .Q (new_AGEMA_signal_26194) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_26197), .Q (new_AGEMA_signal_26198) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_26201), .Q (new_AGEMA_signal_26202) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_26205), .Q (new_AGEMA_signal_26206) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_26209), .Q (new_AGEMA_signal_26210) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_26213), .Q (new_AGEMA_signal_26214) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_26217), .Q (new_AGEMA_signal_26218) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_26221), .Q (new_AGEMA_signal_26222) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_26225), .Q (new_AGEMA_signal_26226) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_26229), .Q (new_AGEMA_signal_26230) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_26233), .Q (new_AGEMA_signal_26234) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_26237), .Q (new_AGEMA_signal_26238) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_26241), .Q (new_AGEMA_signal_26242) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_26245), .Q (new_AGEMA_signal_26246) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_26249), .Q (new_AGEMA_signal_26250) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_26253), .Q (new_AGEMA_signal_26254) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_26257), .Q (new_AGEMA_signal_26258) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_26261), .Q (new_AGEMA_signal_26262) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_26265), .Q (new_AGEMA_signal_26266) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_26269), .Q (new_AGEMA_signal_26270) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_26273), .Q (new_AGEMA_signal_26274) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_26277), .Q (new_AGEMA_signal_26278) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_26281), .Q (new_AGEMA_signal_26282) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_26285), .Q (new_AGEMA_signal_26286) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_26289), .Q (new_AGEMA_signal_26290) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_26293), .Q (new_AGEMA_signal_26294) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_26297), .Q (new_AGEMA_signal_26298) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_26301), .Q (new_AGEMA_signal_26302) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_26305), .Q (new_AGEMA_signal_26306) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_26309), .Q (new_AGEMA_signal_26310) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_26313), .Q (new_AGEMA_signal_26314) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_26317), .Q (new_AGEMA_signal_26318) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_26321), .Q (new_AGEMA_signal_26322) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_26325), .Q (new_AGEMA_signal_26326) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_26329), .Q (new_AGEMA_signal_26330) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_26333), .Q (new_AGEMA_signal_26334) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_26337), .Q (new_AGEMA_signal_26338) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_26341), .Q (new_AGEMA_signal_26342) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_26345), .Q (new_AGEMA_signal_26346) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_26349), .Q (new_AGEMA_signal_26350) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_26353), .Q (new_AGEMA_signal_26354) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_26357), .Q (new_AGEMA_signal_26358) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_26361), .Q (new_AGEMA_signal_26362) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_26365), .Q (new_AGEMA_signal_26366) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_26369), .Q (new_AGEMA_signal_26370) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_26373), .Q (new_AGEMA_signal_26374) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_26377), .Q (new_AGEMA_signal_26378) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_26381), .Q (new_AGEMA_signal_26382) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_26385), .Q (new_AGEMA_signal_26386) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_26389), .Q (new_AGEMA_signal_26390) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_26393), .Q (new_AGEMA_signal_26394) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_26397), .Q (new_AGEMA_signal_26398) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_26401), .Q (new_AGEMA_signal_26402) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_26405), .Q (new_AGEMA_signal_26406) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_26409), .Q (new_AGEMA_signal_26410) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_26413), .Q (new_AGEMA_signal_26414) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_26417), .Q (new_AGEMA_signal_26418) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_26421), .Q (new_AGEMA_signal_26422) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_26425), .Q (new_AGEMA_signal_26426) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_26429), .Q (new_AGEMA_signal_26430) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_26433), .Q (new_AGEMA_signal_26434) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_26437), .Q (new_AGEMA_signal_26438) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_26441), .Q (new_AGEMA_signal_26442) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_26445), .Q (new_AGEMA_signal_26446) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_26449), .Q (new_AGEMA_signal_26450) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_26453), .Q (new_AGEMA_signal_26454) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_26457), .Q (new_AGEMA_signal_26458) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_26461), .Q (new_AGEMA_signal_26462) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_26465), .Q (new_AGEMA_signal_26466) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_26469), .Q (new_AGEMA_signal_26470) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_26473), .Q (new_AGEMA_signal_26474) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_26477), .Q (new_AGEMA_signal_26478) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_26481), .Q (new_AGEMA_signal_26482) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_26485), .Q (new_AGEMA_signal_26486) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_26489), .Q (new_AGEMA_signal_26490) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_26493), .Q (new_AGEMA_signal_26494) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_26497), .Q (new_AGEMA_signal_26498) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_26501), .Q (new_AGEMA_signal_26502) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_26505), .Q (new_AGEMA_signal_26506) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_26509), .Q (new_AGEMA_signal_26510) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_26513), .Q (new_AGEMA_signal_26514) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_26517), .Q (new_AGEMA_signal_26518) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_26521), .Q (new_AGEMA_signal_26522) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_26525), .Q (new_AGEMA_signal_26526) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_26529), .Q (new_AGEMA_signal_26530) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_26533), .Q (new_AGEMA_signal_26534) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_26537), .Q (new_AGEMA_signal_26538) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_26541), .Q (new_AGEMA_signal_26542) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_26545), .Q (new_AGEMA_signal_26546) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_26549), .Q (new_AGEMA_signal_26550) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_26553), .Q (new_AGEMA_signal_26554) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_26557), .Q (new_AGEMA_signal_26558) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_26561), .Q (new_AGEMA_signal_26562) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_26565), .Q (new_AGEMA_signal_26566) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_26569), .Q (new_AGEMA_signal_26570) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_26573), .Q (new_AGEMA_signal_26574) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_26577), .Q (new_AGEMA_signal_26578) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_26581), .Q (new_AGEMA_signal_26582) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_26585), .Q (new_AGEMA_signal_26586) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_26589), .Q (new_AGEMA_signal_26590) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_26593), .Q (new_AGEMA_signal_26594) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_26597), .Q (new_AGEMA_signal_26598) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_26601), .Q (new_AGEMA_signal_26602) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_26605), .Q (new_AGEMA_signal_26606) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_26609), .Q (new_AGEMA_signal_26610) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_26613), .Q (new_AGEMA_signal_26614) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_26617), .Q (new_AGEMA_signal_26618) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_26621), .Q (new_AGEMA_signal_26622) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_26625), .Q (new_AGEMA_signal_26626) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_26629), .Q (new_AGEMA_signal_26630) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_26633), .Q (new_AGEMA_signal_26634) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_26637), .Q (new_AGEMA_signal_26638) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_26641), .Q (new_AGEMA_signal_26642) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_26645), .Q (new_AGEMA_signal_26646) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_26649), .Q (new_AGEMA_signal_26650) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_26653), .Q (new_AGEMA_signal_26654) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_26657), .Q (new_AGEMA_signal_26658) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_26661), .Q (new_AGEMA_signal_26662) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_26665), .Q (new_AGEMA_signal_26666) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_26669), .Q (new_AGEMA_signal_26670) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_26673), .Q (new_AGEMA_signal_26674) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_26677), .Q (new_AGEMA_signal_26678) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_26681), .Q (new_AGEMA_signal_26682) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_26685), .Q (new_AGEMA_signal_26686) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_26689), .Q (new_AGEMA_signal_26690) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_26693), .Q (new_AGEMA_signal_26694) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_26697), .Q (new_AGEMA_signal_26698) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_26701), .Q (new_AGEMA_signal_26702) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_26705), .Q (new_AGEMA_signal_26706) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_26709), .Q (new_AGEMA_signal_26710) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_26713), .Q (new_AGEMA_signal_26714) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_26717), .Q (new_AGEMA_signal_26718) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_26721), .Q (new_AGEMA_signal_26722) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_26725), .Q (new_AGEMA_signal_26726) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_26729), .Q (new_AGEMA_signal_26730) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_26733), .Q (new_AGEMA_signal_26734) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_26737), .Q (new_AGEMA_signal_26738) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_26741), .Q (new_AGEMA_signal_26742) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_26745), .Q (new_AGEMA_signal_26746) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_26749), .Q (new_AGEMA_signal_26750) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_26753), .Q (new_AGEMA_signal_26754) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_26757), .Q (new_AGEMA_signal_26758) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_26761), .Q (new_AGEMA_signal_26762) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_26765), .Q (new_AGEMA_signal_26766) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_26769), .Q (new_AGEMA_signal_26770) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_26773), .Q (new_AGEMA_signal_26774) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_26777), .Q (new_AGEMA_signal_26778) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_26781), .Q (new_AGEMA_signal_26782) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_26785), .Q (new_AGEMA_signal_26786) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_26789), .Q (new_AGEMA_signal_26790) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_26793), .Q (new_AGEMA_signal_26794) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_26797), .Q (new_AGEMA_signal_26798) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_26801), .Q (new_AGEMA_signal_26802) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_26805), .Q (new_AGEMA_signal_26806) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_26809), .Q (new_AGEMA_signal_26810) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_26813), .Q (new_AGEMA_signal_26814) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_26817), .Q (new_AGEMA_signal_26818) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_26821), .Q (new_AGEMA_signal_26822) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_26825), .Q (new_AGEMA_signal_26826) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_26829), .Q (new_AGEMA_signal_26830) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_26833), .Q (new_AGEMA_signal_26834) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_26837), .Q (new_AGEMA_signal_26838) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_26841), .Q (new_AGEMA_signal_26842) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_26845), .Q (new_AGEMA_signal_26846) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_26849), .Q (new_AGEMA_signal_26850) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_26853), .Q (new_AGEMA_signal_26854) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_26857), .Q (new_AGEMA_signal_26858) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_26861), .Q (new_AGEMA_signal_26862) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_26865), .Q (new_AGEMA_signal_26866) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_26869), .Q (new_AGEMA_signal_26870) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_26873), .Q (new_AGEMA_signal_26874) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_26877), .Q (new_AGEMA_signal_26878) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_26881), .Q (new_AGEMA_signal_26882) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_26885), .Q (new_AGEMA_signal_26886) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_26889), .Q (new_AGEMA_signal_26890) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_26893), .Q (new_AGEMA_signal_26894) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_26897), .Q (new_AGEMA_signal_26898) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_26901), .Q (new_AGEMA_signal_26902) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_26905), .Q (new_AGEMA_signal_26906) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_26909), .Q (new_AGEMA_signal_26910) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_26913), .Q (new_AGEMA_signal_26914) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_26917), .Q (new_AGEMA_signal_26918) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_26921), .Q (new_AGEMA_signal_26922) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_26925), .Q (new_AGEMA_signal_26926) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_26929), .Q (new_AGEMA_signal_26930) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_26933), .Q (new_AGEMA_signal_26934) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_26937), .Q (new_AGEMA_signal_26938) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_26941), .Q (new_AGEMA_signal_26942) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_26945), .Q (new_AGEMA_signal_26946) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_26949), .Q (new_AGEMA_signal_26950) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_26953), .Q (new_AGEMA_signal_26954) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_26957), .Q (new_AGEMA_signal_26958) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_26961), .Q (new_AGEMA_signal_26962) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_26965), .Q (new_AGEMA_signal_26966) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_26969), .Q (new_AGEMA_signal_26970) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_26973), .Q (new_AGEMA_signal_26974) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_26977), .Q (new_AGEMA_signal_26978) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_26981), .Q (new_AGEMA_signal_26982) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_26985), .Q (new_AGEMA_signal_26986) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_26989), .Q (new_AGEMA_signal_26990) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_26993), .Q (new_AGEMA_signal_26994) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_26997), .Q (new_AGEMA_signal_26998) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_27001), .Q (new_AGEMA_signal_27002) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_27005), .Q (new_AGEMA_signal_27006) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_27009), .Q (new_AGEMA_signal_27010) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_27013), .Q (new_AGEMA_signal_27014) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_27017), .Q (new_AGEMA_signal_27018) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_27021), .Q (new_AGEMA_signal_27022) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_27025), .Q (new_AGEMA_signal_27026) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_27029), .Q (new_AGEMA_signal_27030) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_27033), .Q (new_AGEMA_signal_27034) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_27037), .Q (new_AGEMA_signal_27038) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_27041), .Q (new_AGEMA_signal_27042) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_27045), .Q (new_AGEMA_signal_27046) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_27049), .Q (new_AGEMA_signal_27050) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_27053), .Q (new_AGEMA_signal_27054) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_27057), .Q (new_AGEMA_signal_27058) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_27061), .Q (new_AGEMA_signal_27062) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_27065), .Q (new_AGEMA_signal_27066) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_27069), .Q (new_AGEMA_signal_27070) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_27073), .Q (new_AGEMA_signal_27074) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_27077), .Q (new_AGEMA_signal_27078) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_27081), .Q (new_AGEMA_signal_27082) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_27085), .Q (new_AGEMA_signal_27086) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_27089), .Q (new_AGEMA_signal_27090) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_27093), .Q (new_AGEMA_signal_27094) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_27097), .Q (new_AGEMA_signal_27098) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_27101), .Q (new_AGEMA_signal_27102) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_27105), .Q (new_AGEMA_signal_27106) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_27109), .Q (new_AGEMA_signal_27110) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_27113), .Q (new_AGEMA_signal_27114) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_27117), .Q (new_AGEMA_signal_27118) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_27121), .Q (new_AGEMA_signal_27122) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_27125), .Q (new_AGEMA_signal_27126) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_27129), .Q (new_AGEMA_signal_27130) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_27133), .Q (new_AGEMA_signal_27134) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_27137), .Q (new_AGEMA_signal_27138) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_27141), .Q (new_AGEMA_signal_27142) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_27145), .Q (new_AGEMA_signal_27146) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_27149), .Q (new_AGEMA_signal_27150) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_27153), .Q (new_AGEMA_signal_27154) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_27157), .Q (new_AGEMA_signal_27158) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_27161), .Q (new_AGEMA_signal_27162) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_27165), .Q (new_AGEMA_signal_27166) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_27169), .Q (new_AGEMA_signal_27170) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_27173), .Q (new_AGEMA_signal_27174) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_27177), .Q (new_AGEMA_signal_27178) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_27181), .Q (new_AGEMA_signal_27182) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_27185), .Q (new_AGEMA_signal_27186) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_27189), .Q (new_AGEMA_signal_27190) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_27193), .Q (new_AGEMA_signal_27194) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_27197), .Q (new_AGEMA_signal_27198) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_27201), .Q (new_AGEMA_signal_27202) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_27205), .Q (new_AGEMA_signal_27206) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_27209), .Q (new_AGEMA_signal_27210) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_27213), .Q (new_AGEMA_signal_27214) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_27217), .Q (new_AGEMA_signal_27218) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_27221), .Q (new_AGEMA_signal_27222) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_27225), .Q (new_AGEMA_signal_27226) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_27229), .Q (new_AGEMA_signal_27230) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_27233), .Q (new_AGEMA_signal_27234) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_27237), .Q (new_AGEMA_signal_27238) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_27241), .Q (new_AGEMA_signal_27242) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_27245), .Q (new_AGEMA_signal_27246) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_27249), .Q (new_AGEMA_signal_27250) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_27253), .Q (new_AGEMA_signal_27254) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_27257), .Q (new_AGEMA_signal_27258) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_27261), .Q (new_AGEMA_signal_27262) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_27265), .Q (new_AGEMA_signal_27266) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_27269), .Q (new_AGEMA_signal_27270) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_27273), .Q (new_AGEMA_signal_27274) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_27277), .Q (new_AGEMA_signal_27278) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_27281), .Q (new_AGEMA_signal_27282) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_27285), .Q (new_AGEMA_signal_27286) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_27289), .Q (new_AGEMA_signal_27290) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_27293), .Q (new_AGEMA_signal_27294) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_27297), .Q (new_AGEMA_signal_27298) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_27301), .Q (new_AGEMA_signal_27302) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_27305), .Q (new_AGEMA_signal_27306) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_27309), .Q (new_AGEMA_signal_27310) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_27313), .Q (new_AGEMA_signal_27314) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_27317), .Q (new_AGEMA_signal_27318) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_27321), .Q (new_AGEMA_signal_27322) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_27325), .Q (new_AGEMA_signal_27326) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_27329), .Q (new_AGEMA_signal_27330) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_27333), .Q (new_AGEMA_signal_27334) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_27337), .Q (new_AGEMA_signal_27338) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_27341), .Q (new_AGEMA_signal_27342) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_27345), .Q (new_AGEMA_signal_27346) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_27349), .Q (new_AGEMA_signal_27350) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_27353), .Q (new_AGEMA_signal_27354) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_27357), .Q (new_AGEMA_signal_27358) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_27361), .Q (new_AGEMA_signal_27362) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_27365), .Q (new_AGEMA_signal_27366) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_27369), .Q (new_AGEMA_signal_27370) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_27373), .Q (new_AGEMA_signal_27374) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_27377), .Q (new_AGEMA_signal_27378) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_27381), .Q (new_AGEMA_signal_27382) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_27385), .Q (new_AGEMA_signal_27386) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_27389), .Q (new_AGEMA_signal_27390) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_27393), .Q (new_AGEMA_signal_27394) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_27397), .Q (new_AGEMA_signal_27398) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_27401), .Q (new_AGEMA_signal_27402) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_27405), .Q (new_AGEMA_signal_27406) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_27409), .Q (new_AGEMA_signal_27410) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_27413), .Q (new_AGEMA_signal_27414) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_27417), .Q (new_AGEMA_signal_27418) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_27421), .Q (new_AGEMA_signal_27422) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_27425), .Q (new_AGEMA_signal_27426) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_27429), .Q (new_AGEMA_signal_27430) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_27433), .Q (new_AGEMA_signal_27434) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_27437), .Q (new_AGEMA_signal_27438) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_27441), .Q (new_AGEMA_signal_27442) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_27445), .Q (new_AGEMA_signal_27446) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_27449), .Q (new_AGEMA_signal_27450) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_27453), .Q (new_AGEMA_signal_27454) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_27457), .Q (new_AGEMA_signal_27458) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C (clk), .D (new_AGEMA_signal_27461), .Q (new_AGEMA_signal_27462) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_27465), .Q (new_AGEMA_signal_27466) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_27469), .Q (new_AGEMA_signal_27470) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C (clk), .D (new_AGEMA_signal_27473), .Q (new_AGEMA_signal_27474) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_27477), .Q (new_AGEMA_signal_27478) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_27481), .Q (new_AGEMA_signal_27482) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_27485), .Q (new_AGEMA_signal_27486) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_27489), .Q (new_AGEMA_signal_27490) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_27493), .Q (new_AGEMA_signal_27494) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C (clk), .D (new_AGEMA_signal_27497), .Q (new_AGEMA_signal_27498) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_27501), .Q (new_AGEMA_signal_27502) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_27505), .Q (new_AGEMA_signal_27506) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_27509), .Q (new_AGEMA_signal_27510) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_27513), .Q (new_AGEMA_signal_27514) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_27517), .Q (new_AGEMA_signal_27518) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_27521), .Q (new_AGEMA_signal_27522) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_27525), .Q (new_AGEMA_signal_27526) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_27529), .Q (new_AGEMA_signal_27530) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C (clk), .D (new_AGEMA_signal_27533), .Q (new_AGEMA_signal_27534) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_27537), .Q (new_AGEMA_signal_27538) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_27541), .Q (new_AGEMA_signal_27542) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_27545), .Q (new_AGEMA_signal_27546) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_27549), .Q (new_AGEMA_signal_27550) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_27553), .Q (new_AGEMA_signal_27554) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_27557), .Q (new_AGEMA_signal_27558) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_27561), .Q (new_AGEMA_signal_27562) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_27565), .Q (new_AGEMA_signal_27566) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C (clk), .D (new_AGEMA_signal_27569), .Q (new_AGEMA_signal_27570) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_27573), .Q (new_AGEMA_signal_27574) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_27577), .Q (new_AGEMA_signal_27578) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_27581), .Q (new_AGEMA_signal_27582) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_27585), .Q (new_AGEMA_signal_27586) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_27589), .Q (new_AGEMA_signal_27590) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_27593), .Q (new_AGEMA_signal_27594) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_27597), .Q (new_AGEMA_signal_27598) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_27601), .Q (new_AGEMA_signal_27602) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C (clk), .D (new_AGEMA_signal_27605), .Q (new_AGEMA_signal_27606) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_27609), .Q (new_AGEMA_signal_27610) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_27613), .Q (new_AGEMA_signal_27614) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_27617), .Q (new_AGEMA_signal_27618) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_27621), .Q (new_AGEMA_signal_27622) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_27625), .Q (new_AGEMA_signal_27626) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_27629), .Q (new_AGEMA_signal_27630) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_27633), .Q (new_AGEMA_signal_27634) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_27637), .Q (new_AGEMA_signal_27638) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C (clk), .D (new_AGEMA_signal_27641), .Q (new_AGEMA_signal_27642) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C (clk), .D (new_AGEMA_signal_27645), .Q (new_AGEMA_signal_27646) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C (clk), .D (new_AGEMA_signal_27649), .Q (new_AGEMA_signal_27650) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C (clk), .D (new_AGEMA_signal_27653), .Q (new_AGEMA_signal_27654) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C (clk), .D (new_AGEMA_signal_27657), .Q (new_AGEMA_signal_27658) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C (clk), .D (new_AGEMA_signal_27661), .Q (new_AGEMA_signal_27662) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C (clk), .D (new_AGEMA_signal_27665), .Q (new_AGEMA_signal_27666) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C (clk), .D (new_AGEMA_signal_27669), .Q (new_AGEMA_signal_27670) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C (clk), .D (new_AGEMA_signal_27673), .Q (new_AGEMA_signal_27674) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C (clk), .D (new_AGEMA_signal_27677), .Q (new_AGEMA_signal_27678) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C (clk), .D (new_AGEMA_signal_27681), .Q (new_AGEMA_signal_27682) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C (clk), .D (new_AGEMA_signal_27685), .Q (new_AGEMA_signal_27686) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C (clk), .D (new_AGEMA_signal_27689), .Q (new_AGEMA_signal_27690) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C (clk), .D (new_AGEMA_signal_27693), .Q (new_AGEMA_signal_27694) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C (clk), .D (new_AGEMA_signal_27697), .Q (new_AGEMA_signal_27698) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C (clk), .D (new_AGEMA_signal_27701), .Q (new_AGEMA_signal_27702) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C (clk), .D (new_AGEMA_signal_27705), .Q (new_AGEMA_signal_27706) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C (clk), .D (new_AGEMA_signal_27709), .Q (new_AGEMA_signal_27710) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C (clk), .D (new_AGEMA_signal_27713), .Q (new_AGEMA_signal_27714) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C (clk), .D (new_AGEMA_signal_27717), .Q (new_AGEMA_signal_27718) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C (clk), .D (new_AGEMA_signal_27721), .Q (new_AGEMA_signal_27722) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C (clk), .D (new_AGEMA_signal_27725), .Q (new_AGEMA_signal_27726) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C (clk), .D (new_AGEMA_signal_27729), .Q (new_AGEMA_signal_27730) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C (clk), .D (new_AGEMA_signal_27733), .Q (new_AGEMA_signal_27734) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C (clk), .D (new_AGEMA_signal_27737), .Q (new_AGEMA_signal_27738) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C (clk), .D (new_AGEMA_signal_27741), .Q (new_AGEMA_signal_27742) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C (clk), .D (new_AGEMA_signal_27745), .Q (new_AGEMA_signal_27746) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C (clk), .D (new_AGEMA_signal_27749), .Q (new_AGEMA_signal_27750) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C (clk), .D (new_AGEMA_signal_27753), .Q (new_AGEMA_signal_27754) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C (clk), .D (new_AGEMA_signal_27757), .Q (new_AGEMA_signal_27758) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C (clk), .D (new_AGEMA_signal_27761), .Q (new_AGEMA_signal_27762) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C (clk), .D (new_AGEMA_signal_27765), .Q (new_AGEMA_signal_27766) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C (clk), .D (new_AGEMA_signal_27769), .Q (new_AGEMA_signal_27770) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C (clk), .D (new_AGEMA_signal_27773), .Q (new_AGEMA_signal_27774) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C (clk), .D (new_AGEMA_signal_27777), .Q (new_AGEMA_signal_27778) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C (clk), .D (new_AGEMA_signal_27781), .Q (new_AGEMA_signal_27782) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C (clk), .D (new_AGEMA_signal_27785), .Q (new_AGEMA_signal_27786) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C (clk), .D (new_AGEMA_signal_27789), .Q (new_AGEMA_signal_27790) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C (clk), .D (new_AGEMA_signal_27793), .Q (new_AGEMA_signal_27794) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C (clk), .D (new_AGEMA_signal_27797), .Q (new_AGEMA_signal_27798) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C (clk), .D (new_AGEMA_signal_27801), .Q (new_AGEMA_signal_27802) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C (clk), .D (new_AGEMA_signal_27805), .Q (new_AGEMA_signal_27806) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C (clk), .D (new_AGEMA_signal_27809), .Q (new_AGEMA_signal_27810) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C (clk), .D (new_AGEMA_signal_27813), .Q (new_AGEMA_signal_27814) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C (clk), .D (new_AGEMA_signal_27817), .Q (new_AGEMA_signal_27818) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C (clk), .D (new_AGEMA_signal_27821), .Q (new_AGEMA_signal_27822) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C (clk), .D (new_AGEMA_signal_27825), .Q (new_AGEMA_signal_27826) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C (clk), .D (new_AGEMA_signal_27829), .Q (new_AGEMA_signal_27830) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C (clk), .D (new_AGEMA_signal_27833), .Q (new_AGEMA_signal_27834) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C (clk), .D (new_AGEMA_signal_27837), .Q (new_AGEMA_signal_27838) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C (clk), .D (new_AGEMA_signal_27841), .Q (new_AGEMA_signal_27842) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C (clk), .D (new_AGEMA_signal_27845), .Q (new_AGEMA_signal_27846) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C (clk), .D (new_AGEMA_signal_27849), .Q (new_AGEMA_signal_27850) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C (clk), .D (new_AGEMA_signal_27853), .Q (new_AGEMA_signal_27854) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C (clk), .D (new_AGEMA_signal_27857), .Q (new_AGEMA_signal_27858) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C (clk), .D (new_AGEMA_signal_27861), .Q (new_AGEMA_signal_27862) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C (clk), .D (new_AGEMA_signal_27865), .Q (new_AGEMA_signal_27866) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C (clk), .D (new_AGEMA_signal_27869), .Q (new_AGEMA_signal_27870) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C (clk), .D (new_AGEMA_signal_27873), .Q (new_AGEMA_signal_27874) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C (clk), .D (new_AGEMA_signal_27877), .Q (new_AGEMA_signal_27878) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C (clk), .D (new_AGEMA_signal_27881), .Q (new_AGEMA_signal_27882) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C (clk), .D (new_AGEMA_signal_27885), .Q (new_AGEMA_signal_27886) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C (clk), .D (new_AGEMA_signal_27889), .Q (new_AGEMA_signal_27890) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C (clk), .D (new_AGEMA_signal_27893), .Q (new_AGEMA_signal_27894) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C (clk), .D (new_AGEMA_signal_27897), .Q (new_AGEMA_signal_27898) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C (clk), .D (new_AGEMA_signal_27901), .Q (new_AGEMA_signal_27902) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C (clk), .D (new_AGEMA_signal_27905), .Q (new_AGEMA_signal_27906) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C (clk), .D (new_AGEMA_signal_27909), .Q (new_AGEMA_signal_27910) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C (clk), .D (new_AGEMA_signal_27913), .Q (new_AGEMA_signal_27914) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C (clk), .D (new_AGEMA_signal_27917), .Q (new_AGEMA_signal_27918) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C (clk), .D (new_AGEMA_signal_27921), .Q (new_AGEMA_signal_27922) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C (clk), .D (new_AGEMA_signal_27925), .Q (new_AGEMA_signal_27926) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C (clk), .D (new_AGEMA_signal_27929), .Q (new_AGEMA_signal_27930) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C (clk), .D (new_AGEMA_signal_27933), .Q (new_AGEMA_signal_27934) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C (clk), .D (new_AGEMA_signal_27937), .Q (new_AGEMA_signal_27938) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C (clk), .D (new_AGEMA_signal_27941), .Q (new_AGEMA_signal_27942) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C (clk), .D (new_AGEMA_signal_27945), .Q (new_AGEMA_signal_27946) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C (clk), .D (new_AGEMA_signal_27949), .Q (new_AGEMA_signal_27950) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C (clk), .D (new_AGEMA_signal_27953), .Q (new_AGEMA_signal_27954) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C (clk), .D (new_AGEMA_signal_27957), .Q (new_AGEMA_signal_27958) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C (clk), .D (new_AGEMA_signal_27961), .Q (new_AGEMA_signal_27962) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C (clk), .D (new_AGEMA_signal_27965), .Q (new_AGEMA_signal_27966) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C (clk), .D (new_AGEMA_signal_27969), .Q (new_AGEMA_signal_27970) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C (clk), .D (new_AGEMA_signal_27973), .Q (new_AGEMA_signal_27974) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C (clk), .D (new_AGEMA_signal_27977), .Q (new_AGEMA_signal_27978) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C (clk), .D (new_AGEMA_signal_27981), .Q (new_AGEMA_signal_27982) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C (clk), .D (new_AGEMA_signal_27985), .Q (new_AGEMA_signal_27986) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C (clk), .D (new_AGEMA_signal_27989), .Q (new_AGEMA_signal_27990) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C (clk), .D (new_AGEMA_signal_27993), .Q (new_AGEMA_signal_27994) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C (clk), .D (new_AGEMA_signal_27997), .Q (new_AGEMA_signal_27998) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C (clk), .D (new_AGEMA_signal_28001), .Q (new_AGEMA_signal_28002) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C (clk), .D (new_AGEMA_signal_28005), .Q (new_AGEMA_signal_28006) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C (clk), .D (new_AGEMA_signal_28009), .Q (new_AGEMA_signal_28010) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C (clk), .D (new_AGEMA_signal_28013), .Q (new_AGEMA_signal_28014) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C (clk), .D (new_AGEMA_signal_28017), .Q (new_AGEMA_signal_28018) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C (clk), .D (new_AGEMA_signal_28021), .Q (new_AGEMA_signal_28022) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C (clk), .D (new_AGEMA_signal_28025), .Q (new_AGEMA_signal_28026) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C (clk), .D (new_AGEMA_signal_28029), .Q (new_AGEMA_signal_28030) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C (clk), .D (new_AGEMA_signal_28033), .Q (new_AGEMA_signal_28034) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C (clk), .D (new_AGEMA_signal_28037), .Q (new_AGEMA_signal_28038) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C (clk), .D (new_AGEMA_signal_28041), .Q (new_AGEMA_signal_28042) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C (clk), .D (new_AGEMA_signal_28045), .Q (new_AGEMA_signal_28046) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C (clk), .D (new_AGEMA_signal_28049), .Q (new_AGEMA_signal_28050) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C (clk), .D (new_AGEMA_signal_28053), .Q (new_AGEMA_signal_28054) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C (clk), .D (new_AGEMA_signal_28057), .Q (new_AGEMA_signal_28058) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C (clk), .D (new_AGEMA_signal_28061), .Q (new_AGEMA_signal_28062) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C (clk), .D (new_AGEMA_signal_28065), .Q (new_AGEMA_signal_28066) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C (clk), .D (new_AGEMA_signal_28069), .Q (new_AGEMA_signal_28070) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C (clk), .D (new_AGEMA_signal_28073), .Q (new_AGEMA_signal_28074) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C (clk), .D (new_AGEMA_signal_28077), .Q (new_AGEMA_signal_28078) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C (clk), .D (new_AGEMA_signal_28081), .Q (new_AGEMA_signal_28082) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C (clk), .D (new_AGEMA_signal_28085), .Q (new_AGEMA_signal_28086) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C (clk), .D (new_AGEMA_signal_28089), .Q (new_AGEMA_signal_28090) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C (clk), .D (new_AGEMA_signal_28093), .Q (new_AGEMA_signal_28094) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C (clk), .D (new_AGEMA_signal_28097), .Q (new_AGEMA_signal_28098) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C (clk), .D (new_AGEMA_signal_28101), .Q (new_AGEMA_signal_28102) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C (clk), .D (new_AGEMA_signal_28105), .Q (new_AGEMA_signal_28106) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C (clk), .D (new_AGEMA_signal_28109), .Q (new_AGEMA_signal_28110) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C (clk), .D (new_AGEMA_signal_28113), .Q (new_AGEMA_signal_28114) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C (clk), .D (new_AGEMA_signal_28117), .Q (new_AGEMA_signal_28118) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C (clk), .D (new_AGEMA_signal_28121), .Q (new_AGEMA_signal_28122) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C (clk), .D (new_AGEMA_signal_28125), .Q (new_AGEMA_signal_28126) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C (clk), .D (new_AGEMA_signal_28129), .Q (new_AGEMA_signal_28130) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C (clk), .D (new_AGEMA_signal_28133), .Q (new_AGEMA_signal_28134) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C (clk), .D (new_AGEMA_signal_28137), .Q (new_AGEMA_signal_28138) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C (clk), .D (new_AGEMA_signal_28141), .Q (new_AGEMA_signal_28142) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C (clk), .D (new_AGEMA_signal_28145), .Q (new_AGEMA_signal_28146) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C (clk), .D (new_AGEMA_signal_28149), .Q (new_AGEMA_signal_28150) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C (clk), .D (new_AGEMA_signal_28153), .Q (new_AGEMA_signal_28154) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C (clk), .D (new_AGEMA_signal_28157), .Q (new_AGEMA_signal_28158) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C (clk), .D (new_AGEMA_signal_28161), .Q (new_AGEMA_signal_28162) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C (clk), .D (new_AGEMA_signal_28165), .Q (new_AGEMA_signal_28166) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C (clk), .D (new_AGEMA_signal_28169), .Q (new_AGEMA_signal_28170) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C (clk), .D (new_AGEMA_signal_28173), .Q (new_AGEMA_signal_28174) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C (clk), .D (new_AGEMA_signal_28177), .Q (new_AGEMA_signal_28178) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C (clk), .D (new_AGEMA_signal_28181), .Q (new_AGEMA_signal_28182) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C (clk), .D (new_AGEMA_signal_28185), .Q (new_AGEMA_signal_28186) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C (clk), .D (new_AGEMA_signal_28189), .Q (new_AGEMA_signal_28190) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C (clk), .D (new_AGEMA_signal_28193), .Q (new_AGEMA_signal_28194) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C (clk), .D (new_AGEMA_signal_28197), .Q (new_AGEMA_signal_28198) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C (clk), .D (new_AGEMA_signal_28201), .Q (new_AGEMA_signal_28202) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C (clk), .D (new_AGEMA_signal_28205), .Q (new_AGEMA_signal_28206) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C (clk), .D (new_AGEMA_signal_28208), .Q (new_AGEMA_signal_28209) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C (clk), .D (new_AGEMA_signal_28211), .Q (new_AGEMA_signal_28212) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C (clk), .D (new_AGEMA_signal_28214), .Q (new_AGEMA_signal_28215) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C (clk), .D (new_AGEMA_signal_28217), .Q (new_AGEMA_signal_28218) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C (clk), .D (new_AGEMA_signal_28220), .Q (new_AGEMA_signal_28221) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C (clk), .D (new_AGEMA_signal_28223), .Q (new_AGEMA_signal_28224) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C (clk), .D (new_AGEMA_signal_28226), .Q (new_AGEMA_signal_28227) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C (clk), .D (new_AGEMA_signal_28229), .Q (new_AGEMA_signal_28230) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C (clk), .D (new_AGEMA_signal_28232), .Q (new_AGEMA_signal_28233) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C (clk), .D (new_AGEMA_signal_28235), .Q (new_AGEMA_signal_28236) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C (clk), .D (new_AGEMA_signal_28238), .Q (new_AGEMA_signal_28239) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C (clk), .D (new_AGEMA_signal_28241), .Q (new_AGEMA_signal_28242) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C (clk), .D (new_AGEMA_signal_28244), .Q (new_AGEMA_signal_28245) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C (clk), .D (new_AGEMA_signal_28247), .Q (new_AGEMA_signal_28248) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C (clk), .D (new_AGEMA_signal_28250), .Q (new_AGEMA_signal_28251) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C (clk), .D (new_AGEMA_signal_28253), .Q (new_AGEMA_signal_28254) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C (clk), .D (new_AGEMA_signal_28256), .Q (new_AGEMA_signal_28257) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C (clk), .D (new_AGEMA_signal_28259), .Q (new_AGEMA_signal_28260) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C (clk), .D (new_AGEMA_signal_28262), .Q (new_AGEMA_signal_28263) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C (clk), .D (new_AGEMA_signal_28265), .Q (new_AGEMA_signal_28266) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C (clk), .D (new_AGEMA_signal_28268), .Q (new_AGEMA_signal_28269) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C (clk), .D (new_AGEMA_signal_28271), .Q (new_AGEMA_signal_28272) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C (clk), .D (new_AGEMA_signal_28274), .Q (new_AGEMA_signal_28275) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C (clk), .D (new_AGEMA_signal_28277), .Q (new_AGEMA_signal_28278) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C (clk), .D (new_AGEMA_signal_28280), .Q (new_AGEMA_signal_28281) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C (clk), .D (new_AGEMA_signal_28283), .Q (new_AGEMA_signal_28284) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C (clk), .D (new_AGEMA_signal_28286), .Q (new_AGEMA_signal_28287) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C (clk), .D (new_AGEMA_signal_28289), .Q (new_AGEMA_signal_28290) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C (clk), .D (new_AGEMA_signal_28292), .Q (new_AGEMA_signal_28293) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C (clk), .D (new_AGEMA_signal_28295), .Q (new_AGEMA_signal_28296) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C (clk), .D (new_AGEMA_signal_28298), .Q (new_AGEMA_signal_28299) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C (clk), .D (new_AGEMA_signal_28301), .Q (new_AGEMA_signal_28302) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C (clk), .D (new_AGEMA_signal_28304), .Q (new_AGEMA_signal_28305) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C (clk), .D (new_AGEMA_signal_28307), .Q (new_AGEMA_signal_28308) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C (clk), .D (new_AGEMA_signal_28310), .Q (new_AGEMA_signal_28311) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C (clk), .D (new_AGEMA_signal_28313), .Q (new_AGEMA_signal_28314) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C (clk), .D (new_AGEMA_signal_28316), .Q (new_AGEMA_signal_28317) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C (clk), .D (new_AGEMA_signal_28319), .Q (new_AGEMA_signal_28320) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C (clk), .D (new_AGEMA_signal_28322), .Q (new_AGEMA_signal_28323) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C (clk), .D (new_AGEMA_signal_28325), .Q (new_AGEMA_signal_28326) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C (clk), .D (new_AGEMA_signal_28328), .Q (new_AGEMA_signal_28329) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C (clk), .D (new_AGEMA_signal_28331), .Q (new_AGEMA_signal_28332) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C (clk), .D (new_AGEMA_signal_28334), .Q (new_AGEMA_signal_28335) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C (clk), .D (new_AGEMA_signal_28337), .Q (new_AGEMA_signal_28338) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C (clk), .D (new_AGEMA_signal_28340), .Q (new_AGEMA_signal_28341) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C (clk), .D (new_AGEMA_signal_28343), .Q (new_AGEMA_signal_28344) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C (clk), .D (new_AGEMA_signal_28346), .Q (new_AGEMA_signal_28347) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C (clk), .D (new_AGEMA_signal_28349), .Q (new_AGEMA_signal_28350) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C (clk), .D (new_AGEMA_signal_28352), .Q (new_AGEMA_signal_28353) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C (clk), .D (new_AGEMA_signal_28355), .Q (new_AGEMA_signal_28356) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C (clk), .D (new_AGEMA_signal_28358), .Q (new_AGEMA_signal_28359) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C (clk), .D (new_AGEMA_signal_28361), .Q (new_AGEMA_signal_28362) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C (clk), .D (new_AGEMA_signal_28364), .Q (new_AGEMA_signal_28365) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C (clk), .D (new_AGEMA_signal_28367), .Q (new_AGEMA_signal_28368) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C (clk), .D (new_AGEMA_signal_28370), .Q (new_AGEMA_signal_28371) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C (clk), .D (new_AGEMA_signal_28373), .Q (new_AGEMA_signal_28374) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C (clk), .D (new_AGEMA_signal_28376), .Q (new_AGEMA_signal_28377) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C (clk), .D (new_AGEMA_signal_28379), .Q (new_AGEMA_signal_28380) ) ;
    buf_clk new_AGEMA_reg_buffer_7427 ( .C (clk), .D (new_AGEMA_signal_28382), .Q (new_AGEMA_signal_28383) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C (clk), .D (new_AGEMA_signal_28385), .Q (new_AGEMA_signal_28386) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C (clk), .D (new_AGEMA_signal_28388), .Q (new_AGEMA_signal_28389) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C (clk), .D (new_AGEMA_signal_28391), .Q (new_AGEMA_signal_28392) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C (clk), .D (new_AGEMA_signal_28394), .Q (new_AGEMA_signal_28395) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C (clk), .D (new_AGEMA_signal_28397), .Q (new_AGEMA_signal_28398) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C (clk), .D (new_AGEMA_signal_28400), .Q (new_AGEMA_signal_28401) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C (clk), .D (new_AGEMA_signal_28403), .Q (new_AGEMA_signal_28404) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C (clk), .D (new_AGEMA_signal_28406), .Q (new_AGEMA_signal_28407) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C (clk), .D (new_AGEMA_signal_28409), .Q (new_AGEMA_signal_28410) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C (clk), .D (new_AGEMA_signal_28412), .Q (new_AGEMA_signal_28413) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C (clk), .D (new_AGEMA_signal_28415), .Q (new_AGEMA_signal_28416) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C (clk), .D (new_AGEMA_signal_28418), .Q (new_AGEMA_signal_28419) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C (clk), .D (new_AGEMA_signal_28421), .Q (new_AGEMA_signal_28422) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C (clk), .D (new_AGEMA_signal_28424), .Q (new_AGEMA_signal_28425) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C (clk), .D (new_AGEMA_signal_28427), .Q (new_AGEMA_signal_28428) ) ;
    buf_clk new_AGEMA_reg_buffer_7475 ( .C (clk), .D (new_AGEMA_signal_28430), .Q (new_AGEMA_signal_28431) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C (clk), .D (new_AGEMA_signal_28433), .Q (new_AGEMA_signal_28434) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C (clk), .D (new_AGEMA_signal_28436), .Q (new_AGEMA_signal_28437) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C (clk), .D (new_AGEMA_signal_28439), .Q (new_AGEMA_signal_28440) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C (clk), .D (new_AGEMA_signal_28442), .Q (new_AGEMA_signal_28443) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C (clk), .D (new_AGEMA_signal_28445), .Q (new_AGEMA_signal_28446) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C (clk), .D (new_AGEMA_signal_28448), .Q (new_AGEMA_signal_28449) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C (clk), .D (new_AGEMA_signal_28451), .Q (new_AGEMA_signal_28452) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C (clk), .D (new_AGEMA_signal_28454), .Q (new_AGEMA_signal_28455) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C (clk), .D (new_AGEMA_signal_28457), .Q (new_AGEMA_signal_28458) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C (clk), .D (new_AGEMA_signal_28460), .Q (new_AGEMA_signal_28461) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C (clk), .D (new_AGEMA_signal_28463), .Q (new_AGEMA_signal_28464) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C (clk), .D (new_AGEMA_signal_28466), .Q (new_AGEMA_signal_28467) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C (clk), .D (new_AGEMA_signal_28469), .Q (new_AGEMA_signal_28470) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C (clk), .D (new_AGEMA_signal_28472), .Q (new_AGEMA_signal_28473) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C (clk), .D (new_AGEMA_signal_28475), .Q (new_AGEMA_signal_28476) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C (clk), .D (new_AGEMA_signal_28478), .Q (new_AGEMA_signal_28479) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C (clk), .D (new_AGEMA_signal_28481), .Q (new_AGEMA_signal_28482) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C (clk), .D (new_AGEMA_signal_28484), .Q (new_AGEMA_signal_28485) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C (clk), .D (new_AGEMA_signal_28487), .Q (new_AGEMA_signal_28488) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C (clk), .D (new_AGEMA_signal_28490), .Q (new_AGEMA_signal_28491) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C (clk), .D (new_AGEMA_signal_28493), .Q (new_AGEMA_signal_28494) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C (clk), .D (new_AGEMA_signal_28496), .Q (new_AGEMA_signal_28497) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C (clk), .D (new_AGEMA_signal_28499), .Q (new_AGEMA_signal_28500) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C (clk), .D (new_AGEMA_signal_28502), .Q (new_AGEMA_signal_28503) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C (clk), .D (new_AGEMA_signal_28505), .Q (new_AGEMA_signal_28506) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C (clk), .D (new_AGEMA_signal_28508), .Q (new_AGEMA_signal_28509) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C (clk), .D (new_AGEMA_signal_28511), .Q (new_AGEMA_signal_28512) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C (clk), .D (new_AGEMA_signal_28514), .Q (new_AGEMA_signal_28515) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C (clk), .D (new_AGEMA_signal_28517), .Q (new_AGEMA_signal_28518) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C (clk), .D (new_AGEMA_signal_28520), .Q (new_AGEMA_signal_28521) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C (clk), .D (new_AGEMA_signal_28523), .Q (new_AGEMA_signal_28524) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C (clk), .D (new_AGEMA_signal_28526), .Q (new_AGEMA_signal_28527) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C (clk), .D (new_AGEMA_signal_28529), .Q (new_AGEMA_signal_28530) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C (clk), .D (new_AGEMA_signal_28532), .Q (new_AGEMA_signal_28533) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C (clk), .D (new_AGEMA_signal_28535), .Q (new_AGEMA_signal_28536) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C (clk), .D (new_AGEMA_signal_28538), .Q (new_AGEMA_signal_28539) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C (clk), .D (new_AGEMA_signal_28541), .Q (new_AGEMA_signal_28542) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C (clk), .D (new_AGEMA_signal_28544), .Q (new_AGEMA_signal_28545) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C (clk), .D (new_AGEMA_signal_28547), .Q (new_AGEMA_signal_28548) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C (clk), .D (new_AGEMA_signal_28550), .Q (new_AGEMA_signal_28551) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C (clk), .D (new_AGEMA_signal_28553), .Q (new_AGEMA_signal_28554) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C (clk), .D (new_AGEMA_signal_28556), .Q (new_AGEMA_signal_28557) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C (clk), .D (new_AGEMA_signal_28559), .Q (new_AGEMA_signal_28560) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C (clk), .D (new_AGEMA_signal_28562), .Q (new_AGEMA_signal_28563) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C (clk), .D (new_AGEMA_signal_28565), .Q (new_AGEMA_signal_28566) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C (clk), .D (new_AGEMA_signal_28568), .Q (new_AGEMA_signal_28569) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C (clk), .D (new_AGEMA_signal_28571), .Q (new_AGEMA_signal_28572) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C (clk), .D (new_AGEMA_signal_28574), .Q (new_AGEMA_signal_28575) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C (clk), .D (new_AGEMA_signal_28577), .Q (new_AGEMA_signal_28578) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C (clk), .D (new_AGEMA_signal_28580), .Q (new_AGEMA_signal_28581) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C (clk), .D (new_AGEMA_signal_28583), .Q (new_AGEMA_signal_28584) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C (clk), .D (new_AGEMA_signal_28586), .Q (new_AGEMA_signal_28587) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C (clk), .D (new_AGEMA_signal_28589), .Q (new_AGEMA_signal_28590) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C (clk), .D (new_AGEMA_signal_28592), .Q (new_AGEMA_signal_28593) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C (clk), .D (new_AGEMA_signal_28595), .Q (new_AGEMA_signal_28596) ) ;
    buf_clk new_AGEMA_reg_buffer_7643 ( .C (clk), .D (new_AGEMA_signal_28598), .Q (new_AGEMA_signal_28599) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C (clk), .D (new_AGEMA_signal_28601), .Q (new_AGEMA_signal_28602) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C (clk), .D (new_AGEMA_signal_28604), .Q (new_AGEMA_signal_28605) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C (clk), .D (new_AGEMA_signal_28607), .Q (new_AGEMA_signal_28608) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C (clk), .D (new_AGEMA_signal_28610), .Q (new_AGEMA_signal_28611) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C (clk), .D (new_AGEMA_signal_28613), .Q (new_AGEMA_signal_28614) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C (clk), .D (new_AGEMA_signal_28616), .Q (new_AGEMA_signal_28617) ) ;
    buf_clk new_AGEMA_reg_buffer_7664 ( .C (clk), .D (new_AGEMA_signal_28619), .Q (new_AGEMA_signal_28620) ) ;
    buf_clk new_AGEMA_reg_buffer_7667 ( .C (clk), .D (new_AGEMA_signal_28622), .Q (new_AGEMA_signal_28623) ) ;
    buf_clk new_AGEMA_reg_buffer_7670 ( .C (clk), .D (new_AGEMA_signal_28625), .Q (new_AGEMA_signal_28626) ) ;
    buf_clk new_AGEMA_reg_buffer_7673 ( .C (clk), .D (new_AGEMA_signal_28628), .Q (new_AGEMA_signal_28629) ) ;
    buf_clk new_AGEMA_reg_buffer_7676 ( .C (clk), .D (new_AGEMA_signal_28631), .Q (new_AGEMA_signal_28632) ) ;
    buf_clk new_AGEMA_reg_buffer_7679 ( .C (clk), .D (new_AGEMA_signal_28634), .Q (new_AGEMA_signal_28635) ) ;
    buf_clk new_AGEMA_reg_buffer_7682 ( .C (clk), .D (new_AGEMA_signal_28637), .Q (new_AGEMA_signal_28638) ) ;
    buf_clk new_AGEMA_reg_buffer_7685 ( .C (clk), .D (new_AGEMA_signal_28640), .Q (new_AGEMA_signal_28641) ) ;
    buf_clk new_AGEMA_reg_buffer_7688 ( .C (clk), .D (new_AGEMA_signal_28643), .Q (new_AGEMA_signal_28644) ) ;
    buf_clk new_AGEMA_reg_buffer_7691 ( .C (clk), .D (new_AGEMA_signal_28646), .Q (new_AGEMA_signal_28647) ) ;
    buf_clk new_AGEMA_reg_buffer_7694 ( .C (clk), .D (new_AGEMA_signal_28649), .Q (new_AGEMA_signal_28650) ) ;
    buf_clk new_AGEMA_reg_buffer_7697 ( .C (clk), .D (new_AGEMA_signal_28652), .Q (new_AGEMA_signal_28653) ) ;
    buf_clk new_AGEMA_reg_buffer_7700 ( .C (clk), .D (new_AGEMA_signal_28655), .Q (new_AGEMA_signal_28656) ) ;
    buf_clk new_AGEMA_reg_buffer_7703 ( .C (clk), .D (new_AGEMA_signal_28658), .Q (new_AGEMA_signal_28659) ) ;
    buf_clk new_AGEMA_reg_buffer_7706 ( .C (clk), .D (new_AGEMA_signal_28661), .Q (new_AGEMA_signal_28662) ) ;
    buf_clk new_AGEMA_reg_buffer_7709 ( .C (clk), .D (new_AGEMA_signal_28664), .Q (new_AGEMA_signal_28665) ) ;
    buf_clk new_AGEMA_reg_buffer_7712 ( .C (clk), .D (new_AGEMA_signal_28667), .Q (new_AGEMA_signal_28668) ) ;
    buf_clk new_AGEMA_reg_buffer_7715 ( .C (clk), .D (new_AGEMA_signal_28670), .Q (new_AGEMA_signal_28671) ) ;
    buf_clk new_AGEMA_reg_buffer_7718 ( .C (clk), .D (new_AGEMA_signal_28673), .Q (new_AGEMA_signal_28674) ) ;
    buf_clk new_AGEMA_reg_buffer_7721 ( .C (clk), .D (new_AGEMA_signal_28676), .Q (new_AGEMA_signal_28677) ) ;
    buf_clk new_AGEMA_reg_buffer_7724 ( .C (clk), .D (new_AGEMA_signal_28679), .Q (new_AGEMA_signal_28680) ) ;
    buf_clk new_AGEMA_reg_buffer_7727 ( .C (clk), .D (new_AGEMA_signal_28682), .Q (new_AGEMA_signal_28683) ) ;
    buf_clk new_AGEMA_reg_buffer_7730 ( .C (clk), .D (new_AGEMA_signal_28685), .Q (new_AGEMA_signal_28686) ) ;
    buf_clk new_AGEMA_reg_buffer_7733 ( .C (clk), .D (new_AGEMA_signal_28688), .Q (new_AGEMA_signal_28689) ) ;
    buf_clk new_AGEMA_reg_buffer_7736 ( .C (clk), .D (new_AGEMA_signal_28691), .Q (new_AGEMA_signal_28692) ) ;
    buf_clk new_AGEMA_reg_buffer_7739 ( .C (clk), .D (new_AGEMA_signal_28694), .Q (new_AGEMA_signal_28695) ) ;
    buf_clk new_AGEMA_reg_buffer_7742 ( .C (clk), .D (new_AGEMA_signal_28697), .Q (new_AGEMA_signal_28698) ) ;
    buf_clk new_AGEMA_reg_buffer_7745 ( .C (clk), .D (new_AGEMA_signal_28700), .Q (new_AGEMA_signal_28701) ) ;
    buf_clk new_AGEMA_reg_buffer_7748 ( .C (clk), .D (new_AGEMA_signal_28703), .Q (new_AGEMA_signal_28704) ) ;
    buf_clk new_AGEMA_reg_buffer_7751 ( .C (clk), .D (new_AGEMA_signal_28706), .Q (new_AGEMA_signal_28707) ) ;
    buf_clk new_AGEMA_reg_buffer_7754 ( .C (clk), .D (new_AGEMA_signal_28709), .Q (new_AGEMA_signal_28710) ) ;
    buf_clk new_AGEMA_reg_buffer_7757 ( .C (clk), .D (new_AGEMA_signal_28712), .Q (new_AGEMA_signal_28713) ) ;
    buf_clk new_AGEMA_reg_buffer_7760 ( .C (clk), .D (new_AGEMA_signal_28715), .Q (new_AGEMA_signal_28716) ) ;
    buf_clk new_AGEMA_reg_buffer_7763 ( .C (clk), .D (new_AGEMA_signal_28718), .Q (new_AGEMA_signal_28719) ) ;
    buf_clk new_AGEMA_reg_buffer_7766 ( .C (clk), .D (new_AGEMA_signal_28721), .Q (new_AGEMA_signal_28722) ) ;
    buf_clk new_AGEMA_reg_buffer_7769 ( .C (clk), .D (new_AGEMA_signal_28724), .Q (new_AGEMA_signal_28725) ) ;
    buf_clk new_AGEMA_reg_buffer_7772 ( .C (clk), .D (new_AGEMA_signal_28727), .Q (new_AGEMA_signal_28728) ) ;
    buf_clk new_AGEMA_reg_buffer_7775 ( .C (clk), .D (new_AGEMA_signal_28730), .Q (new_AGEMA_signal_28731) ) ;
    buf_clk new_AGEMA_reg_buffer_7778 ( .C (clk), .D (new_AGEMA_signal_28733), .Q (new_AGEMA_signal_28734) ) ;
    buf_clk new_AGEMA_reg_buffer_7781 ( .C (clk), .D (new_AGEMA_signal_28736), .Q (new_AGEMA_signal_28737) ) ;
    buf_clk new_AGEMA_reg_buffer_7784 ( .C (clk), .D (new_AGEMA_signal_28739), .Q (new_AGEMA_signal_28740) ) ;
    buf_clk new_AGEMA_reg_buffer_7787 ( .C (clk), .D (new_AGEMA_signal_28742), .Q (new_AGEMA_signal_28743) ) ;
    buf_clk new_AGEMA_reg_buffer_7790 ( .C (clk), .D (new_AGEMA_signal_28745), .Q (new_AGEMA_signal_28746) ) ;
    buf_clk new_AGEMA_reg_buffer_7793 ( .C (clk), .D (new_AGEMA_signal_28748), .Q (new_AGEMA_signal_28749) ) ;
    buf_clk new_AGEMA_reg_buffer_7796 ( .C (clk), .D (new_AGEMA_signal_28751), .Q (new_AGEMA_signal_28752) ) ;
    buf_clk new_AGEMA_reg_buffer_7799 ( .C (clk), .D (new_AGEMA_signal_28754), .Q (new_AGEMA_signal_28755) ) ;
    buf_clk new_AGEMA_reg_buffer_7802 ( .C (clk), .D (new_AGEMA_signal_28757), .Q (new_AGEMA_signal_28758) ) ;
    buf_clk new_AGEMA_reg_buffer_7805 ( .C (clk), .D (new_AGEMA_signal_28760), .Q (new_AGEMA_signal_28761) ) ;
    buf_clk new_AGEMA_reg_buffer_7808 ( .C (clk), .D (new_AGEMA_signal_28763), .Q (new_AGEMA_signal_28764) ) ;
    buf_clk new_AGEMA_reg_buffer_7811 ( .C (clk), .D (new_AGEMA_signal_28766), .Q (new_AGEMA_signal_28767) ) ;
    buf_clk new_AGEMA_reg_buffer_7814 ( .C (clk), .D (new_AGEMA_signal_28769), .Q (new_AGEMA_signal_28770) ) ;
    buf_clk new_AGEMA_reg_buffer_7817 ( .C (clk), .D (new_AGEMA_signal_28772), .Q (new_AGEMA_signal_28773) ) ;
    buf_clk new_AGEMA_reg_buffer_7820 ( .C (clk), .D (new_AGEMA_signal_28775), .Q (new_AGEMA_signal_28776) ) ;
    buf_clk new_AGEMA_reg_buffer_7823 ( .C (clk), .D (new_AGEMA_signal_28778), .Q (new_AGEMA_signal_28779) ) ;
    buf_clk new_AGEMA_reg_buffer_7826 ( .C (clk), .D (new_AGEMA_signal_28781), .Q (new_AGEMA_signal_28782) ) ;
    buf_clk new_AGEMA_reg_buffer_7829 ( .C (clk), .D (new_AGEMA_signal_28784), .Q (new_AGEMA_signal_28785) ) ;
    buf_clk new_AGEMA_reg_buffer_7832 ( .C (clk), .D (new_AGEMA_signal_28787), .Q (new_AGEMA_signal_28788) ) ;
    buf_clk new_AGEMA_reg_buffer_7835 ( .C (clk), .D (new_AGEMA_signal_28790), .Q (new_AGEMA_signal_28791) ) ;
    buf_clk new_AGEMA_reg_buffer_7838 ( .C (clk), .D (new_AGEMA_signal_28793), .Q (new_AGEMA_signal_28794) ) ;
    buf_clk new_AGEMA_reg_buffer_7841 ( .C (clk), .D (new_AGEMA_signal_28796), .Q (new_AGEMA_signal_28797) ) ;
    buf_clk new_AGEMA_reg_buffer_7844 ( .C (clk), .D (new_AGEMA_signal_28799), .Q (new_AGEMA_signal_28800) ) ;
    buf_clk new_AGEMA_reg_buffer_7847 ( .C (clk), .D (new_AGEMA_signal_28802), .Q (new_AGEMA_signal_28803) ) ;
    buf_clk new_AGEMA_reg_buffer_7850 ( .C (clk), .D (new_AGEMA_signal_28805), .Q (new_AGEMA_signal_28806) ) ;
    buf_clk new_AGEMA_reg_buffer_7853 ( .C (clk), .D (new_AGEMA_signal_28808), .Q (new_AGEMA_signal_28809) ) ;
    buf_clk new_AGEMA_reg_buffer_7856 ( .C (clk), .D (new_AGEMA_signal_28811), .Q (new_AGEMA_signal_28812) ) ;
    buf_clk new_AGEMA_reg_buffer_7859 ( .C (clk), .D (new_AGEMA_signal_28814), .Q (new_AGEMA_signal_28815) ) ;
    buf_clk new_AGEMA_reg_buffer_7862 ( .C (clk), .D (new_AGEMA_signal_28817), .Q (new_AGEMA_signal_28818) ) ;
    buf_clk new_AGEMA_reg_buffer_7865 ( .C (clk), .D (new_AGEMA_signal_28820), .Q (new_AGEMA_signal_28821) ) ;
    buf_clk new_AGEMA_reg_buffer_7868 ( .C (clk), .D (new_AGEMA_signal_28823), .Q (new_AGEMA_signal_28824) ) ;
    buf_clk new_AGEMA_reg_buffer_7871 ( .C (clk), .D (new_AGEMA_signal_28826), .Q (new_AGEMA_signal_28827) ) ;
    buf_clk new_AGEMA_reg_buffer_7874 ( .C (clk), .D (new_AGEMA_signal_28829), .Q (new_AGEMA_signal_28830) ) ;
    buf_clk new_AGEMA_reg_buffer_7877 ( .C (clk), .D (new_AGEMA_signal_28832), .Q (new_AGEMA_signal_28833) ) ;
    buf_clk new_AGEMA_reg_buffer_7880 ( .C (clk), .D (new_AGEMA_signal_28835), .Q (new_AGEMA_signal_28836) ) ;
    buf_clk new_AGEMA_reg_buffer_7883 ( .C (clk), .D (new_AGEMA_signal_28838), .Q (new_AGEMA_signal_28839) ) ;
    buf_clk new_AGEMA_reg_buffer_7886 ( .C (clk), .D (new_AGEMA_signal_28841), .Q (new_AGEMA_signal_28842) ) ;
    buf_clk new_AGEMA_reg_buffer_7889 ( .C (clk), .D (new_AGEMA_signal_28844), .Q (new_AGEMA_signal_28845) ) ;
    buf_clk new_AGEMA_reg_buffer_7892 ( .C (clk), .D (new_AGEMA_signal_28847), .Q (new_AGEMA_signal_28848) ) ;
    buf_clk new_AGEMA_reg_buffer_7895 ( .C (clk), .D (new_AGEMA_signal_28850), .Q (new_AGEMA_signal_28851) ) ;
    buf_clk new_AGEMA_reg_buffer_7898 ( .C (clk), .D (new_AGEMA_signal_28853), .Q (new_AGEMA_signal_28854) ) ;
    buf_clk new_AGEMA_reg_buffer_7901 ( .C (clk), .D (new_AGEMA_signal_28856), .Q (new_AGEMA_signal_28857) ) ;
    buf_clk new_AGEMA_reg_buffer_7904 ( .C (clk), .D (new_AGEMA_signal_28859), .Q (new_AGEMA_signal_28860) ) ;
    buf_clk new_AGEMA_reg_buffer_7907 ( .C (clk), .D (new_AGEMA_signal_28862), .Q (new_AGEMA_signal_28863) ) ;
    buf_clk new_AGEMA_reg_buffer_7910 ( .C (clk), .D (new_AGEMA_signal_28865), .Q (new_AGEMA_signal_28866) ) ;
    buf_clk new_AGEMA_reg_buffer_7913 ( .C (clk), .D (new_AGEMA_signal_28868), .Q (new_AGEMA_signal_28869) ) ;
    buf_clk new_AGEMA_reg_buffer_7916 ( .C (clk), .D (new_AGEMA_signal_28871), .Q (new_AGEMA_signal_28872) ) ;
    buf_clk new_AGEMA_reg_buffer_7919 ( .C (clk), .D (new_AGEMA_signal_28874), .Q (new_AGEMA_signal_28875) ) ;
    buf_clk new_AGEMA_reg_buffer_7922 ( .C (clk), .D (new_AGEMA_signal_28877), .Q (new_AGEMA_signal_28878) ) ;
    buf_clk new_AGEMA_reg_buffer_7925 ( .C (clk), .D (new_AGEMA_signal_28880), .Q (new_AGEMA_signal_28881) ) ;
    buf_clk new_AGEMA_reg_buffer_7928 ( .C (clk), .D (new_AGEMA_signal_28883), .Q (new_AGEMA_signal_28884) ) ;
    buf_clk new_AGEMA_reg_buffer_7931 ( .C (clk), .D (new_AGEMA_signal_28886), .Q (new_AGEMA_signal_28887) ) ;
    buf_clk new_AGEMA_reg_buffer_7934 ( .C (clk), .D (new_AGEMA_signal_28889), .Q (new_AGEMA_signal_28890) ) ;
    buf_clk new_AGEMA_reg_buffer_7937 ( .C (clk), .D (new_AGEMA_signal_28892), .Q (new_AGEMA_signal_28893) ) ;
    buf_clk new_AGEMA_reg_buffer_7940 ( .C (clk), .D (new_AGEMA_signal_28895), .Q (new_AGEMA_signal_28896) ) ;
    buf_clk new_AGEMA_reg_buffer_7943 ( .C (clk), .D (new_AGEMA_signal_28898), .Q (new_AGEMA_signal_28899) ) ;
    buf_clk new_AGEMA_reg_buffer_7946 ( .C (clk), .D (new_AGEMA_signal_28901), .Q (new_AGEMA_signal_28902) ) ;
    buf_clk new_AGEMA_reg_buffer_7949 ( .C (clk), .D (new_AGEMA_signal_28904), .Q (new_AGEMA_signal_28905) ) ;
    buf_clk new_AGEMA_reg_buffer_7952 ( .C (clk), .D (new_AGEMA_signal_28907), .Q (new_AGEMA_signal_28908) ) ;
    buf_clk new_AGEMA_reg_buffer_7955 ( .C (clk), .D (new_AGEMA_signal_28910), .Q (new_AGEMA_signal_28911) ) ;
    buf_clk new_AGEMA_reg_buffer_7958 ( .C (clk), .D (new_AGEMA_signal_28913), .Q (new_AGEMA_signal_28914) ) ;
    buf_clk new_AGEMA_reg_buffer_7961 ( .C (clk), .D (new_AGEMA_signal_28916), .Q (new_AGEMA_signal_28917) ) ;
    buf_clk new_AGEMA_reg_buffer_7964 ( .C (clk), .D (new_AGEMA_signal_28919), .Q (new_AGEMA_signal_28920) ) ;
    buf_clk new_AGEMA_reg_buffer_7967 ( .C (clk), .D (new_AGEMA_signal_28922), .Q (new_AGEMA_signal_28923) ) ;
    buf_clk new_AGEMA_reg_buffer_7970 ( .C (clk), .D (new_AGEMA_signal_28925), .Q (new_AGEMA_signal_28926) ) ;
    buf_clk new_AGEMA_reg_buffer_7973 ( .C (clk), .D (new_AGEMA_signal_28928), .Q (new_AGEMA_signal_28929) ) ;
    buf_clk new_AGEMA_reg_buffer_7976 ( .C (clk), .D (new_AGEMA_signal_28931), .Q (new_AGEMA_signal_28932) ) ;
    buf_clk new_AGEMA_reg_buffer_7979 ( .C (clk), .D (new_AGEMA_signal_28934), .Q (new_AGEMA_signal_28935) ) ;
    buf_clk new_AGEMA_reg_buffer_7982 ( .C (clk), .D (new_AGEMA_signal_28937), .Q (new_AGEMA_signal_28938) ) ;
    buf_clk new_AGEMA_reg_buffer_7985 ( .C (clk), .D (new_AGEMA_signal_28940), .Q (new_AGEMA_signal_28941) ) ;
    buf_clk new_AGEMA_reg_buffer_7988 ( .C (clk), .D (new_AGEMA_signal_28943), .Q (new_AGEMA_signal_28944) ) ;
    buf_clk new_AGEMA_reg_buffer_7991 ( .C (clk), .D (new_AGEMA_signal_28946), .Q (new_AGEMA_signal_28947) ) ;
    buf_clk new_AGEMA_reg_buffer_7994 ( .C (clk), .D (new_AGEMA_signal_28949), .Q (new_AGEMA_signal_28950) ) ;
    buf_clk new_AGEMA_reg_buffer_7997 ( .C (clk), .D (new_AGEMA_signal_28952), .Q (new_AGEMA_signal_28953) ) ;
    buf_clk new_AGEMA_reg_buffer_8000 ( .C (clk), .D (new_AGEMA_signal_28955), .Q (new_AGEMA_signal_28956) ) ;
    buf_clk new_AGEMA_reg_buffer_8003 ( .C (clk), .D (new_AGEMA_signal_28958), .Q (new_AGEMA_signal_28959) ) ;
    buf_clk new_AGEMA_reg_buffer_8006 ( .C (clk), .D (new_AGEMA_signal_28961), .Q (new_AGEMA_signal_28962) ) ;
    buf_clk new_AGEMA_reg_buffer_8009 ( .C (clk), .D (new_AGEMA_signal_28964), .Q (new_AGEMA_signal_28965) ) ;
    buf_clk new_AGEMA_reg_buffer_8012 ( .C (clk), .D (new_AGEMA_signal_28967), .Q (new_AGEMA_signal_28968) ) ;
    buf_clk new_AGEMA_reg_buffer_8015 ( .C (clk), .D (new_AGEMA_signal_28970), .Q (new_AGEMA_signal_28971) ) ;
    buf_clk new_AGEMA_reg_buffer_8018 ( .C (clk), .D (new_AGEMA_signal_28973), .Q (new_AGEMA_signal_28974) ) ;
    buf_clk new_AGEMA_reg_buffer_8021 ( .C (clk), .D (new_AGEMA_signal_28976), .Q (new_AGEMA_signal_28977) ) ;
    buf_clk new_AGEMA_reg_buffer_8024 ( .C (clk), .D (new_AGEMA_signal_28979), .Q (new_AGEMA_signal_28980) ) ;
    buf_clk new_AGEMA_reg_buffer_8027 ( .C (clk), .D (new_AGEMA_signal_28982), .Q (new_AGEMA_signal_28983) ) ;
    buf_clk new_AGEMA_reg_buffer_8030 ( .C (clk), .D (new_AGEMA_signal_28985), .Q (new_AGEMA_signal_28986) ) ;
    buf_clk new_AGEMA_reg_buffer_8033 ( .C (clk), .D (new_AGEMA_signal_28988), .Q (new_AGEMA_signal_28989) ) ;
    buf_clk new_AGEMA_reg_buffer_8036 ( .C (clk), .D (new_AGEMA_signal_28991), .Q (new_AGEMA_signal_28992) ) ;
    buf_clk new_AGEMA_reg_buffer_8039 ( .C (clk), .D (new_AGEMA_signal_28994), .Q (new_AGEMA_signal_28995) ) ;
    buf_clk new_AGEMA_reg_buffer_8042 ( .C (clk), .D (new_AGEMA_signal_28997), .Q (new_AGEMA_signal_28998) ) ;
    buf_clk new_AGEMA_reg_buffer_8045 ( .C (clk), .D (new_AGEMA_signal_29000), .Q (new_AGEMA_signal_29001) ) ;
    buf_clk new_AGEMA_reg_buffer_8048 ( .C (clk), .D (new_AGEMA_signal_29003), .Q (new_AGEMA_signal_29004) ) ;
    buf_clk new_AGEMA_reg_buffer_8051 ( .C (clk), .D (new_AGEMA_signal_29006), .Q (new_AGEMA_signal_29007) ) ;
    buf_clk new_AGEMA_reg_buffer_8054 ( .C (clk), .D (new_AGEMA_signal_29009), .Q (new_AGEMA_signal_29010) ) ;
    buf_clk new_AGEMA_reg_buffer_8057 ( .C (clk), .D (new_AGEMA_signal_29012), .Q (new_AGEMA_signal_29013) ) ;
    buf_clk new_AGEMA_reg_buffer_8060 ( .C (clk), .D (new_AGEMA_signal_29015), .Q (new_AGEMA_signal_29016) ) ;
    buf_clk new_AGEMA_reg_buffer_8063 ( .C (clk), .D (new_AGEMA_signal_29018), .Q (new_AGEMA_signal_29019) ) ;
    buf_clk new_AGEMA_reg_buffer_8066 ( .C (clk), .D (new_AGEMA_signal_29021), .Q (new_AGEMA_signal_29022) ) ;
    buf_clk new_AGEMA_reg_buffer_8069 ( .C (clk), .D (new_AGEMA_signal_29024), .Q (new_AGEMA_signal_29025) ) ;
    buf_clk new_AGEMA_reg_buffer_8072 ( .C (clk), .D (new_AGEMA_signal_29027), .Q (new_AGEMA_signal_29028) ) ;
    buf_clk new_AGEMA_reg_buffer_8075 ( .C (clk), .D (new_AGEMA_signal_29030), .Q (new_AGEMA_signal_29031) ) ;
    buf_clk new_AGEMA_reg_buffer_8078 ( .C (clk), .D (new_AGEMA_signal_29033), .Q (new_AGEMA_signal_29034) ) ;
    buf_clk new_AGEMA_reg_buffer_8081 ( .C (clk), .D (new_AGEMA_signal_29036), .Q (new_AGEMA_signal_29037) ) ;
    buf_clk new_AGEMA_reg_buffer_8084 ( .C (clk), .D (new_AGEMA_signal_29039), .Q (new_AGEMA_signal_29040) ) ;
    buf_clk new_AGEMA_reg_buffer_8087 ( .C (clk), .D (new_AGEMA_signal_29042), .Q (new_AGEMA_signal_29043) ) ;
    buf_clk new_AGEMA_reg_buffer_8090 ( .C (clk), .D (new_AGEMA_signal_29045), .Q (new_AGEMA_signal_29046) ) ;
    buf_clk new_AGEMA_reg_buffer_8093 ( .C (clk), .D (new_AGEMA_signal_29048), .Q (new_AGEMA_signal_29049) ) ;
    buf_clk new_AGEMA_reg_buffer_8096 ( .C (clk), .D (new_AGEMA_signal_29051), .Q (new_AGEMA_signal_29052) ) ;
    buf_clk new_AGEMA_reg_buffer_8099 ( .C (clk), .D (new_AGEMA_signal_29054), .Q (new_AGEMA_signal_29055) ) ;
    buf_clk new_AGEMA_reg_buffer_8102 ( .C (clk), .D (new_AGEMA_signal_29057), .Q (new_AGEMA_signal_29058) ) ;
    buf_clk new_AGEMA_reg_buffer_8105 ( .C (clk), .D (new_AGEMA_signal_29060), .Q (new_AGEMA_signal_29061) ) ;
    buf_clk new_AGEMA_reg_buffer_8108 ( .C (clk), .D (new_AGEMA_signal_29063), .Q (new_AGEMA_signal_29064) ) ;
    buf_clk new_AGEMA_reg_buffer_8111 ( .C (clk), .D (new_AGEMA_signal_29066), .Q (new_AGEMA_signal_29067) ) ;
    buf_clk new_AGEMA_reg_buffer_8114 ( .C (clk), .D (new_AGEMA_signal_29069), .Q (new_AGEMA_signal_29070) ) ;
    buf_clk new_AGEMA_reg_buffer_8117 ( .C (clk), .D (new_AGEMA_signal_29072), .Q (new_AGEMA_signal_29073) ) ;
    buf_clk new_AGEMA_reg_buffer_8120 ( .C (clk), .D (new_AGEMA_signal_29075), .Q (new_AGEMA_signal_29076) ) ;
    buf_clk new_AGEMA_reg_buffer_8123 ( .C (clk), .D (new_AGEMA_signal_29078), .Q (new_AGEMA_signal_29079) ) ;
    buf_clk new_AGEMA_reg_buffer_8126 ( .C (clk), .D (new_AGEMA_signal_29081), .Q (new_AGEMA_signal_29082) ) ;
    buf_clk new_AGEMA_reg_buffer_8129 ( .C (clk), .D (new_AGEMA_signal_29084), .Q (new_AGEMA_signal_29085) ) ;
    buf_clk new_AGEMA_reg_buffer_8132 ( .C (clk), .D (new_AGEMA_signal_29087), .Q (new_AGEMA_signal_29088) ) ;
    buf_clk new_AGEMA_reg_buffer_8135 ( .C (clk), .D (new_AGEMA_signal_29090), .Q (new_AGEMA_signal_29091) ) ;
    buf_clk new_AGEMA_reg_buffer_8138 ( .C (clk), .D (new_AGEMA_signal_29093), .Q (new_AGEMA_signal_29094) ) ;
    buf_clk new_AGEMA_reg_buffer_8141 ( .C (clk), .D (new_AGEMA_signal_29096), .Q (new_AGEMA_signal_29097) ) ;
    buf_clk new_AGEMA_reg_buffer_8144 ( .C (clk), .D (new_AGEMA_signal_29099), .Q (new_AGEMA_signal_29100) ) ;
    buf_clk new_AGEMA_reg_buffer_8147 ( .C (clk), .D (new_AGEMA_signal_29102), .Q (new_AGEMA_signal_29103) ) ;
    buf_clk new_AGEMA_reg_buffer_8150 ( .C (clk), .D (new_AGEMA_signal_29105), .Q (new_AGEMA_signal_29106) ) ;
    buf_clk new_AGEMA_reg_buffer_8153 ( .C (clk), .D (new_AGEMA_signal_29108), .Q (new_AGEMA_signal_29109) ) ;
    buf_clk new_AGEMA_reg_buffer_8156 ( .C (clk), .D (new_AGEMA_signal_29111), .Q (new_AGEMA_signal_29112) ) ;
    buf_clk new_AGEMA_reg_buffer_8159 ( .C (clk), .D (new_AGEMA_signal_29114), .Q (new_AGEMA_signal_29115) ) ;
    buf_clk new_AGEMA_reg_buffer_8162 ( .C (clk), .D (new_AGEMA_signal_29117), .Q (new_AGEMA_signal_29118) ) ;
    buf_clk new_AGEMA_reg_buffer_8165 ( .C (clk), .D (new_AGEMA_signal_29120), .Q (new_AGEMA_signal_29121) ) ;
    buf_clk new_AGEMA_reg_buffer_8168 ( .C (clk), .D (new_AGEMA_signal_29123), .Q (new_AGEMA_signal_29124) ) ;
    buf_clk new_AGEMA_reg_buffer_8171 ( .C (clk), .D (new_AGEMA_signal_29126), .Q (new_AGEMA_signal_29127) ) ;
    buf_clk new_AGEMA_reg_buffer_8174 ( .C (clk), .D (new_AGEMA_signal_29129), .Q (new_AGEMA_signal_29130) ) ;
    buf_clk new_AGEMA_reg_buffer_8177 ( .C (clk), .D (new_AGEMA_signal_29132), .Q (new_AGEMA_signal_29133) ) ;
    buf_clk new_AGEMA_reg_buffer_8180 ( .C (clk), .D (new_AGEMA_signal_29135), .Q (new_AGEMA_signal_29136) ) ;
    buf_clk new_AGEMA_reg_buffer_8183 ( .C (clk), .D (new_AGEMA_signal_29138), .Q (new_AGEMA_signal_29139) ) ;
    buf_clk new_AGEMA_reg_buffer_8186 ( .C (clk), .D (new_AGEMA_signal_29141), .Q (new_AGEMA_signal_29142) ) ;
    buf_clk new_AGEMA_reg_buffer_8189 ( .C (clk), .D (new_AGEMA_signal_29144), .Q (new_AGEMA_signal_29145) ) ;
    buf_clk new_AGEMA_reg_buffer_8192 ( .C (clk), .D (new_AGEMA_signal_29147), .Q (new_AGEMA_signal_29148) ) ;
    buf_clk new_AGEMA_reg_buffer_8195 ( .C (clk), .D (new_AGEMA_signal_29150), .Q (new_AGEMA_signal_29151) ) ;
    buf_clk new_AGEMA_reg_buffer_8198 ( .C (clk), .D (new_AGEMA_signal_29153), .Q (new_AGEMA_signal_29154) ) ;
    buf_clk new_AGEMA_reg_buffer_8201 ( .C (clk), .D (new_AGEMA_signal_29156), .Q (new_AGEMA_signal_29157) ) ;
    buf_clk new_AGEMA_reg_buffer_8204 ( .C (clk), .D (new_AGEMA_signal_29159), .Q (new_AGEMA_signal_29160) ) ;
    buf_clk new_AGEMA_reg_buffer_8207 ( .C (clk), .D (new_AGEMA_signal_29162), .Q (new_AGEMA_signal_29163) ) ;
    buf_clk new_AGEMA_reg_buffer_8210 ( .C (clk), .D (new_AGEMA_signal_29165), .Q (new_AGEMA_signal_29166) ) ;
    buf_clk new_AGEMA_reg_buffer_8213 ( .C (clk), .D (new_AGEMA_signal_29168), .Q (new_AGEMA_signal_29169) ) ;
    buf_clk new_AGEMA_reg_buffer_8216 ( .C (clk), .D (new_AGEMA_signal_29171), .Q (new_AGEMA_signal_29172) ) ;
    buf_clk new_AGEMA_reg_buffer_8219 ( .C (clk), .D (new_AGEMA_signal_29174), .Q (new_AGEMA_signal_29175) ) ;
    buf_clk new_AGEMA_reg_buffer_8222 ( .C (clk), .D (new_AGEMA_signal_29177), .Q (new_AGEMA_signal_29178) ) ;
    buf_clk new_AGEMA_reg_buffer_8225 ( .C (clk), .D (new_AGEMA_signal_29180), .Q (new_AGEMA_signal_29181) ) ;
    buf_clk new_AGEMA_reg_buffer_8228 ( .C (clk), .D (new_AGEMA_signal_29183), .Q (new_AGEMA_signal_29184) ) ;
    buf_clk new_AGEMA_reg_buffer_8231 ( .C (clk), .D (new_AGEMA_signal_29186), .Q (new_AGEMA_signal_29187) ) ;
    buf_clk new_AGEMA_reg_buffer_8234 ( .C (clk), .D (new_AGEMA_signal_29189), .Q (new_AGEMA_signal_29190) ) ;
    buf_clk new_AGEMA_reg_buffer_8237 ( .C (clk), .D (new_AGEMA_signal_29192), .Q (new_AGEMA_signal_29193) ) ;
    buf_clk new_AGEMA_reg_buffer_8240 ( .C (clk), .D (new_AGEMA_signal_29195), .Q (new_AGEMA_signal_29196) ) ;
    buf_clk new_AGEMA_reg_buffer_8243 ( .C (clk), .D (new_AGEMA_signal_29198), .Q (new_AGEMA_signal_29199) ) ;
    buf_clk new_AGEMA_reg_buffer_8246 ( .C (clk), .D (new_AGEMA_signal_29201), .Q (new_AGEMA_signal_29202) ) ;
    buf_clk new_AGEMA_reg_buffer_8249 ( .C (clk), .D (new_AGEMA_signal_29204), .Q (new_AGEMA_signal_29205) ) ;
    buf_clk new_AGEMA_reg_buffer_8252 ( .C (clk), .D (new_AGEMA_signal_29207), .Q (new_AGEMA_signal_29208) ) ;
    buf_clk new_AGEMA_reg_buffer_8255 ( .C (clk), .D (new_AGEMA_signal_29210), .Q (new_AGEMA_signal_29211) ) ;
    buf_clk new_AGEMA_reg_buffer_8258 ( .C (clk), .D (new_AGEMA_signal_29213), .Q (new_AGEMA_signal_29214) ) ;
    buf_clk new_AGEMA_reg_buffer_8261 ( .C (clk), .D (new_AGEMA_signal_29216), .Q (new_AGEMA_signal_29217) ) ;
    buf_clk new_AGEMA_reg_buffer_8264 ( .C (clk), .D (new_AGEMA_signal_29219), .Q (new_AGEMA_signal_29220) ) ;
    buf_clk new_AGEMA_reg_buffer_8267 ( .C (clk), .D (new_AGEMA_signal_29222), .Q (new_AGEMA_signal_29223) ) ;
    buf_clk new_AGEMA_reg_buffer_8270 ( .C (clk), .D (new_AGEMA_signal_29225), .Q (new_AGEMA_signal_29226) ) ;
    buf_clk new_AGEMA_reg_buffer_8273 ( .C (clk), .D (new_AGEMA_signal_29228), .Q (new_AGEMA_signal_29229) ) ;
    buf_clk new_AGEMA_reg_buffer_8276 ( .C (clk), .D (new_AGEMA_signal_29231), .Q (new_AGEMA_signal_29232) ) ;
    buf_clk new_AGEMA_reg_buffer_8279 ( .C (clk), .D (new_AGEMA_signal_29234), .Q (new_AGEMA_signal_29235) ) ;
    buf_clk new_AGEMA_reg_buffer_8282 ( .C (clk), .D (new_AGEMA_signal_29237), .Q (new_AGEMA_signal_29238) ) ;
    buf_clk new_AGEMA_reg_buffer_8285 ( .C (clk), .D (new_AGEMA_signal_29240), .Q (new_AGEMA_signal_29241) ) ;
    buf_clk new_AGEMA_reg_buffer_8288 ( .C (clk), .D (new_AGEMA_signal_29243), .Q (new_AGEMA_signal_29244) ) ;
    buf_clk new_AGEMA_reg_buffer_8291 ( .C (clk), .D (new_AGEMA_signal_29246), .Q (new_AGEMA_signal_29247) ) ;
    buf_clk new_AGEMA_reg_buffer_8294 ( .C (clk), .D (new_AGEMA_signal_29249), .Q (new_AGEMA_signal_29250) ) ;
    buf_clk new_AGEMA_reg_buffer_8297 ( .C (clk), .D (new_AGEMA_signal_29252), .Q (new_AGEMA_signal_29253) ) ;
    buf_clk new_AGEMA_reg_buffer_8300 ( .C (clk), .D (new_AGEMA_signal_29255), .Q (new_AGEMA_signal_29256) ) ;
    buf_clk new_AGEMA_reg_buffer_8303 ( .C (clk), .D (new_AGEMA_signal_29258), .Q (new_AGEMA_signal_29259) ) ;
    buf_clk new_AGEMA_reg_buffer_8306 ( .C (clk), .D (new_AGEMA_signal_29261), .Q (new_AGEMA_signal_29262) ) ;
    buf_clk new_AGEMA_reg_buffer_8309 ( .C (clk), .D (new_AGEMA_signal_29264), .Q (new_AGEMA_signal_29265) ) ;
    buf_clk new_AGEMA_reg_buffer_8312 ( .C (clk), .D (new_AGEMA_signal_29267), .Q (new_AGEMA_signal_29268) ) ;
    buf_clk new_AGEMA_reg_buffer_8315 ( .C (clk), .D (new_AGEMA_signal_29270), .Q (new_AGEMA_signal_29271) ) ;
    buf_clk new_AGEMA_reg_buffer_8318 ( .C (clk), .D (new_AGEMA_signal_29273), .Q (new_AGEMA_signal_29274) ) ;
    buf_clk new_AGEMA_reg_buffer_8321 ( .C (clk), .D (new_AGEMA_signal_29276), .Q (new_AGEMA_signal_29277) ) ;
    buf_clk new_AGEMA_reg_buffer_8324 ( .C (clk), .D (new_AGEMA_signal_29279), .Q (new_AGEMA_signal_29280) ) ;
    buf_clk new_AGEMA_reg_buffer_8327 ( .C (clk), .D (new_AGEMA_signal_29282), .Q (new_AGEMA_signal_29283) ) ;
    buf_clk new_AGEMA_reg_buffer_8330 ( .C (clk), .D (new_AGEMA_signal_29285), .Q (new_AGEMA_signal_29286) ) ;
    buf_clk new_AGEMA_reg_buffer_8333 ( .C (clk), .D (new_AGEMA_signal_29288), .Q (new_AGEMA_signal_29289) ) ;
    buf_clk new_AGEMA_reg_buffer_8336 ( .C (clk), .D (new_AGEMA_signal_29291), .Q (new_AGEMA_signal_29292) ) ;
    buf_clk new_AGEMA_reg_buffer_8339 ( .C (clk), .D (new_AGEMA_signal_29294), .Q (new_AGEMA_signal_29295) ) ;
    buf_clk new_AGEMA_reg_buffer_8342 ( .C (clk), .D (new_AGEMA_signal_29297), .Q (new_AGEMA_signal_29298) ) ;
    buf_clk new_AGEMA_reg_buffer_8345 ( .C (clk), .D (new_AGEMA_signal_29300), .Q (new_AGEMA_signal_29301) ) ;
    buf_clk new_AGEMA_reg_buffer_8348 ( .C (clk), .D (new_AGEMA_signal_29303), .Q (new_AGEMA_signal_29304) ) ;
    buf_clk new_AGEMA_reg_buffer_8351 ( .C (clk), .D (new_AGEMA_signal_29306), .Q (new_AGEMA_signal_29307) ) ;
    buf_clk new_AGEMA_reg_buffer_8354 ( .C (clk), .D (new_AGEMA_signal_29309), .Q (new_AGEMA_signal_29310) ) ;
    buf_clk new_AGEMA_reg_buffer_8357 ( .C (clk), .D (new_AGEMA_signal_29312), .Q (new_AGEMA_signal_29313) ) ;
    buf_clk new_AGEMA_reg_buffer_8360 ( .C (clk), .D (new_AGEMA_signal_29315), .Q (new_AGEMA_signal_29316) ) ;
    buf_clk new_AGEMA_reg_buffer_8363 ( .C (clk), .D (new_AGEMA_signal_29318), .Q (new_AGEMA_signal_29319) ) ;
    buf_clk new_AGEMA_reg_buffer_8366 ( .C (clk), .D (new_AGEMA_signal_29321), .Q (new_AGEMA_signal_29322) ) ;
    buf_clk new_AGEMA_reg_buffer_8369 ( .C (clk), .D (new_AGEMA_signal_29324), .Q (new_AGEMA_signal_29325) ) ;
    buf_clk new_AGEMA_reg_buffer_8372 ( .C (clk), .D (new_AGEMA_signal_29327), .Q (new_AGEMA_signal_29328) ) ;
    buf_clk new_AGEMA_reg_buffer_8375 ( .C (clk), .D (new_AGEMA_signal_29330), .Q (new_AGEMA_signal_29331) ) ;
    buf_clk new_AGEMA_reg_buffer_8378 ( .C (clk), .D (new_AGEMA_signal_29333), .Q (new_AGEMA_signal_29334) ) ;
    buf_clk new_AGEMA_reg_buffer_8381 ( .C (clk), .D (new_AGEMA_signal_29336), .Q (new_AGEMA_signal_29337) ) ;
    buf_clk new_AGEMA_reg_buffer_8384 ( .C (clk), .D (new_AGEMA_signal_29339), .Q (new_AGEMA_signal_29340) ) ;
    buf_clk new_AGEMA_reg_buffer_8387 ( .C (clk), .D (new_AGEMA_signal_29342), .Q (new_AGEMA_signal_29343) ) ;
    buf_clk new_AGEMA_reg_buffer_8390 ( .C (clk), .D (new_AGEMA_signal_29345), .Q (new_AGEMA_signal_29346) ) ;
    buf_clk new_AGEMA_reg_buffer_8393 ( .C (clk), .D (new_AGEMA_signal_29348), .Q (new_AGEMA_signal_29349) ) ;
    buf_clk new_AGEMA_reg_buffer_8396 ( .C (clk), .D (new_AGEMA_signal_29351), .Q (new_AGEMA_signal_29352) ) ;
    buf_clk new_AGEMA_reg_buffer_8399 ( .C (clk), .D (new_AGEMA_signal_29354), .Q (new_AGEMA_signal_29355) ) ;
    buf_clk new_AGEMA_reg_buffer_8402 ( .C (clk), .D (new_AGEMA_signal_29357), .Q (new_AGEMA_signal_29358) ) ;
    buf_clk new_AGEMA_reg_buffer_8405 ( .C (clk), .D (new_AGEMA_signal_29360), .Q (new_AGEMA_signal_29361) ) ;
    buf_clk new_AGEMA_reg_buffer_8408 ( .C (clk), .D (new_AGEMA_signal_29363), .Q (new_AGEMA_signal_29364) ) ;
    buf_clk new_AGEMA_reg_buffer_8411 ( .C (clk), .D (new_AGEMA_signal_29366), .Q (new_AGEMA_signal_29367) ) ;
    buf_clk new_AGEMA_reg_buffer_8414 ( .C (clk), .D (new_AGEMA_signal_29369), .Q (new_AGEMA_signal_29370) ) ;
    buf_clk new_AGEMA_reg_buffer_8417 ( .C (clk), .D (new_AGEMA_signal_29372), .Q (new_AGEMA_signal_29373) ) ;
    buf_clk new_AGEMA_reg_buffer_8420 ( .C (clk), .D (new_AGEMA_signal_29375), .Q (new_AGEMA_signal_29376) ) ;
    buf_clk new_AGEMA_reg_buffer_8423 ( .C (clk), .D (new_AGEMA_signal_29378), .Q (new_AGEMA_signal_29379) ) ;
    buf_clk new_AGEMA_reg_buffer_8426 ( .C (clk), .D (new_AGEMA_signal_29381), .Q (new_AGEMA_signal_29382) ) ;
    buf_clk new_AGEMA_reg_buffer_8429 ( .C (clk), .D (new_AGEMA_signal_29384), .Q (new_AGEMA_signal_29385) ) ;
    buf_clk new_AGEMA_reg_buffer_8432 ( .C (clk), .D (new_AGEMA_signal_29387), .Q (new_AGEMA_signal_29388) ) ;
    buf_clk new_AGEMA_reg_buffer_8435 ( .C (clk), .D (new_AGEMA_signal_29390), .Q (new_AGEMA_signal_29391) ) ;
    buf_clk new_AGEMA_reg_buffer_8438 ( .C (clk), .D (new_AGEMA_signal_29393), .Q (new_AGEMA_signal_29394) ) ;
    buf_clk new_AGEMA_reg_buffer_8441 ( .C (clk), .D (new_AGEMA_signal_29396), .Q (new_AGEMA_signal_29397) ) ;
    buf_clk new_AGEMA_reg_buffer_8444 ( .C (clk), .D (new_AGEMA_signal_29399), .Q (new_AGEMA_signal_29400) ) ;
    buf_clk new_AGEMA_reg_buffer_8447 ( .C (clk), .D (new_AGEMA_signal_29402), .Q (new_AGEMA_signal_29403) ) ;
    buf_clk new_AGEMA_reg_buffer_8450 ( .C (clk), .D (new_AGEMA_signal_29405), .Q (new_AGEMA_signal_29406) ) ;
    buf_clk new_AGEMA_reg_buffer_8453 ( .C (clk), .D (new_AGEMA_signal_29408), .Q (new_AGEMA_signal_29409) ) ;
    buf_clk new_AGEMA_reg_buffer_8456 ( .C (clk), .D (new_AGEMA_signal_29411), .Q (new_AGEMA_signal_29412) ) ;
    buf_clk new_AGEMA_reg_buffer_8459 ( .C (clk), .D (new_AGEMA_signal_29414), .Q (new_AGEMA_signal_29415) ) ;
    buf_clk new_AGEMA_reg_buffer_8462 ( .C (clk), .D (new_AGEMA_signal_29417), .Q (new_AGEMA_signal_29418) ) ;
    buf_clk new_AGEMA_reg_buffer_8465 ( .C (clk), .D (new_AGEMA_signal_29420), .Q (new_AGEMA_signal_29421) ) ;
    buf_clk new_AGEMA_reg_buffer_8468 ( .C (clk), .D (new_AGEMA_signal_29423), .Q (new_AGEMA_signal_29424) ) ;
    buf_clk new_AGEMA_reg_buffer_8471 ( .C (clk), .D (new_AGEMA_signal_29426), .Q (new_AGEMA_signal_29427) ) ;
    buf_clk new_AGEMA_reg_buffer_8474 ( .C (clk), .D (new_AGEMA_signal_29429), .Q (new_AGEMA_signal_29430) ) ;
    buf_clk new_AGEMA_reg_buffer_8477 ( .C (clk), .D (new_AGEMA_signal_29432), .Q (new_AGEMA_signal_29433) ) ;
    buf_clk new_AGEMA_reg_buffer_8480 ( .C (clk), .D (new_AGEMA_signal_29435), .Q (new_AGEMA_signal_29436) ) ;
    buf_clk new_AGEMA_reg_buffer_8483 ( .C (clk), .D (new_AGEMA_signal_29438), .Q (new_AGEMA_signal_29439) ) ;
    buf_clk new_AGEMA_reg_buffer_8486 ( .C (clk), .D (new_AGEMA_signal_29441), .Q (new_AGEMA_signal_29442) ) ;
    buf_clk new_AGEMA_reg_buffer_8489 ( .C (clk), .D (new_AGEMA_signal_29444), .Q (new_AGEMA_signal_29445) ) ;
    buf_clk new_AGEMA_reg_buffer_8492 ( .C (clk), .D (new_AGEMA_signal_29447), .Q (new_AGEMA_signal_29448) ) ;
    buf_clk new_AGEMA_reg_buffer_8495 ( .C (clk), .D (new_AGEMA_signal_29450), .Q (new_AGEMA_signal_29451) ) ;
    buf_clk new_AGEMA_reg_buffer_8498 ( .C (clk), .D (new_AGEMA_signal_29453), .Q (new_AGEMA_signal_29454) ) ;
    buf_clk new_AGEMA_reg_buffer_8501 ( .C (clk), .D (new_AGEMA_signal_29456), .Q (new_AGEMA_signal_29457) ) ;
    buf_clk new_AGEMA_reg_buffer_8504 ( .C (clk), .D (new_AGEMA_signal_29459), .Q (new_AGEMA_signal_29460) ) ;
    buf_clk new_AGEMA_reg_buffer_8507 ( .C (clk), .D (new_AGEMA_signal_29462), .Q (new_AGEMA_signal_29463) ) ;
    buf_clk new_AGEMA_reg_buffer_8510 ( .C (clk), .D (new_AGEMA_signal_29465), .Q (new_AGEMA_signal_29466) ) ;
    buf_clk new_AGEMA_reg_buffer_8513 ( .C (clk), .D (new_AGEMA_signal_29468), .Q (new_AGEMA_signal_29469) ) ;
    buf_clk new_AGEMA_reg_buffer_8516 ( .C (clk), .D (new_AGEMA_signal_29471), .Q (new_AGEMA_signal_29472) ) ;
    buf_clk new_AGEMA_reg_buffer_8519 ( .C (clk), .D (new_AGEMA_signal_29474), .Q (new_AGEMA_signal_29475) ) ;
    buf_clk new_AGEMA_reg_buffer_8522 ( .C (clk), .D (new_AGEMA_signal_29477), .Q (new_AGEMA_signal_29478) ) ;
    buf_clk new_AGEMA_reg_buffer_8525 ( .C (clk), .D (new_AGEMA_signal_29480), .Q (new_AGEMA_signal_29481) ) ;
    buf_clk new_AGEMA_reg_buffer_8528 ( .C (clk), .D (new_AGEMA_signal_29483), .Q (new_AGEMA_signal_29484) ) ;
    buf_clk new_AGEMA_reg_buffer_8531 ( .C (clk), .D (new_AGEMA_signal_29486), .Q (new_AGEMA_signal_29487) ) ;
    buf_clk new_AGEMA_reg_buffer_8534 ( .C (clk), .D (new_AGEMA_signal_29489), .Q (new_AGEMA_signal_29490) ) ;
    buf_clk new_AGEMA_reg_buffer_8537 ( .C (clk), .D (new_AGEMA_signal_29492), .Q (new_AGEMA_signal_29493) ) ;
    buf_clk new_AGEMA_reg_buffer_8540 ( .C (clk), .D (new_AGEMA_signal_29495), .Q (new_AGEMA_signal_29496) ) ;
    buf_clk new_AGEMA_reg_buffer_8543 ( .C (clk), .D (new_AGEMA_signal_29498), .Q (new_AGEMA_signal_29499) ) ;
    buf_clk new_AGEMA_reg_buffer_8546 ( .C (clk), .D (new_AGEMA_signal_29501), .Q (new_AGEMA_signal_29502) ) ;
    buf_clk new_AGEMA_reg_buffer_8549 ( .C (clk), .D (new_AGEMA_signal_29504), .Q (new_AGEMA_signal_29505) ) ;
    buf_clk new_AGEMA_reg_buffer_8552 ( .C (clk), .D (new_AGEMA_signal_29507), .Q (new_AGEMA_signal_29508) ) ;
    buf_clk new_AGEMA_reg_buffer_8555 ( .C (clk), .D (new_AGEMA_signal_29510), .Q (new_AGEMA_signal_29511) ) ;
    buf_clk new_AGEMA_reg_buffer_8558 ( .C (clk), .D (new_AGEMA_signal_29513), .Q (new_AGEMA_signal_29514) ) ;
    buf_clk new_AGEMA_reg_buffer_8561 ( .C (clk), .D (new_AGEMA_signal_29516), .Q (new_AGEMA_signal_29517) ) ;
    buf_clk new_AGEMA_reg_buffer_8564 ( .C (clk), .D (new_AGEMA_signal_29519), .Q (new_AGEMA_signal_29520) ) ;
    buf_clk new_AGEMA_reg_buffer_8567 ( .C (clk), .D (new_AGEMA_signal_29522), .Q (new_AGEMA_signal_29523) ) ;
    buf_clk new_AGEMA_reg_buffer_8570 ( .C (clk), .D (new_AGEMA_signal_29525), .Q (new_AGEMA_signal_29526) ) ;
    buf_clk new_AGEMA_reg_buffer_8573 ( .C (clk), .D (new_AGEMA_signal_29528), .Q (new_AGEMA_signal_29529) ) ;
    buf_clk new_AGEMA_reg_buffer_8576 ( .C (clk), .D (new_AGEMA_signal_29531), .Q (new_AGEMA_signal_29532) ) ;
    buf_clk new_AGEMA_reg_buffer_8579 ( .C (clk), .D (new_AGEMA_signal_29534), .Q (new_AGEMA_signal_29535) ) ;
    buf_clk new_AGEMA_reg_buffer_8582 ( .C (clk), .D (new_AGEMA_signal_29537), .Q (new_AGEMA_signal_29538) ) ;
    buf_clk new_AGEMA_reg_buffer_8585 ( .C (clk), .D (new_AGEMA_signal_29540), .Q (new_AGEMA_signal_29541) ) ;
    buf_clk new_AGEMA_reg_buffer_8588 ( .C (clk), .D (new_AGEMA_signal_29543), .Q (new_AGEMA_signal_29544) ) ;
    buf_clk new_AGEMA_reg_buffer_8591 ( .C (clk), .D (new_AGEMA_signal_29546), .Q (new_AGEMA_signal_29547) ) ;
    buf_clk new_AGEMA_reg_buffer_8594 ( .C (clk), .D (new_AGEMA_signal_29549), .Q (new_AGEMA_signal_29550) ) ;
    buf_clk new_AGEMA_reg_buffer_8597 ( .C (clk), .D (new_AGEMA_signal_29552), .Q (new_AGEMA_signal_29553) ) ;
    buf_clk new_AGEMA_reg_buffer_8600 ( .C (clk), .D (new_AGEMA_signal_29555), .Q (new_AGEMA_signal_29556) ) ;
    buf_clk new_AGEMA_reg_buffer_8603 ( .C (clk), .D (new_AGEMA_signal_29558), .Q (new_AGEMA_signal_29559) ) ;
    buf_clk new_AGEMA_reg_buffer_8606 ( .C (clk), .D (new_AGEMA_signal_29561), .Q (new_AGEMA_signal_29562) ) ;
    buf_clk new_AGEMA_reg_buffer_8609 ( .C (clk), .D (new_AGEMA_signal_29564), .Q (new_AGEMA_signal_29565) ) ;
    buf_clk new_AGEMA_reg_buffer_8612 ( .C (clk), .D (new_AGEMA_signal_29567), .Q (new_AGEMA_signal_29568) ) ;
    buf_clk new_AGEMA_reg_buffer_8615 ( .C (clk), .D (new_AGEMA_signal_29570), .Q (new_AGEMA_signal_29571) ) ;
    buf_clk new_AGEMA_reg_buffer_8618 ( .C (clk), .D (new_AGEMA_signal_29573), .Q (new_AGEMA_signal_29574) ) ;
    buf_clk new_AGEMA_reg_buffer_8621 ( .C (clk), .D (new_AGEMA_signal_29576), .Q (new_AGEMA_signal_29577) ) ;
    buf_clk new_AGEMA_reg_buffer_8624 ( .C (clk), .D (new_AGEMA_signal_29579), .Q (new_AGEMA_signal_29580) ) ;
    buf_clk new_AGEMA_reg_buffer_8627 ( .C (clk), .D (new_AGEMA_signal_29582), .Q (new_AGEMA_signal_29583) ) ;
    buf_clk new_AGEMA_reg_buffer_8630 ( .C (clk), .D (new_AGEMA_signal_29585), .Q (new_AGEMA_signal_29586) ) ;
    buf_clk new_AGEMA_reg_buffer_8633 ( .C (clk), .D (new_AGEMA_signal_29588), .Q (new_AGEMA_signal_29589) ) ;
    buf_clk new_AGEMA_reg_buffer_8636 ( .C (clk), .D (new_AGEMA_signal_29591), .Q (new_AGEMA_signal_29592) ) ;
    buf_clk new_AGEMA_reg_buffer_8639 ( .C (clk), .D (new_AGEMA_signal_29594), .Q (new_AGEMA_signal_29595) ) ;
    buf_clk new_AGEMA_reg_buffer_8642 ( .C (clk), .D (new_AGEMA_signal_29597), .Q (new_AGEMA_signal_29598) ) ;
    buf_clk new_AGEMA_reg_buffer_8645 ( .C (clk), .D (new_AGEMA_signal_29600), .Q (new_AGEMA_signal_29601) ) ;
    buf_clk new_AGEMA_reg_buffer_8648 ( .C (clk), .D (new_AGEMA_signal_29603), .Q (new_AGEMA_signal_29604) ) ;
    buf_clk new_AGEMA_reg_buffer_8651 ( .C (clk), .D (new_AGEMA_signal_29606), .Q (new_AGEMA_signal_29607) ) ;
    buf_clk new_AGEMA_reg_buffer_8654 ( .C (clk), .D (new_AGEMA_signal_29609), .Q (new_AGEMA_signal_29610) ) ;
    buf_clk new_AGEMA_reg_buffer_8657 ( .C (clk), .D (new_AGEMA_signal_29612), .Q (new_AGEMA_signal_29613) ) ;
    buf_clk new_AGEMA_reg_buffer_8660 ( .C (clk), .D (new_AGEMA_signal_29615), .Q (new_AGEMA_signal_29616) ) ;
    buf_clk new_AGEMA_reg_buffer_8663 ( .C (clk), .D (new_AGEMA_signal_29618), .Q (new_AGEMA_signal_29619) ) ;
    buf_clk new_AGEMA_reg_buffer_8666 ( .C (clk), .D (new_AGEMA_signal_29621), .Q (new_AGEMA_signal_29622) ) ;
    buf_clk new_AGEMA_reg_buffer_8669 ( .C (clk), .D (new_AGEMA_signal_29624), .Q (new_AGEMA_signal_29625) ) ;
    buf_clk new_AGEMA_reg_buffer_8672 ( .C (clk), .D (new_AGEMA_signal_29627), .Q (new_AGEMA_signal_29628) ) ;
    buf_clk new_AGEMA_reg_buffer_8675 ( .C (clk), .D (new_AGEMA_signal_29630), .Q (new_AGEMA_signal_29631) ) ;
    buf_clk new_AGEMA_reg_buffer_8678 ( .C (clk), .D (new_AGEMA_signal_29633), .Q (new_AGEMA_signal_29634) ) ;
    buf_clk new_AGEMA_reg_buffer_8681 ( .C (clk), .D (new_AGEMA_signal_29636), .Q (new_AGEMA_signal_29637) ) ;
    buf_clk new_AGEMA_reg_buffer_8684 ( .C (clk), .D (new_AGEMA_signal_29639), .Q (new_AGEMA_signal_29640) ) ;
    buf_clk new_AGEMA_reg_buffer_8687 ( .C (clk), .D (new_AGEMA_signal_29642), .Q (new_AGEMA_signal_29643) ) ;
    buf_clk new_AGEMA_reg_buffer_8690 ( .C (clk), .D (new_AGEMA_signal_29645), .Q (new_AGEMA_signal_29646) ) ;
    buf_clk new_AGEMA_reg_buffer_8693 ( .C (clk), .D (new_AGEMA_signal_29648), .Q (new_AGEMA_signal_29649) ) ;
    buf_clk new_AGEMA_reg_buffer_8696 ( .C (clk), .D (new_AGEMA_signal_29651), .Q (new_AGEMA_signal_29652) ) ;
    buf_clk new_AGEMA_reg_buffer_8699 ( .C (clk), .D (new_AGEMA_signal_29654), .Q (new_AGEMA_signal_29655) ) ;
    buf_clk new_AGEMA_reg_buffer_8702 ( .C (clk), .D (new_AGEMA_signal_29657), .Q (new_AGEMA_signal_29658) ) ;
    buf_clk new_AGEMA_reg_buffer_8705 ( .C (clk), .D (new_AGEMA_signal_29660), .Q (new_AGEMA_signal_29661) ) ;
    buf_clk new_AGEMA_reg_buffer_8708 ( .C (clk), .D (new_AGEMA_signal_29663), .Q (new_AGEMA_signal_29664) ) ;
    buf_clk new_AGEMA_reg_buffer_8711 ( .C (clk), .D (new_AGEMA_signal_29666), .Q (new_AGEMA_signal_29667) ) ;
    buf_clk new_AGEMA_reg_buffer_8714 ( .C (clk), .D (new_AGEMA_signal_29669), .Q (new_AGEMA_signal_29670) ) ;
    buf_clk new_AGEMA_reg_buffer_8717 ( .C (clk), .D (new_AGEMA_signal_29672), .Q (new_AGEMA_signal_29673) ) ;
    buf_clk new_AGEMA_reg_buffer_8720 ( .C (clk), .D (new_AGEMA_signal_29675), .Q (new_AGEMA_signal_29676) ) ;
    buf_clk new_AGEMA_reg_buffer_8723 ( .C (clk), .D (new_AGEMA_signal_29678), .Q (new_AGEMA_signal_29679) ) ;
    buf_clk new_AGEMA_reg_buffer_8726 ( .C (clk), .D (new_AGEMA_signal_29681), .Q (new_AGEMA_signal_29682) ) ;
    buf_clk new_AGEMA_reg_buffer_8729 ( .C (clk), .D (new_AGEMA_signal_29684), .Q (new_AGEMA_signal_29685) ) ;
    buf_clk new_AGEMA_reg_buffer_8732 ( .C (clk), .D (new_AGEMA_signal_29687), .Q (new_AGEMA_signal_29688) ) ;
    buf_clk new_AGEMA_reg_buffer_8735 ( .C (clk), .D (new_AGEMA_signal_29690), .Q (new_AGEMA_signal_29691) ) ;
    buf_clk new_AGEMA_reg_buffer_8738 ( .C (clk), .D (new_AGEMA_signal_29693), .Q (new_AGEMA_signal_29694) ) ;
    buf_clk new_AGEMA_reg_buffer_8741 ( .C (clk), .D (new_AGEMA_signal_29696), .Q (new_AGEMA_signal_29697) ) ;
    buf_clk new_AGEMA_reg_buffer_8744 ( .C (clk), .D (new_AGEMA_signal_29699), .Q (new_AGEMA_signal_29700) ) ;
    buf_clk new_AGEMA_reg_buffer_8747 ( .C (clk), .D (new_AGEMA_signal_29702), .Q (new_AGEMA_signal_29703) ) ;
    buf_clk new_AGEMA_reg_buffer_8750 ( .C (clk), .D (new_AGEMA_signal_29705), .Q (new_AGEMA_signal_29706) ) ;
    buf_clk new_AGEMA_reg_buffer_8753 ( .C (clk), .D (new_AGEMA_signal_29708), .Q (new_AGEMA_signal_29709) ) ;
    buf_clk new_AGEMA_reg_buffer_8756 ( .C (clk), .D (new_AGEMA_signal_29711), .Q (new_AGEMA_signal_29712) ) ;
    buf_clk new_AGEMA_reg_buffer_8759 ( .C (clk), .D (new_AGEMA_signal_29714), .Q (new_AGEMA_signal_29715) ) ;
    buf_clk new_AGEMA_reg_buffer_8762 ( .C (clk), .D (new_AGEMA_signal_29717), .Q (new_AGEMA_signal_29718) ) ;
    buf_clk new_AGEMA_reg_buffer_8765 ( .C (clk), .D (new_AGEMA_signal_29720), .Q (new_AGEMA_signal_29721) ) ;
    buf_clk new_AGEMA_reg_buffer_8768 ( .C (clk), .D (new_AGEMA_signal_29723), .Q (new_AGEMA_signal_29724) ) ;
    buf_clk new_AGEMA_reg_buffer_8771 ( .C (clk), .D (new_AGEMA_signal_29726), .Q (new_AGEMA_signal_29727) ) ;
    buf_clk new_AGEMA_reg_buffer_8774 ( .C (clk), .D (new_AGEMA_signal_29729), .Q (new_AGEMA_signal_29730) ) ;
    buf_clk new_AGEMA_reg_buffer_8777 ( .C (clk), .D (new_AGEMA_signal_29732), .Q (new_AGEMA_signal_29733) ) ;
    buf_clk new_AGEMA_reg_buffer_8780 ( .C (clk), .D (new_AGEMA_signal_29735), .Q (new_AGEMA_signal_29736) ) ;
    buf_clk new_AGEMA_reg_buffer_8783 ( .C (clk), .D (new_AGEMA_signal_29738), .Q (new_AGEMA_signal_29739) ) ;
    buf_clk new_AGEMA_reg_buffer_8786 ( .C (clk), .D (new_AGEMA_signal_29741), .Q (new_AGEMA_signal_29742) ) ;
    buf_clk new_AGEMA_reg_buffer_8789 ( .C (clk), .D (new_AGEMA_signal_29744), .Q (new_AGEMA_signal_29745) ) ;
    buf_clk new_AGEMA_reg_buffer_8792 ( .C (clk), .D (new_AGEMA_signal_29747), .Q (new_AGEMA_signal_29748) ) ;
    buf_clk new_AGEMA_reg_buffer_8795 ( .C (clk), .D (new_AGEMA_signal_29750), .Q (new_AGEMA_signal_29751) ) ;
    buf_clk new_AGEMA_reg_buffer_8798 ( .C (clk), .D (new_AGEMA_signal_29753), .Q (new_AGEMA_signal_29754) ) ;
    buf_clk new_AGEMA_reg_buffer_8801 ( .C (clk), .D (new_AGEMA_signal_29756), .Q (new_AGEMA_signal_29757) ) ;
    buf_clk new_AGEMA_reg_buffer_8804 ( .C (clk), .D (new_AGEMA_signal_29759), .Q (new_AGEMA_signal_29760) ) ;
    buf_clk new_AGEMA_reg_buffer_8807 ( .C (clk), .D (new_AGEMA_signal_29762), .Q (new_AGEMA_signal_29763) ) ;
    buf_clk new_AGEMA_reg_buffer_8810 ( .C (clk), .D (new_AGEMA_signal_29765), .Q (new_AGEMA_signal_29766) ) ;
    buf_clk new_AGEMA_reg_buffer_8813 ( .C (clk), .D (new_AGEMA_signal_29768), .Q (new_AGEMA_signal_29769) ) ;
    buf_clk new_AGEMA_reg_buffer_8816 ( .C (clk), .D (new_AGEMA_signal_29771), .Q (new_AGEMA_signal_29772) ) ;
    buf_clk new_AGEMA_reg_buffer_8819 ( .C (clk), .D (new_AGEMA_signal_29774), .Q (new_AGEMA_signal_29775) ) ;
    buf_clk new_AGEMA_reg_buffer_8822 ( .C (clk), .D (new_AGEMA_signal_29777), .Q (new_AGEMA_signal_29778) ) ;
    buf_clk new_AGEMA_reg_buffer_8825 ( .C (clk), .D (new_AGEMA_signal_29780), .Q (new_AGEMA_signal_29781) ) ;
    buf_clk new_AGEMA_reg_buffer_8828 ( .C (clk), .D (new_AGEMA_signal_29783), .Q (new_AGEMA_signal_29784) ) ;
    buf_clk new_AGEMA_reg_buffer_8831 ( .C (clk), .D (new_AGEMA_signal_29786), .Q (new_AGEMA_signal_29787) ) ;
    buf_clk new_AGEMA_reg_buffer_8834 ( .C (clk), .D (new_AGEMA_signal_29789), .Q (new_AGEMA_signal_29790) ) ;
    buf_clk new_AGEMA_reg_buffer_8837 ( .C (clk), .D (new_AGEMA_signal_29792), .Q (new_AGEMA_signal_29793) ) ;
    buf_clk new_AGEMA_reg_buffer_8840 ( .C (clk), .D (new_AGEMA_signal_29795), .Q (new_AGEMA_signal_29796) ) ;
    buf_clk new_AGEMA_reg_buffer_8843 ( .C (clk), .D (new_AGEMA_signal_29798), .Q (new_AGEMA_signal_29799) ) ;
    buf_clk new_AGEMA_reg_buffer_8846 ( .C (clk), .D (new_AGEMA_signal_29801), .Q (new_AGEMA_signal_29802) ) ;
    buf_clk new_AGEMA_reg_buffer_8849 ( .C (clk), .D (new_AGEMA_signal_29804), .Q (new_AGEMA_signal_29805) ) ;
    buf_clk new_AGEMA_reg_buffer_8852 ( .C (clk), .D (new_AGEMA_signal_29807), .Q (new_AGEMA_signal_29808) ) ;
    buf_clk new_AGEMA_reg_buffer_8855 ( .C (clk), .D (new_AGEMA_signal_29810), .Q (new_AGEMA_signal_29811) ) ;
    buf_clk new_AGEMA_reg_buffer_8858 ( .C (clk), .D (new_AGEMA_signal_29813), .Q (new_AGEMA_signal_29814) ) ;
    buf_clk new_AGEMA_reg_buffer_8861 ( .C (clk), .D (new_AGEMA_signal_29816), .Q (new_AGEMA_signal_29817) ) ;
    buf_clk new_AGEMA_reg_buffer_8864 ( .C (clk), .D (new_AGEMA_signal_29819), .Q (new_AGEMA_signal_29820) ) ;
    buf_clk new_AGEMA_reg_buffer_8867 ( .C (clk), .D (new_AGEMA_signal_29822), .Q (new_AGEMA_signal_29823) ) ;
    buf_clk new_AGEMA_reg_buffer_8870 ( .C (clk), .D (new_AGEMA_signal_29825), .Q (new_AGEMA_signal_29826) ) ;
    buf_clk new_AGEMA_reg_buffer_8873 ( .C (clk), .D (new_AGEMA_signal_29828), .Q (new_AGEMA_signal_29829) ) ;
    buf_clk new_AGEMA_reg_buffer_8876 ( .C (clk), .D (new_AGEMA_signal_29831), .Q (new_AGEMA_signal_29832) ) ;
    buf_clk new_AGEMA_reg_buffer_8879 ( .C (clk), .D (new_AGEMA_signal_29834), .Q (new_AGEMA_signal_29835) ) ;
    buf_clk new_AGEMA_reg_buffer_8882 ( .C (clk), .D (new_AGEMA_signal_29837), .Q (new_AGEMA_signal_29838) ) ;
    buf_clk new_AGEMA_reg_buffer_8885 ( .C (clk), .D (new_AGEMA_signal_29840), .Q (new_AGEMA_signal_29841) ) ;
    buf_clk new_AGEMA_reg_buffer_8888 ( .C (clk), .D (new_AGEMA_signal_29843), .Q (new_AGEMA_signal_29844) ) ;
    buf_clk new_AGEMA_reg_buffer_8891 ( .C (clk), .D (new_AGEMA_signal_29846), .Q (new_AGEMA_signal_29847) ) ;
    buf_clk new_AGEMA_reg_buffer_8894 ( .C (clk), .D (new_AGEMA_signal_29849), .Q (new_AGEMA_signal_29850) ) ;
    buf_clk new_AGEMA_reg_buffer_8897 ( .C (clk), .D (new_AGEMA_signal_29852), .Q (new_AGEMA_signal_29853) ) ;
    buf_clk new_AGEMA_reg_buffer_8900 ( .C (clk), .D (new_AGEMA_signal_29855), .Q (new_AGEMA_signal_29856) ) ;
    buf_clk new_AGEMA_reg_buffer_8903 ( .C (clk), .D (new_AGEMA_signal_29858), .Q (new_AGEMA_signal_29859) ) ;
    buf_clk new_AGEMA_reg_buffer_8906 ( .C (clk), .D (new_AGEMA_signal_29861), .Q (new_AGEMA_signal_29862) ) ;
    buf_clk new_AGEMA_reg_buffer_8909 ( .C (clk), .D (new_AGEMA_signal_29864), .Q (new_AGEMA_signal_29865) ) ;
    buf_clk new_AGEMA_reg_buffer_8912 ( .C (clk), .D (new_AGEMA_signal_29867), .Q (new_AGEMA_signal_29868) ) ;
    buf_clk new_AGEMA_reg_buffer_8915 ( .C (clk), .D (new_AGEMA_signal_29870), .Q (new_AGEMA_signal_29871) ) ;
    buf_clk new_AGEMA_reg_buffer_8918 ( .C (clk), .D (new_AGEMA_signal_29873), .Q (new_AGEMA_signal_29874) ) ;
    buf_clk new_AGEMA_reg_buffer_8921 ( .C (clk), .D (new_AGEMA_signal_29876), .Q (new_AGEMA_signal_29877) ) ;
    buf_clk new_AGEMA_reg_buffer_8924 ( .C (clk), .D (new_AGEMA_signal_29879), .Q (new_AGEMA_signal_29880) ) ;
    buf_clk new_AGEMA_reg_buffer_8927 ( .C (clk), .D (new_AGEMA_signal_29882), .Q (new_AGEMA_signal_29883) ) ;
    buf_clk new_AGEMA_reg_buffer_8930 ( .C (clk), .D (new_AGEMA_signal_29885), .Q (new_AGEMA_signal_29886) ) ;
    buf_clk new_AGEMA_reg_buffer_8933 ( .C (clk), .D (new_AGEMA_signal_29888), .Q (new_AGEMA_signal_29889) ) ;
    buf_clk new_AGEMA_reg_buffer_8936 ( .C (clk), .D (new_AGEMA_signal_29891), .Q (new_AGEMA_signal_29892) ) ;
    buf_clk new_AGEMA_reg_buffer_8939 ( .C (clk), .D (new_AGEMA_signal_29894), .Q (new_AGEMA_signal_29895) ) ;
    buf_clk new_AGEMA_reg_buffer_8942 ( .C (clk), .D (new_AGEMA_signal_29897), .Q (new_AGEMA_signal_29898) ) ;
    buf_clk new_AGEMA_reg_buffer_8945 ( .C (clk), .D (new_AGEMA_signal_29900), .Q (new_AGEMA_signal_29901) ) ;
    buf_clk new_AGEMA_reg_buffer_8948 ( .C (clk), .D (new_AGEMA_signal_29903), .Q (new_AGEMA_signal_29904) ) ;
    buf_clk new_AGEMA_reg_buffer_8951 ( .C (clk), .D (new_AGEMA_signal_29906), .Q (new_AGEMA_signal_29907) ) ;
    buf_clk new_AGEMA_reg_buffer_8954 ( .C (clk), .D (new_AGEMA_signal_29909), .Q (new_AGEMA_signal_29910) ) ;
    buf_clk new_AGEMA_reg_buffer_8957 ( .C (clk), .D (new_AGEMA_signal_29912), .Q (new_AGEMA_signal_29913) ) ;
    buf_clk new_AGEMA_reg_buffer_8960 ( .C (clk), .D (new_AGEMA_signal_29915), .Q (new_AGEMA_signal_29916) ) ;
    buf_clk new_AGEMA_reg_buffer_8963 ( .C (clk), .D (new_AGEMA_signal_29918), .Q (new_AGEMA_signal_29919) ) ;
    buf_clk new_AGEMA_reg_buffer_8966 ( .C (clk), .D (new_AGEMA_signal_29921), .Q (new_AGEMA_signal_29922) ) ;
    buf_clk new_AGEMA_reg_buffer_8969 ( .C (clk), .D (new_AGEMA_signal_29924), .Q (new_AGEMA_signal_29925) ) ;
    buf_clk new_AGEMA_reg_buffer_8972 ( .C (clk), .D (new_AGEMA_signal_29927), .Q (new_AGEMA_signal_29928) ) ;
    buf_clk new_AGEMA_reg_buffer_8975 ( .C (clk), .D (new_AGEMA_signal_29930), .Q (new_AGEMA_signal_29931) ) ;
    buf_clk new_AGEMA_reg_buffer_8978 ( .C (clk), .D (new_AGEMA_signal_29933), .Q (new_AGEMA_signal_29934) ) ;
    buf_clk new_AGEMA_reg_buffer_8981 ( .C (clk), .D (new_AGEMA_signal_29936), .Q (new_AGEMA_signal_29937) ) ;
    buf_clk new_AGEMA_reg_buffer_8984 ( .C (clk), .D (new_AGEMA_signal_29939), .Q (new_AGEMA_signal_29940) ) ;
    buf_clk new_AGEMA_reg_buffer_8987 ( .C (clk), .D (new_AGEMA_signal_29942), .Q (new_AGEMA_signal_29943) ) ;
    buf_clk new_AGEMA_reg_buffer_8990 ( .C (clk), .D (new_AGEMA_signal_29945), .Q (new_AGEMA_signal_29946) ) ;
    buf_clk new_AGEMA_reg_buffer_8993 ( .C (clk), .D (new_AGEMA_signal_29948), .Q (new_AGEMA_signal_29949) ) ;
    buf_clk new_AGEMA_reg_buffer_8996 ( .C (clk), .D (new_AGEMA_signal_29951), .Q (new_AGEMA_signal_29952) ) ;
    buf_clk new_AGEMA_reg_buffer_8999 ( .C (clk), .D (new_AGEMA_signal_29954), .Q (new_AGEMA_signal_29955) ) ;
    buf_clk new_AGEMA_reg_buffer_9002 ( .C (clk), .D (new_AGEMA_signal_29957), .Q (new_AGEMA_signal_29958) ) ;
    buf_clk new_AGEMA_reg_buffer_9005 ( .C (clk), .D (new_AGEMA_signal_29960), .Q (new_AGEMA_signal_29961) ) ;
    buf_clk new_AGEMA_reg_buffer_9008 ( .C (clk), .D (new_AGEMA_signal_29963), .Q (new_AGEMA_signal_29964) ) ;
    buf_clk new_AGEMA_reg_buffer_9011 ( .C (clk), .D (new_AGEMA_signal_29966), .Q (new_AGEMA_signal_29967) ) ;
    buf_clk new_AGEMA_reg_buffer_9014 ( .C (clk), .D (new_AGEMA_signal_29969), .Q (new_AGEMA_signal_29970) ) ;
    buf_clk new_AGEMA_reg_buffer_9017 ( .C (clk), .D (new_AGEMA_signal_29972), .Q (new_AGEMA_signal_29973) ) ;
    buf_clk new_AGEMA_reg_buffer_9020 ( .C (clk), .D (new_AGEMA_signal_29975), .Q (new_AGEMA_signal_29976) ) ;
    buf_clk new_AGEMA_reg_buffer_9023 ( .C (clk), .D (new_AGEMA_signal_29978), .Q (new_AGEMA_signal_29979) ) ;
    buf_clk new_AGEMA_reg_buffer_9026 ( .C (clk), .D (new_AGEMA_signal_29981), .Q (new_AGEMA_signal_29982) ) ;
    buf_clk new_AGEMA_reg_buffer_9029 ( .C (clk), .D (new_AGEMA_signal_29984), .Q (new_AGEMA_signal_29985) ) ;
    buf_clk new_AGEMA_reg_buffer_9032 ( .C (clk), .D (new_AGEMA_signal_29987), .Q (new_AGEMA_signal_29988) ) ;
    buf_clk new_AGEMA_reg_buffer_9035 ( .C (clk), .D (new_AGEMA_signal_29990), .Q (new_AGEMA_signal_29991) ) ;
    buf_clk new_AGEMA_reg_buffer_9038 ( .C (clk), .D (new_AGEMA_signal_29993), .Q (new_AGEMA_signal_29994) ) ;
    buf_clk new_AGEMA_reg_buffer_9041 ( .C (clk), .D (new_AGEMA_signal_29996), .Q (new_AGEMA_signal_29997) ) ;
    buf_clk new_AGEMA_reg_buffer_9044 ( .C (clk), .D (new_AGEMA_signal_29999), .Q (new_AGEMA_signal_30000) ) ;
    buf_clk new_AGEMA_reg_buffer_9047 ( .C (clk), .D (new_AGEMA_signal_30002), .Q (new_AGEMA_signal_30003) ) ;
    buf_clk new_AGEMA_reg_buffer_9050 ( .C (clk), .D (new_AGEMA_signal_30005), .Q (new_AGEMA_signal_30006) ) ;
    buf_clk new_AGEMA_reg_buffer_9053 ( .C (clk), .D (new_AGEMA_signal_30008), .Q (new_AGEMA_signal_30009) ) ;
    buf_clk new_AGEMA_reg_buffer_9056 ( .C (clk), .D (new_AGEMA_signal_30011), .Q (new_AGEMA_signal_30012) ) ;
    buf_clk new_AGEMA_reg_buffer_9059 ( .C (clk), .D (new_AGEMA_signal_30014), .Q (new_AGEMA_signal_30015) ) ;
    buf_clk new_AGEMA_reg_buffer_9062 ( .C (clk), .D (new_AGEMA_signal_30017), .Q (new_AGEMA_signal_30018) ) ;
    buf_clk new_AGEMA_reg_buffer_9065 ( .C (clk), .D (new_AGEMA_signal_30020), .Q (new_AGEMA_signal_30021) ) ;
    buf_clk new_AGEMA_reg_buffer_9068 ( .C (clk), .D (new_AGEMA_signal_30023), .Q (new_AGEMA_signal_30024) ) ;
    buf_clk new_AGEMA_reg_buffer_9071 ( .C (clk), .D (new_AGEMA_signal_30026), .Q (new_AGEMA_signal_30027) ) ;
    buf_clk new_AGEMA_reg_buffer_9074 ( .C (clk), .D (new_AGEMA_signal_30029), .Q (new_AGEMA_signal_30030) ) ;
    buf_clk new_AGEMA_reg_buffer_9077 ( .C (clk), .D (new_AGEMA_signal_30032), .Q (new_AGEMA_signal_30033) ) ;
    buf_clk new_AGEMA_reg_buffer_9080 ( .C (clk), .D (new_AGEMA_signal_30035), .Q (new_AGEMA_signal_30036) ) ;
    buf_clk new_AGEMA_reg_buffer_9083 ( .C (clk), .D (new_AGEMA_signal_30038), .Q (new_AGEMA_signal_30039) ) ;
    buf_clk new_AGEMA_reg_buffer_9086 ( .C (clk), .D (new_AGEMA_signal_30041), .Q (new_AGEMA_signal_30042) ) ;
    buf_clk new_AGEMA_reg_buffer_9089 ( .C (clk), .D (new_AGEMA_signal_30044), .Q (new_AGEMA_signal_30045) ) ;
    buf_clk new_AGEMA_reg_buffer_9092 ( .C (clk), .D (new_AGEMA_signal_30047), .Q (new_AGEMA_signal_30048) ) ;
    buf_clk new_AGEMA_reg_buffer_9095 ( .C (clk), .D (new_AGEMA_signal_30050), .Q (new_AGEMA_signal_30051) ) ;
    buf_clk new_AGEMA_reg_buffer_9098 ( .C (clk), .D (new_AGEMA_signal_30053), .Q (new_AGEMA_signal_30054) ) ;
    buf_clk new_AGEMA_reg_buffer_9101 ( .C (clk), .D (new_AGEMA_signal_30056), .Q (new_AGEMA_signal_30057) ) ;
    buf_clk new_AGEMA_reg_buffer_9104 ( .C (clk), .D (new_AGEMA_signal_30059), .Q (new_AGEMA_signal_30060) ) ;
    buf_clk new_AGEMA_reg_buffer_9107 ( .C (clk), .D (new_AGEMA_signal_30062), .Q (new_AGEMA_signal_30063) ) ;
    buf_clk new_AGEMA_reg_buffer_9110 ( .C (clk), .D (new_AGEMA_signal_30065), .Q (new_AGEMA_signal_30066) ) ;
    buf_clk new_AGEMA_reg_buffer_9113 ( .C (clk), .D (new_AGEMA_signal_30068), .Q (new_AGEMA_signal_30069) ) ;
    buf_clk new_AGEMA_reg_buffer_9116 ( .C (clk), .D (new_AGEMA_signal_30071), .Q (new_AGEMA_signal_30072) ) ;
    buf_clk new_AGEMA_reg_buffer_9119 ( .C (clk), .D (new_AGEMA_signal_30074), .Q (new_AGEMA_signal_30075) ) ;
    buf_clk new_AGEMA_reg_buffer_9122 ( .C (clk), .D (new_AGEMA_signal_30077), .Q (new_AGEMA_signal_30078) ) ;
    buf_clk new_AGEMA_reg_buffer_9125 ( .C (clk), .D (new_AGEMA_signal_30080), .Q (new_AGEMA_signal_30081) ) ;
    buf_clk new_AGEMA_reg_buffer_9128 ( .C (clk), .D (new_AGEMA_signal_30083), .Q (new_AGEMA_signal_30084) ) ;
    buf_clk new_AGEMA_reg_buffer_9131 ( .C (clk), .D (new_AGEMA_signal_30086), .Q (new_AGEMA_signal_30087) ) ;
    buf_clk new_AGEMA_reg_buffer_9134 ( .C (clk), .D (new_AGEMA_signal_30089), .Q (new_AGEMA_signal_30090) ) ;
    buf_clk new_AGEMA_reg_buffer_9137 ( .C (clk), .D (new_AGEMA_signal_30092), .Q (new_AGEMA_signal_30093) ) ;
    buf_clk new_AGEMA_reg_buffer_9140 ( .C (clk), .D (new_AGEMA_signal_30095), .Q (new_AGEMA_signal_30096) ) ;
    buf_clk new_AGEMA_reg_buffer_9143 ( .C (clk), .D (new_AGEMA_signal_30098), .Q (new_AGEMA_signal_30099) ) ;
    buf_clk new_AGEMA_reg_buffer_9146 ( .C (clk), .D (new_AGEMA_signal_30101), .Q (new_AGEMA_signal_30102) ) ;
    buf_clk new_AGEMA_reg_buffer_9149 ( .C (clk), .D (new_AGEMA_signal_30104), .Q (new_AGEMA_signal_30105) ) ;
    buf_clk new_AGEMA_reg_buffer_9152 ( .C (clk), .D (new_AGEMA_signal_30107), .Q (new_AGEMA_signal_30108) ) ;
    buf_clk new_AGEMA_reg_buffer_9155 ( .C (clk), .D (new_AGEMA_signal_30110), .Q (new_AGEMA_signal_30111) ) ;
    buf_clk new_AGEMA_reg_buffer_9158 ( .C (clk), .D (new_AGEMA_signal_30113), .Q (new_AGEMA_signal_30114) ) ;
    buf_clk new_AGEMA_reg_buffer_9161 ( .C (clk), .D (new_AGEMA_signal_30116), .Q (new_AGEMA_signal_30117) ) ;
    buf_clk new_AGEMA_reg_buffer_9164 ( .C (clk), .D (new_AGEMA_signal_30119), .Q (new_AGEMA_signal_30120) ) ;
    buf_clk new_AGEMA_reg_buffer_9167 ( .C (clk), .D (new_AGEMA_signal_30122), .Q (new_AGEMA_signal_30123) ) ;
    buf_clk new_AGEMA_reg_buffer_9170 ( .C (clk), .D (new_AGEMA_signal_30125), .Q (new_AGEMA_signal_30126) ) ;
    buf_clk new_AGEMA_reg_buffer_9173 ( .C (clk), .D (new_AGEMA_signal_30128), .Q (new_AGEMA_signal_30129) ) ;
    buf_clk new_AGEMA_reg_buffer_9176 ( .C (clk), .D (new_AGEMA_signal_30131), .Q (new_AGEMA_signal_30132) ) ;
    buf_clk new_AGEMA_reg_buffer_9179 ( .C (clk), .D (new_AGEMA_signal_30134), .Q (new_AGEMA_signal_30135) ) ;
    buf_clk new_AGEMA_reg_buffer_9182 ( .C (clk), .D (new_AGEMA_signal_30137), .Q (new_AGEMA_signal_30138) ) ;
    buf_clk new_AGEMA_reg_buffer_9185 ( .C (clk), .D (new_AGEMA_signal_30140), .Q (new_AGEMA_signal_30141) ) ;
    buf_clk new_AGEMA_reg_buffer_9188 ( .C (clk), .D (new_AGEMA_signal_30143), .Q (new_AGEMA_signal_30144) ) ;
    buf_clk new_AGEMA_reg_buffer_9191 ( .C (clk), .D (new_AGEMA_signal_30146), .Q (new_AGEMA_signal_30147) ) ;
    buf_clk new_AGEMA_reg_buffer_9194 ( .C (clk), .D (new_AGEMA_signal_30149), .Q (new_AGEMA_signal_30150) ) ;
    buf_clk new_AGEMA_reg_buffer_9197 ( .C (clk), .D (new_AGEMA_signal_30152), .Q (new_AGEMA_signal_30153) ) ;
    buf_clk new_AGEMA_reg_buffer_9200 ( .C (clk), .D (new_AGEMA_signal_30155), .Q (new_AGEMA_signal_30156) ) ;
    buf_clk new_AGEMA_reg_buffer_9203 ( .C (clk), .D (new_AGEMA_signal_30158), .Q (new_AGEMA_signal_30159) ) ;
    buf_clk new_AGEMA_reg_buffer_9206 ( .C (clk), .D (new_AGEMA_signal_30161), .Q (new_AGEMA_signal_30162) ) ;
    buf_clk new_AGEMA_reg_buffer_9209 ( .C (clk), .D (new_AGEMA_signal_30164), .Q (new_AGEMA_signal_30165) ) ;
    buf_clk new_AGEMA_reg_buffer_9212 ( .C (clk), .D (new_AGEMA_signal_30167), .Q (new_AGEMA_signal_30168) ) ;
    buf_clk new_AGEMA_reg_buffer_9215 ( .C (clk), .D (new_AGEMA_signal_30170), .Q (new_AGEMA_signal_30171) ) ;
    buf_clk new_AGEMA_reg_buffer_9218 ( .C (clk), .D (new_AGEMA_signal_30173), .Q (new_AGEMA_signal_30174) ) ;
    buf_clk new_AGEMA_reg_buffer_9221 ( .C (clk), .D (new_AGEMA_signal_30176), .Q (new_AGEMA_signal_30177) ) ;
    buf_clk new_AGEMA_reg_buffer_9224 ( .C (clk), .D (new_AGEMA_signal_30179), .Q (new_AGEMA_signal_30180) ) ;
    buf_clk new_AGEMA_reg_buffer_9227 ( .C (clk), .D (new_AGEMA_signal_30182), .Q (new_AGEMA_signal_30183) ) ;
    buf_clk new_AGEMA_reg_buffer_9230 ( .C (clk), .D (new_AGEMA_signal_30185), .Q (new_AGEMA_signal_30186) ) ;
    buf_clk new_AGEMA_reg_buffer_9233 ( .C (clk), .D (new_AGEMA_signal_30188), .Q (new_AGEMA_signal_30189) ) ;
    buf_clk new_AGEMA_reg_buffer_9236 ( .C (clk), .D (new_AGEMA_signal_30191), .Q (new_AGEMA_signal_30192) ) ;
    buf_clk new_AGEMA_reg_buffer_9239 ( .C (clk), .D (new_AGEMA_signal_30194), .Q (new_AGEMA_signal_30195) ) ;
    buf_clk new_AGEMA_reg_buffer_9242 ( .C (clk), .D (new_AGEMA_signal_30197), .Q (new_AGEMA_signal_30198) ) ;
    buf_clk new_AGEMA_reg_buffer_9245 ( .C (clk), .D (new_AGEMA_signal_30200), .Q (new_AGEMA_signal_30201) ) ;
    buf_clk new_AGEMA_reg_buffer_9248 ( .C (clk), .D (new_AGEMA_signal_30203), .Q (new_AGEMA_signal_30204) ) ;
    buf_clk new_AGEMA_reg_buffer_9251 ( .C (clk), .D (new_AGEMA_signal_30206), .Q (new_AGEMA_signal_30207) ) ;
    buf_clk new_AGEMA_reg_buffer_9254 ( .C (clk), .D (new_AGEMA_signal_30209), .Q (new_AGEMA_signal_30210) ) ;
    buf_clk new_AGEMA_reg_buffer_9257 ( .C (clk), .D (new_AGEMA_signal_30212), .Q (new_AGEMA_signal_30213) ) ;
    buf_clk new_AGEMA_reg_buffer_9260 ( .C (clk), .D (new_AGEMA_signal_30215), .Q (new_AGEMA_signal_30216) ) ;
    buf_clk new_AGEMA_reg_buffer_9263 ( .C (clk), .D (new_AGEMA_signal_30218), .Q (new_AGEMA_signal_30219) ) ;
    buf_clk new_AGEMA_reg_buffer_9266 ( .C (clk), .D (new_AGEMA_signal_30221), .Q (new_AGEMA_signal_30222) ) ;
    buf_clk new_AGEMA_reg_buffer_9269 ( .C (clk), .D (new_AGEMA_signal_30224), .Q (new_AGEMA_signal_30225) ) ;
    buf_clk new_AGEMA_reg_buffer_9272 ( .C (clk), .D (new_AGEMA_signal_30227), .Q (new_AGEMA_signal_30228) ) ;
    buf_clk new_AGEMA_reg_buffer_9275 ( .C (clk), .D (new_AGEMA_signal_30230), .Q (new_AGEMA_signal_30231) ) ;
    buf_clk new_AGEMA_reg_buffer_9278 ( .C (clk), .D (new_AGEMA_signal_30233), .Q (new_AGEMA_signal_30234) ) ;
    buf_clk new_AGEMA_reg_buffer_9281 ( .C (clk), .D (new_AGEMA_signal_30236), .Q (new_AGEMA_signal_30237) ) ;
    buf_clk new_AGEMA_reg_buffer_9284 ( .C (clk), .D (new_AGEMA_signal_30239), .Q (new_AGEMA_signal_30240) ) ;
    buf_clk new_AGEMA_reg_buffer_9287 ( .C (clk), .D (new_AGEMA_signal_30242), .Q (new_AGEMA_signal_30243) ) ;
    buf_clk new_AGEMA_reg_buffer_9290 ( .C (clk), .D (new_AGEMA_signal_30245), .Q (new_AGEMA_signal_30246) ) ;
    buf_clk new_AGEMA_reg_buffer_9293 ( .C (clk), .D (new_AGEMA_signal_30248), .Q (new_AGEMA_signal_30249) ) ;
    buf_clk new_AGEMA_reg_buffer_9296 ( .C (clk), .D (new_AGEMA_signal_30251), .Q (new_AGEMA_signal_30252) ) ;
    buf_clk new_AGEMA_reg_buffer_9299 ( .C (clk), .D (new_AGEMA_signal_30254), .Q (new_AGEMA_signal_30255) ) ;
    buf_clk new_AGEMA_reg_buffer_9302 ( .C (clk), .D (new_AGEMA_signal_30257), .Q (new_AGEMA_signal_30258) ) ;
    buf_clk new_AGEMA_reg_buffer_9305 ( .C (clk), .D (new_AGEMA_signal_30260), .Q (new_AGEMA_signal_30261) ) ;
    buf_clk new_AGEMA_reg_buffer_9308 ( .C (clk), .D (new_AGEMA_signal_30263), .Q (new_AGEMA_signal_30264) ) ;
    buf_clk new_AGEMA_reg_buffer_9311 ( .C (clk), .D (new_AGEMA_signal_30266), .Q (new_AGEMA_signal_30267) ) ;
    buf_clk new_AGEMA_reg_buffer_9314 ( .C (clk), .D (new_AGEMA_signal_30269), .Q (new_AGEMA_signal_30270) ) ;
    buf_clk new_AGEMA_reg_buffer_9317 ( .C (clk), .D (new_AGEMA_signal_30272), .Q (new_AGEMA_signal_30273) ) ;
    buf_clk new_AGEMA_reg_buffer_9320 ( .C (clk), .D (new_AGEMA_signal_30275), .Q (new_AGEMA_signal_30276) ) ;
    buf_clk new_AGEMA_reg_buffer_9323 ( .C (clk), .D (new_AGEMA_signal_30278), .Q (new_AGEMA_signal_30279) ) ;
    buf_clk new_AGEMA_reg_buffer_9326 ( .C (clk), .D (new_AGEMA_signal_30281), .Q (new_AGEMA_signal_30282) ) ;
    buf_clk new_AGEMA_reg_buffer_9329 ( .C (clk), .D (new_AGEMA_signal_30284), .Q (new_AGEMA_signal_30285) ) ;
    buf_clk new_AGEMA_reg_buffer_9332 ( .C (clk), .D (new_AGEMA_signal_30287), .Q (new_AGEMA_signal_30288) ) ;
    buf_clk new_AGEMA_reg_buffer_9335 ( .C (clk), .D (new_AGEMA_signal_30290), .Q (new_AGEMA_signal_30291) ) ;
    buf_clk new_AGEMA_reg_buffer_9338 ( .C (clk), .D (new_AGEMA_signal_30293), .Q (new_AGEMA_signal_30294) ) ;
    buf_clk new_AGEMA_reg_buffer_9341 ( .C (clk), .D (new_AGEMA_signal_30296), .Q (new_AGEMA_signal_30297) ) ;
    buf_clk new_AGEMA_reg_buffer_9344 ( .C (clk), .D (new_AGEMA_signal_30299), .Q (new_AGEMA_signal_30300) ) ;
    buf_clk new_AGEMA_reg_buffer_9347 ( .C (clk), .D (new_AGEMA_signal_30302), .Q (new_AGEMA_signal_30303) ) ;
    buf_clk new_AGEMA_reg_buffer_9350 ( .C (clk), .D (new_AGEMA_signal_30305), .Q (new_AGEMA_signal_30306) ) ;
    buf_clk new_AGEMA_reg_buffer_9353 ( .C (clk), .D (new_AGEMA_signal_30308), .Q (new_AGEMA_signal_30309) ) ;
    buf_clk new_AGEMA_reg_buffer_9356 ( .C (clk), .D (new_AGEMA_signal_30311), .Q (new_AGEMA_signal_30312) ) ;
    buf_clk new_AGEMA_reg_buffer_9359 ( .C (clk), .D (new_AGEMA_signal_30314), .Q (new_AGEMA_signal_30315) ) ;
    buf_clk new_AGEMA_reg_buffer_9362 ( .C (clk), .D (new_AGEMA_signal_30317), .Q (new_AGEMA_signal_30318) ) ;
    buf_clk new_AGEMA_reg_buffer_9365 ( .C (clk), .D (new_AGEMA_signal_30320), .Q (new_AGEMA_signal_30321) ) ;
    buf_clk new_AGEMA_reg_buffer_9368 ( .C (clk), .D (new_AGEMA_signal_30323), .Q (new_AGEMA_signal_30324) ) ;
    buf_clk new_AGEMA_reg_buffer_9371 ( .C (clk), .D (new_AGEMA_signal_30326), .Q (new_AGEMA_signal_30327) ) ;
    buf_clk new_AGEMA_reg_buffer_9374 ( .C (clk), .D (new_AGEMA_signal_30329), .Q (new_AGEMA_signal_30330) ) ;
    buf_clk new_AGEMA_reg_buffer_9377 ( .C (clk), .D (new_AGEMA_signal_30332), .Q (new_AGEMA_signal_30333) ) ;
    buf_clk new_AGEMA_reg_buffer_9380 ( .C (clk), .D (new_AGEMA_signal_30335), .Q (new_AGEMA_signal_30336) ) ;
    buf_clk new_AGEMA_reg_buffer_9383 ( .C (clk), .D (new_AGEMA_signal_30338), .Q (new_AGEMA_signal_30339) ) ;
    buf_clk new_AGEMA_reg_buffer_9386 ( .C (clk), .D (new_AGEMA_signal_30341), .Q (new_AGEMA_signal_30342) ) ;
    buf_clk new_AGEMA_reg_buffer_9389 ( .C (clk), .D (new_AGEMA_signal_30344), .Q (new_AGEMA_signal_30345) ) ;
    buf_clk new_AGEMA_reg_buffer_9392 ( .C (clk), .D (new_AGEMA_signal_30347), .Q (new_AGEMA_signal_30348) ) ;
    buf_clk new_AGEMA_reg_buffer_9395 ( .C (clk), .D (new_AGEMA_signal_30350), .Q (new_AGEMA_signal_30351) ) ;
    buf_clk new_AGEMA_reg_buffer_9398 ( .C (clk), .D (new_AGEMA_signal_30353), .Q (new_AGEMA_signal_30354) ) ;
    buf_clk new_AGEMA_reg_buffer_9401 ( .C (clk), .D (new_AGEMA_signal_30356), .Q (new_AGEMA_signal_30357) ) ;
    buf_clk new_AGEMA_reg_buffer_9404 ( .C (clk), .D (new_AGEMA_signal_30359), .Q (new_AGEMA_signal_30360) ) ;
    buf_clk new_AGEMA_reg_buffer_9407 ( .C (clk), .D (new_AGEMA_signal_30362), .Q (new_AGEMA_signal_30363) ) ;
    buf_clk new_AGEMA_reg_buffer_9410 ( .C (clk), .D (new_AGEMA_signal_30365), .Q (new_AGEMA_signal_30366) ) ;
    buf_clk new_AGEMA_reg_buffer_9413 ( .C (clk), .D (new_AGEMA_signal_30368), .Q (new_AGEMA_signal_30369) ) ;
    buf_clk new_AGEMA_reg_buffer_9416 ( .C (clk), .D (new_AGEMA_signal_30371), .Q (new_AGEMA_signal_30372) ) ;
    buf_clk new_AGEMA_reg_buffer_9419 ( .C (clk), .D (new_AGEMA_signal_30374), .Q (new_AGEMA_signal_30375) ) ;
    buf_clk new_AGEMA_reg_buffer_9422 ( .C (clk), .D (new_AGEMA_signal_30377), .Q (new_AGEMA_signal_30378) ) ;
    buf_clk new_AGEMA_reg_buffer_9425 ( .C (clk), .D (new_AGEMA_signal_30380), .Q (new_AGEMA_signal_30381) ) ;
    buf_clk new_AGEMA_reg_buffer_9428 ( .C (clk), .D (new_AGEMA_signal_30383), .Q (new_AGEMA_signal_30384) ) ;
    buf_clk new_AGEMA_reg_buffer_9431 ( .C (clk), .D (new_AGEMA_signal_30386), .Q (new_AGEMA_signal_30387) ) ;
    buf_clk new_AGEMA_reg_buffer_9434 ( .C (clk), .D (new_AGEMA_signal_30389), .Q (new_AGEMA_signal_30390) ) ;
    buf_clk new_AGEMA_reg_buffer_9437 ( .C (clk), .D (new_AGEMA_signal_30392), .Q (new_AGEMA_signal_30393) ) ;
    buf_clk new_AGEMA_reg_buffer_9440 ( .C (clk), .D (new_AGEMA_signal_30395), .Q (new_AGEMA_signal_30396) ) ;
    buf_clk new_AGEMA_reg_buffer_9443 ( .C (clk), .D (new_AGEMA_signal_30398), .Q (new_AGEMA_signal_30399) ) ;
    buf_clk new_AGEMA_reg_buffer_9446 ( .C (clk), .D (new_AGEMA_signal_30401), .Q (new_AGEMA_signal_30402) ) ;
    buf_clk new_AGEMA_reg_buffer_9449 ( .C (clk), .D (new_AGEMA_signal_30404), .Q (new_AGEMA_signal_30405) ) ;
    buf_clk new_AGEMA_reg_buffer_9452 ( .C (clk), .D (new_AGEMA_signal_30407), .Q (new_AGEMA_signal_30408) ) ;
    buf_clk new_AGEMA_reg_buffer_9455 ( .C (clk), .D (new_AGEMA_signal_30410), .Q (new_AGEMA_signal_30411) ) ;
    buf_clk new_AGEMA_reg_buffer_9458 ( .C (clk), .D (new_AGEMA_signal_30413), .Q (new_AGEMA_signal_30414) ) ;
    buf_clk new_AGEMA_reg_buffer_9461 ( .C (clk), .D (new_AGEMA_signal_30416), .Q (new_AGEMA_signal_30417) ) ;
    buf_clk new_AGEMA_reg_buffer_9464 ( .C (clk), .D (new_AGEMA_signal_30419), .Q (new_AGEMA_signal_30420) ) ;
    buf_clk new_AGEMA_reg_buffer_9467 ( .C (clk), .D (new_AGEMA_signal_30422), .Q (new_AGEMA_signal_30423) ) ;
    buf_clk new_AGEMA_reg_buffer_9470 ( .C (clk), .D (new_AGEMA_signal_30425), .Q (new_AGEMA_signal_30426) ) ;
    buf_clk new_AGEMA_reg_buffer_9473 ( .C (clk), .D (new_AGEMA_signal_30428), .Q (new_AGEMA_signal_30429) ) ;
    buf_clk new_AGEMA_reg_buffer_9476 ( .C (clk), .D (new_AGEMA_signal_30431), .Q (new_AGEMA_signal_30432) ) ;
    buf_clk new_AGEMA_reg_buffer_9479 ( .C (clk), .D (new_AGEMA_signal_30434), .Q (new_AGEMA_signal_30435) ) ;
    buf_clk new_AGEMA_reg_buffer_9482 ( .C (clk), .D (new_AGEMA_signal_30437), .Q (new_AGEMA_signal_30438) ) ;
    buf_clk new_AGEMA_reg_buffer_9485 ( .C (clk), .D (new_AGEMA_signal_30440), .Q (new_AGEMA_signal_30441) ) ;
    buf_clk new_AGEMA_reg_buffer_9488 ( .C (clk), .D (new_AGEMA_signal_30443), .Q (new_AGEMA_signal_30444) ) ;
    buf_clk new_AGEMA_reg_buffer_9491 ( .C (clk), .D (new_AGEMA_signal_30446), .Q (new_AGEMA_signal_30447) ) ;
    buf_clk new_AGEMA_reg_buffer_9494 ( .C (clk), .D (new_AGEMA_signal_30449), .Q (new_AGEMA_signal_30450) ) ;
    buf_clk new_AGEMA_reg_buffer_9497 ( .C (clk), .D (new_AGEMA_signal_30452), .Q (new_AGEMA_signal_30453) ) ;
    buf_clk new_AGEMA_reg_buffer_9500 ( .C (clk), .D (new_AGEMA_signal_30455), .Q (new_AGEMA_signal_30456) ) ;
    buf_clk new_AGEMA_reg_buffer_9503 ( .C (clk), .D (new_AGEMA_signal_30458), .Q (new_AGEMA_signal_30459) ) ;
    buf_clk new_AGEMA_reg_buffer_9506 ( .C (clk), .D (new_AGEMA_signal_30461), .Q (new_AGEMA_signal_30462) ) ;
    buf_clk new_AGEMA_reg_buffer_9509 ( .C (clk), .D (new_AGEMA_signal_30464), .Q (new_AGEMA_signal_30465) ) ;
    buf_clk new_AGEMA_reg_buffer_9512 ( .C (clk), .D (new_AGEMA_signal_30467), .Q (new_AGEMA_signal_30468) ) ;
    buf_clk new_AGEMA_reg_buffer_9515 ( .C (clk), .D (new_AGEMA_signal_30470), .Q (new_AGEMA_signal_30471) ) ;
    buf_clk new_AGEMA_reg_buffer_9518 ( .C (clk), .D (new_AGEMA_signal_30473), .Q (new_AGEMA_signal_30474) ) ;
    buf_clk new_AGEMA_reg_buffer_9521 ( .C (clk), .D (new_AGEMA_signal_30476), .Q (new_AGEMA_signal_30477) ) ;
    buf_clk new_AGEMA_reg_buffer_9524 ( .C (clk), .D (new_AGEMA_signal_30479), .Q (new_AGEMA_signal_30480) ) ;
    buf_clk new_AGEMA_reg_buffer_9527 ( .C (clk), .D (new_AGEMA_signal_30482), .Q (new_AGEMA_signal_30483) ) ;
    buf_clk new_AGEMA_reg_buffer_9530 ( .C (clk), .D (new_AGEMA_signal_30485), .Q (new_AGEMA_signal_30486) ) ;
    buf_clk new_AGEMA_reg_buffer_9533 ( .C (clk), .D (new_AGEMA_signal_30488), .Q (new_AGEMA_signal_30489) ) ;
    buf_clk new_AGEMA_reg_buffer_9536 ( .C (clk), .D (new_AGEMA_signal_30491), .Q (new_AGEMA_signal_30492) ) ;
    buf_clk new_AGEMA_reg_buffer_9539 ( .C (clk), .D (new_AGEMA_signal_30494), .Q (new_AGEMA_signal_30495) ) ;
    buf_clk new_AGEMA_reg_buffer_9542 ( .C (clk), .D (new_AGEMA_signal_30497), .Q (new_AGEMA_signal_30498) ) ;
    buf_clk new_AGEMA_reg_buffer_9545 ( .C (clk), .D (new_AGEMA_signal_30500), .Q (new_AGEMA_signal_30501) ) ;
    buf_clk new_AGEMA_reg_buffer_9548 ( .C (clk), .D (new_AGEMA_signal_30503), .Q (new_AGEMA_signal_30504) ) ;
    buf_clk new_AGEMA_reg_buffer_9551 ( .C (clk), .D (new_AGEMA_signal_30506), .Q (new_AGEMA_signal_30507) ) ;
    buf_clk new_AGEMA_reg_buffer_9554 ( .C (clk), .D (new_AGEMA_signal_30509), .Q (new_AGEMA_signal_30510) ) ;
    buf_clk new_AGEMA_reg_buffer_9557 ( .C (clk), .D (new_AGEMA_signal_30512), .Q (new_AGEMA_signal_30513) ) ;
    buf_clk new_AGEMA_reg_buffer_9560 ( .C (clk), .D (new_AGEMA_signal_30515), .Q (new_AGEMA_signal_30516) ) ;
    buf_clk new_AGEMA_reg_buffer_9563 ( .C (clk), .D (new_AGEMA_signal_30518), .Q (new_AGEMA_signal_30519) ) ;
    buf_clk new_AGEMA_reg_buffer_9566 ( .C (clk), .D (new_AGEMA_signal_30521), .Q (new_AGEMA_signal_30522) ) ;
    buf_clk new_AGEMA_reg_buffer_9569 ( .C (clk), .D (new_AGEMA_signal_30524), .Q (new_AGEMA_signal_30525) ) ;
    buf_clk new_AGEMA_reg_buffer_9572 ( .C (clk), .D (new_AGEMA_signal_30527), .Q (new_AGEMA_signal_30528) ) ;
    buf_clk new_AGEMA_reg_buffer_9575 ( .C (clk), .D (new_AGEMA_signal_30530), .Q (new_AGEMA_signal_30531) ) ;
    buf_clk new_AGEMA_reg_buffer_9578 ( .C (clk), .D (new_AGEMA_signal_30533), .Q (new_AGEMA_signal_30534) ) ;
    buf_clk new_AGEMA_reg_buffer_9581 ( .C (clk), .D (new_AGEMA_signal_30536), .Q (new_AGEMA_signal_30537) ) ;
    buf_clk new_AGEMA_reg_buffer_9584 ( .C (clk), .D (new_AGEMA_signal_30539), .Q (new_AGEMA_signal_30540) ) ;
    buf_clk new_AGEMA_reg_buffer_9587 ( .C (clk), .D (new_AGEMA_signal_30542), .Q (new_AGEMA_signal_30543) ) ;
    buf_clk new_AGEMA_reg_buffer_9590 ( .C (clk), .D (new_AGEMA_signal_30545), .Q (new_AGEMA_signal_30546) ) ;
    buf_clk new_AGEMA_reg_buffer_9593 ( .C (clk), .D (new_AGEMA_signal_30548), .Q (new_AGEMA_signal_30549) ) ;
    buf_clk new_AGEMA_reg_buffer_9596 ( .C (clk), .D (new_AGEMA_signal_30551), .Q (new_AGEMA_signal_30552) ) ;
    buf_clk new_AGEMA_reg_buffer_9599 ( .C (clk), .D (new_AGEMA_signal_30554), .Q (new_AGEMA_signal_30555) ) ;
    buf_clk new_AGEMA_reg_buffer_9602 ( .C (clk), .D (new_AGEMA_signal_30557), .Q (new_AGEMA_signal_30558) ) ;
    buf_clk new_AGEMA_reg_buffer_9605 ( .C (clk), .D (new_AGEMA_signal_30560), .Q (new_AGEMA_signal_30561) ) ;
    buf_clk new_AGEMA_reg_buffer_9608 ( .C (clk), .D (new_AGEMA_signal_30563), .Q (new_AGEMA_signal_30564) ) ;
    buf_clk new_AGEMA_reg_buffer_9611 ( .C (clk), .D (new_AGEMA_signal_30566), .Q (new_AGEMA_signal_30567) ) ;
    buf_clk new_AGEMA_reg_buffer_9614 ( .C (clk), .D (new_AGEMA_signal_30569), .Q (new_AGEMA_signal_30570) ) ;
    buf_clk new_AGEMA_reg_buffer_9617 ( .C (clk), .D (new_AGEMA_signal_30572), .Q (new_AGEMA_signal_30573) ) ;
    buf_clk new_AGEMA_reg_buffer_9620 ( .C (clk), .D (new_AGEMA_signal_30575), .Q (new_AGEMA_signal_30576) ) ;
    buf_clk new_AGEMA_reg_buffer_9623 ( .C (clk), .D (new_AGEMA_signal_30578), .Q (new_AGEMA_signal_30579) ) ;
    buf_clk new_AGEMA_reg_buffer_9626 ( .C (clk), .D (new_AGEMA_signal_30581), .Q (new_AGEMA_signal_30582) ) ;
    buf_clk new_AGEMA_reg_buffer_9629 ( .C (clk), .D (new_AGEMA_signal_30584), .Q (new_AGEMA_signal_30585) ) ;
    buf_clk new_AGEMA_reg_buffer_9632 ( .C (clk), .D (new_AGEMA_signal_30587), .Q (new_AGEMA_signal_30588) ) ;
    buf_clk new_AGEMA_reg_buffer_9635 ( .C (clk), .D (new_AGEMA_signal_30590), .Q (new_AGEMA_signal_30591) ) ;
    buf_clk new_AGEMA_reg_buffer_9638 ( .C (clk), .D (new_AGEMA_signal_30593), .Q (new_AGEMA_signal_30594) ) ;
    buf_clk new_AGEMA_reg_buffer_9641 ( .C (clk), .D (new_AGEMA_signal_30596), .Q (new_AGEMA_signal_30597) ) ;
    buf_clk new_AGEMA_reg_buffer_9644 ( .C (clk), .D (new_AGEMA_signal_30599), .Q (new_AGEMA_signal_30600) ) ;
    buf_clk new_AGEMA_reg_buffer_9647 ( .C (clk), .D (new_AGEMA_signal_30602), .Q (new_AGEMA_signal_30603) ) ;
    buf_clk new_AGEMA_reg_buffer_9650 ( .C (clk), .D (new_AGEMA_signal_30605), .Q (new_AGEMA_signal_30606) ) ;
    buf_clk new_AGEMA_reg_buffer_9653 ( .C (clk), .D (new_AGEMA_signal_30608), .Q (new_AGEMA_signal_30609) ) ;
    buf_clk new_AGEMA_reg_buffer_9656 ( .C (clk), .D (new_AGEMA_signal_30611), .Q (new_AGEMA_signal_30612) ) ;
    buf_clk new_AGEMA_reg_buffer_9659 ( .C (clk), .D (new_AGEMA_signal_30614), .Q (new_AGEMA_signal_30615) ) ;
    buf_clk new_AGEMA_reg_buffer_9662 ( .C (clk), .D (new_AGEMA_signal_30617), .Q (new_AGEMA_signal_30618) ) ;
    buf_clk new_AGEMA_reg_buffer_9665 ( .C (clk), .D (new_AGEMA_signal_30620), .Q (new_AGEMA_signal_30621) ) ;
    buf_clk new_AGEMA_reg_buffer_9668 ( .C (clk), .D (new_AGEMA_signal_30623), .Q (new_AGEMA_signal_30624) ) ;
    buf_clk new_AGEMA_reg_buffer_9671 ( .C (clk), .D (new_AGEMA_signal_30626), .Q (new_AGEMA_signal_30627) ) ;
    buf_clk new_AGEMA_reg_buffer_9674 ( .C (clk), .D (new_AGEMA_signal_30629), .Q (new_AGEMA_signal_30630) ) ;
    buf_clk new_AGEMA_reg_buffer_9677 ( .C (clk), .D (new_AGEMA_signal_30632), .Q (new_AGEMA_signal_30633) ) ;
    buf_clk new_AGEMA_reg_buffer_9680 ( .C (clk), .D (new_AGEMA_signal_30635), .Q (new_AGEMA_signal_30636) ) ;
    buf_clk new_AGEMA_reg_buffer_9683 ( .C (clk), .D (new_AGEMA_signal_30638), .Q (new_AGEMA_signal_30639) ) ;
    buf_clk new_AGEMA_reg_buffer_9686 ( .C (clk), .D (new_AGEMA_signal_30641), .Q (new_AGEMA_signal_30642) ) ;
    buf_clk new_AGEMA_reg_buffer_9689 ( .C (clk), .D (new_AGEMA_signal_30644), .Q (new_AGEMA_signal_30645) ) ;
    buf_clk new_AGEMA_reg_buffer_9692 ( .C (clk), .D (new_AGEMA_signal_30647), .Q (new_AGEMA_signal_30648) ) ;
    buf_clk new_AGEMA_reg_buffer_9695 ( .C (clk), .D (new_AGEMA_signal_30650), .Q (new_AGEMA_signal_30651) ) ;
    buf_clk new_AGEMA_reg_buffer_9698 ( .C (clk), .D (new_AGEMA_signal_30653), .Q (new_AGEMA_signal_30654) ) ;
    buf_clk new_AGEMA_reg_buffer_9701 ( .C (clk), .D (new_AGEMA_signal_30656), .Q (new_AGEMA_signal_30657) ) ;
    buf_clk new_AGEMA_reg_buffer_9704 ( .C (clk), .D (new_AGEMA_signal_30659), .Q (new_AGEMA_signal_30660) ) ;
    buf_clk new_AGEMA_reg_buffer_9707 ( .C (clk), .D (new_AGEMA_signal_30662), .Q (new_AGEMA_signal_30663) ) ;
    buf_clk new_AGEMA_reg_buffer_9710 ( .C (clk), .D (new_AGEMA_signal_30665), .Q (new_AGEMA_signal_30666) ) ;
    buf_clk new_AGEMA_reg_buffer_9713 ( .C (clk), .D (new_AGEMA_signal_30668), .Q (new_AGEMA_signal_30669) ) ;
    buf_clk new_AGEMA_reg_buffer_9716 ( .C (clk), .D (new_AGEMA_signal_30671), .Q (new_AGEMA_signal_30672) ) ;
    buf_clk new_AGEMA_reg_buffer_9719 ( .C (clk), .D (new_AGEMA_signal_30674), .Q (new_AGEMA_signal_30675) ) ;
    buf_clk new_AGEMA_reg_buffer_9722 ( .C (clk), .D (new_AGEMA_signal_30677), .Q (new_AGEMA_signal_30678) ) ;
    buf_clk new_AGEMA_reg_buffer_9725 ( .C (clk), .D (new_AGEMA_signal_30680), .Q (new_AGEMA_signal_30681) ) ;
    buf_clk new_AGEMA_reg_buffer_9728 ( .C (clk), .D (new_AGEMA_signal_30683), .Q (new_AGEMA_signal_30684) ) ;
    buf_clk new_AGEMA_reg_buffer_9731 ( .C (clk), .D (new_AGEMA_signal_30686), .Q (new_AGEMA_signal_30687) ) ;
    buf_clk new_AGEMA_reg_buffer_9734 ( .C (clk), .D (new_AGEMA_signal_30689), .Q (new_AGEMA_signal_30690) ) ;
    buf_clk new_AGEMA_reg_buffer_9737 ( .C (clk), .D (new_AGEMA_signal_30692), .Q (new_AGEMA_signal_30693) ) ;
    buf_clk new_AGEMA_reg_buffer_9740 ( .C (clk), .D (new_AGEMA_signal_30695), .Q (new_AGEMA_signal_30696) ) ;
    buf_clk new_AGEMA_reg_buffer_9743 ( .C (clk), .D (new_AGEMA_signal_30698), .Q (new_AGEMA_signal_30699) ) ;
    buf_clk new_AGEMA_reg_buffer_9746 ( .C (clk), .D (new_AGEMA_signal_30701), .Q (new_AGEMA_signal_30702) ) ;
    buf_clk new_AGEMA_reg_buffer_9749 ( .C (clk), .D (new_AGEMA_signal_30704), .Q (new_AGEMA_signal_30705) ) ;
    buf_clk new_AGEMA_reg_buffer_9752 ( .C (clk), .D (new_AGEMA_signal_30707), .Q (new_AGEMA_signal_30708) ) ;
    buf_clk new_AGEMA_reg_buffer_9755 ( .C (clk), .D (new_AGEMA_signal_30710), .Q (new_AGEMA_signal_30711) ) ;
    buf_clk new_AGEMA_reg_buffer_9758 ( .C (clk), .D (new_AGEMA_signal_30713), .Q (new_AGEMA_signal_30714) ) ;
    buf_clk new_AGEMA_reg_buffer_9761 ( .C (clk), .D (new_AGEMA_signal_30716), .Q (new_AGEMA_signal_30717) ) ;
    buf_clk new_AGEMA_reg_buffer_9764 ( .C (clk), .D (new_AGEMA_signal_30719), .Q (new_AGEMA_signal_30720) ) ;
    buf_clk new_AGEMA_reg_buffer_9767 ( .C (clk), .D (new_AGEMA_signal_30722), .Q (new_AGEMA_signal_30723) ) ;
    buf_clk new_AGEMA_reg_buffer_9770 ( .C (clk), .D (new_AGEMA_signal_30725), .Q (new_AGEMA_signal_30726) ) ;
    buf_clk new_AGEMA_reg_buffer_9773 ( .C (clk), .D (new_AGEMA_signal_30728), .Q (new_AGEMA_signal_30729) ) ;
    buf_clk new_AGEMA_reg_buffer_9776 ( .C (clk), .D (new_AGEMA_signal_30731), .Q (new_AGEMA_signal_30732) ) ;
    buf_clk new_AGEMA_reg_buffer_9779 ( .C (clk), .D (new_AGEMA_signal_30734), .Q (new_AGEMA_signal_30735) ) ;
    buf_clk new_AGEMA_reg_buffer_9782 ( .C (clk), .D (new_AGEMA_signal_30737), .Q (new_AGEMA_signal_30738) ) ;
    buf_clk new_AGEMA_reg_buffer_9785 ( .C (clk), .D (new_AGEMA_signal_30740), .Q (new_AGEMA_signal_30741) ) ;
    buf_clk new_AGEMA_reg_buffer_9788 ( .C (clk), .D (new_AGEMA_signal_30743), .Q (new_AGEMA_signal_30744) ) ;
    buf_clk new_AGEMA_reg_buffer_9791 ( .C (clk), .D (new_AGEMA_signal_30746), .Q (new_AGEMA_signal_30747) ) ;
    buf_clk new_AGEMA_reg_buffer_9794 ( .C (clk), .D (new_AGEMA_signal_30749), .Q (new_AGEMA_signal_30750) ) ;
    buf_clk new_AGEMA_reg_buffer_9797 ( .C (clk), .D (new_AGEMA_signal_30752), .Q (new_AGEMA_signal_30753) ) ;
    buf_clk new_AGEMA_reg_buffer_9800 ( .C (clk), .D (new_AGEMA_signal_30755), .Q (new_AGEMA_signal_30756) ) ;
    buf_clk new_AGEMA_reg_buffer_9803 ( .C (clk), .D (new_AGEMA_signal_30758), .Q (new_AGEMA_signal_30759) ) ;
    buf_clk new_AGEMA_reg_buffer_9806 ( .C (clk), .D (new_AGEMA_signal_30761), .Q (new_AGEMA_signal_30762) ) ;
    buf_clk new_AGEMA_reg_buffer_9809 ( .C (clk), .D (new_AGEMA_signal_30764), .Q (new_AGEMA_signal_30765) ) ;
    buf_clk new_AGEMA_reg_buffer_9812 ( .C (clk), .D (new_AGEMA_signal_30767), .Q (new_AGEMA_signal_30768) ) ;
    buf_clk new_AGEMA_reg_buffer_9815 ( .C (clk), .D (new_AGEMA_signal_30770), .Q (new_AGEMA_signal_30771) ) ;
    buf_clk new_AGEMA_reg_buffer_9818 ( .C (clk), .D (new_AGEMA_signal_30773), .Q (new_AGEMA_signal_30774) ) ;
    buf_clk new_AGEMA_reg_buffer_9821 ( .C (clk), .D (new_AGEMA_signal_30776), .Q (new_AGEMA_signal_30777) ) ;
    buf_clk new_AGEMA_reg_buffer_9824 ( .C (clk), .D (new_AGEMA_signal_30779), .Q (new_AGEMA_signal_30780) ) ;
    buf_clk new_AGEMA_reg_buffer_9827 ( .C (clk), .D (new_AGEMA_signal_30782), .Q (new_AGEMA_signal_30783) ) ;
    buf_clk new_AGEMA_reg_buffer_9830 ( .C (clk), .D (new_AGEMA_signal_30785), .Q (new_AGEMA_signal_30786) ) ;
    buf_clk new_AGEMA_reg_buffer_9833 ( .C (clk), .D (new_AGEMA_signal_30788), .Q (new_AGEMA_signal_30789) ) ;
    buf_clk new_AGEMA_reg_buffer_9836 ( .C (clk), .D (new_AGEMA_signal_30791), .Q (new_AGEMA_signal_30792) ) ;
    buf_clk new_AGEMA_reg_buffer_9839 ( .C (clk), .D (new_AGEMA_signal_30794), .Q (new_AGEMA_signal_30795) ) ;
    buf_clk new_AGEMA_reg_buffer_9842 ( .C (clk), .D (new_AGEMA_signal_30797), .Q (new_AGEMA_signal_30798) ) ;
    buf_clk new_AGEMA_reg_buffer_9845 ( .C (clk), .D (new_AGEMA_signal_30800), .Q (new_AGEMA_signal_30801) ) ;
    buf_clk new_AGEMA_reg_buffer_9848 ( .C (clk), .D (new_AGEMA_signal_30803), .Q (new_AGEMA_signal_30804) ) ;
    buf_clk new_AGEMA_reg_buffer_9851 ( .C (clk), .D (new_AGEMA_signal_30806), .Q (new_AGEMA_signal_30807) ) ;
    buf_clk new_AGEMA_reg_buffer_9854 ( .C (clk), .D (new_AGEMA_signal_30809), .Q (new_AGEMA_signal_30810) ) ;
    buf_clk new_AGEMA_reg_buffer_9857 ( .C (clk), .D (new_AGEMA_signal_30812), .Q (new_AGEMA_signal_30813) ) ;
    buf_clk new_AGEMA_reg_buffer_9860 ( .C (clk), .D (new_AGEMA_signal_30815), .Q (new_AGEMA_signal_30816) ) ;
    buf_clk new_AGEMA_reg_buffer_9863 ( .C (clk), .D (new_AGEMA_signal_30818), .Q (new_AGEMA_signal_30819) ) ;
    buf_clk new_AGEMA_reg_buffer_9866 ( .C (clk), .D (new_AGEMA_signal_30821), .Q (new_AGEMA_signal_30822) ) ;
    buf_clk new_AGEMA_reg_buffer_9869 ( .C (clk), .D (new_AGEMA_signal_30824), .Q (new_AGEMA_signal_30825) ) ;
    buf_clk new_AGEMA_reg_buffer_9872 ( .C (clk), .D (new_AGEMA_signal_30827), .Q (new_AGEMA_signal_30828) ) ;
    buf_clk new_AGEMA_reg_buffer_9875 ( .C (clk), .D (new_AGEMA_signal_30830), .Q (new_AGEMA_signal_30831) ) ;
    buf_clk new_AGEMA_reg_buffer_9878 ( .C (clk), .D (new_AGEMA_signal_30833), .Q (new_AGEMA_signal_30834) ) ;
    buf_clk new_AGEMA_reg_buffer_9881 ( .C (clk), .D (new_AGEMA_signal_30836), .Q (new_AGEMA_signal_30837) ) ;
    buf_clk new_AGEMA_reg_buffer_9884 ( .C (clk), .D (new_AGEMA_signal_30839), .Q (new_AGEMA_signal_30840) ) ;
    buf_clk new_AGEMA_reg_buffer_9887 ( .C (clk), .D (new_AGEMA_signal_30842), .Q (new_AGEMA_signal_30843) ) ;
    buf_clk new_AGEMA_reg_buffer_9890 ( .C (clk), .D (new_AGEMA_signal_30845), .Q (new_AGEMA_signal_30846) ) ;
    buf_clk new_AGEMA_reg_buffer_9893 ( .C (clk), .D (new_AGEMA_signal_30848), .Q (new_AGEMA_signal_30849) ) ;
    buf_clk new_AGEMA_reg_buffer_9896 ( .C (clk), .D (new_AGEMA_signal_30851), .Q (new_AGEMA_signal_30852) ) ;
    buf_clk new_AGEMA_reg_buffer_9899 ( .C (clk), .D (new_AGEMA_signal_30854), .Q (new_AGEMA_signal_30855) ) ;
    buf_clk new_AGEMA_reg_buffer_9902 ( .C (clk), .D (new_AGEMA_signal_30857), .Q (new_AGEMA_signal_30858) ) ;
    buf_clk new_AGEMA_reg_buffer_9905 ( .C (clk), .D (new_AGEMA_signal_30860), .Q (new_AGEMA_signal_30861) ) ;
    buf_clk new_AGEMA_reg_buffer_9908 ( .C (clk), .D (new_AGEMA_signal_30863), .Q (new_AGEMA_signal_30864) ) ;
    buf_clk new_AGEMA_reg_buffer_9911 ( .C (clk), .D (new_AGEMA_signal_30866), .Q (new_AGEMA_signal_30867) ) ;
    buf_clk new_AGEMA_reg_buffer_9914 ( .C (clk), .D (new_AGEMA_signal_30869), .Q (new_AGEMA_signal_30870) ) ;
    buf_clk new_AGEMA_reg_buffer_9917 ( .C (clk), .D (new_AGEMA_signal_30872), .Q (new_AGEMA_signal_30873) ) ;
    buf_clk new_AGEMA_reg_buffer_9920 ( .C (clk), .D (new_AGEMA_signal_30875), .Q (new_AGEMA_signal_30876) ) ;
    buf_clk new_AGEMA_reg_buffer_9923 ( .C (clk), .D (new_AGEMA_signal_30878), .Q (new_AGEMA_signal_30879) ) ;
    buf_clk new_AGEMA_reg_buffer_9926 ( .C (clk), .D (new_AGEMA_signal_30881), .Q (new_AGEMA_signal_30882) ) ;
    buf_clk new_AGEMA_reg_buffer_9929 ( .C (clk), .D (new_AGEMA_signal_30884), .Q (new_AGEMA_signal_30885) ) ;
    buf_clk new_AGEMA_reg_buffer_9932 ( .C (clk), .D (new_AGEMA_signal_30887), .Q (new_AGEMA_signal_30888) ) ;
    buf_clk new_AGEMA_reg_buffer_9935 ( .C (clk), .D (new_AGEMA_signal_30890), .Q (new_AGEMA_signal_30891) ) ;
    buf_clk new_AGEMA_reg_buffer_9938 ( .C (clk), .D (new_AGEMA_signal_30893), .Q (new_AGEMA_signal_30894) ) ;
    buf_clk new_AGEMA_reg_buffer_9941 ( .C (clk), .D (new_AGEMA_signal_30896), .Q (new_AGEMA_signal_30897) ) ;
    buf_clk new_AGEMA_reg_buffer_9944 ( .C (clk), .D (new_AGEMA_signal_30899), .Q (new_AGEMA_signal_30900) ) ;
    buf_clk new_AGEMA_reg_buffer_9947 ( .C (clk), .D (new_AGEMA_signal_30902), .Q (new_AGEMA_signal_30903) ) ;
    buf_clk new_AGEMA_reg_buffer_9950 ( .C (clk), .D (new_AGEMA_signal_30905), .Q (new_AGEMA_signal_30906) ) ;
    buf_clk new_AGEMA_reg_buffer_9953 ( .C (clk), .D (new_AGEMA_signal_30908), .Q (new_AGEMA_signal_30909) ) ;
    buf_clk new_AGEMA_reg_buffer_9956 ( .C (clk), .D (new_AGEMA_signal_30911), .Q (new_AGEMA_signal_30912) ) ;
    buf_clk new_AGEMA_reg_buffer_9959 ( .C (clk), .D (new_AGEMA_signal_30914), .Q (new_AGEMA_signal_30915) ) ;
    buf_clk new_AGEMA_reg_buffer_9962 ( .C (clk), .D (new_AGEMA_signal_30917), .Q (new_AGEMA_signal_30918) ) ;
    buf_clk new_AGEMA_reg_buffer_9965 ( .C (clk), .D (new_AGEMA_signal_30920), .Q (new_AGEMA_signal_30921) ) ;
    buf_clk new_AGEMA_reg_buffer_9968 ( .C (clk), .D (new_AGEMA_signal_30923), .Q (new_AGEMA_signal_30924) ) ;
    buf_clk new_AGEMA_reg_buffer_9971 ( .C (clk), .D (new_AGEMA_signal_30926), .Q (new_AGEMA_signal_30927) ) ;
    buf_clk new_AGEMA_reg_buffer_9974 ( .C (clk), .D (new_AGEMA_signal_30929), .Q (new_AGEMA_signal_30930) ) ;
    buf_clk new_AGEMA_reg_buffer_9977 ( .C (clk), .D (new_AGEMA_signal_30932), .Q (new_AGEMA_signal_30933) ) ;
    buf_clk new_AGEMA_reg_buffer_9980 ( .C (clk), .D (new_AGEMA_signal_30935), .Q (new_AGEMA_signal_30936) ) ;
    buf_clk new_AGEMA_reg_buffer_9983 ( .C (clk), .D (new_AGEMA_signal_30938), .Q (new_AGEMA_signal_30939) ) ;
    buf_clk new_AGEMA_reg_buffer_9986 ( .C (clk), .D (new_AGEMA_signal_30941), .Q (new_AGEMA_signal_30942) ) ;
    buf_clk new_AGEMA_reg_buffer_9989 ( .C (clk), .D (new_AGEMA_signal_30944), .Q (new_AGEMA_signal_30945) ) ;
    buf_clk new_AGEMA_reg_buffer_9992 ( .C (clk), .D (new_AGEMA_signal_30947), .Q (new_AGEMA_signal_30948) ) ;
    buf_clk new_AGEMA_reg_buffer_9995 ( .C (clk), .D (new_AGEMA_signal_30950), .Q (new_AGEMA_signal_30951) ) ;
    buf_clk new_AGEMA_reg_buffer_9998 ( .C (clk), .D (new_AGEMA_signal_30953), .Q (new_AGEMA_signal_30954) ) ;
    buf_clk new_AGEMA_reg_buffer_10001 ( .C (clk), .D (new_AGEMA_signal_30956), .Q (new_AGEMA_signal_30957) ) ;
    buf_clk new_AGEMA_reg_buffer_10004 ( .C (clk), .D (new_AGEMA_signal_30959), .Q (new_AGEMA_signal_30960) ) ;
    buf_clk new_AGEMA_reg_buffer_10007 ( .C (clk), .D (new_AGEMA_signal_30962), .Q (new_AGEMA_signal_30963) ) ;
    buf_clk new_AGEMA_reg_buffer_10010 ( .C (clk), .D (new_AGEMA_signal_30965), .Q (new_AGEMA_signal_30966) ) ;
    buf_clk new_AGEMA_reg_buffer_10013 ( .C (clk), .D (new_AGEMA_signal_30968), .Q (new_AGEMA_signal_30969) ) ;
    buf_clk new_AGEMA_reg_buffer_10016 ( .C (clk), .D (new_AGEMA_signal_30971), .Q (new_AGEMA_signal_30972) ) ;
    buf_clk new_AGEMA_reg_buffer_10019 ( .C (clk), .D (new_AGEMA_signal_30974), .Q (new_AGEMA_signal_30975) ) ;
    buf_clk new_AGEMA_reg_buffer_10022 ( .C (clk), .D (new_AGEMA_signal_30977), .Q (new_AGEMA_signal_30978) ) ;
    buf_clk new_AGEMA_reg_buffer_10025 ( .C (clk), .D (new_AGEMA_signal_30980), .Q (new_AGEMA_signal_30981) ) ;
    buf_clk new_AGEMA_reg_buffer_10028 ( .C (clk), .D (new_AGEMA_signal_30983), .Q (new_AGEMA_signal_30984) ) ;
    buf_clk new_AGEMA_reg_buffer_10031 ( .C (clk), .D (new_AGEMA_signal_30986), .Q (new_AGEMA_signal_30987) ) ;
    buf_clk new_AGEMA_reg_buffer_10034 ( .C (clk), .D (new_AGEMA_signal_30989), .Q (new_AGEMA_signal_30990) ) ;
    buf_clk new_AGEMA_reg_buffer_10037 ( .C (clk), .D (new_AGEMA_signal_30992), .Q (new_AGEMA_signal_30993) ) ;
    buf_clk new_AGEMA_reg_buffer_10040 ( .C (clk), .D (new_AGEMA_signal_30995), .Q (new_AGEMA_signal_30996) ) ;
    buf_clk new_AGEMA_reg_buffer_10043 ( .C (clk), .D (new_AGEMA_signal_30998), .Q (new_AGEMA_signal_30999) ) ;
    buf_clk new_AGEMA_reg_buffer_10046 ( .C (clk), .D (new_AGEMA_signal_31001), .Q (new_AGEMA_signal_31002) ) ;
    buf_clk new_AGEMA_reg_buffer_10049 ( .C (clk), .D (new_AGEMA_signal_31004), .Q (new_AGEMA_signal_31005) ) ;
    buf_clk new_AGEMA_reg_buffer_10052 ( .C (clk), .D (new_AGEMA_signal_31007), .Q (new_AGEMA_signal_31008) ) ;
    buf_clk new_AGEMA_reg_buffer_10055 ( .C (clk), .D (new_AGEMA_signal_31010), .Q (new_AGEMA_signal_31011) ) ;
    buf_clk new_AGEMA_reg_buffer_10058 ( .C (clk), .D (new_AGEMA_signal_31013), .Q (new_AGEMA_signal_31014) ) ;
    buf_clk new_AGEMA_reg_buffer_10061 ( .C (clk), .D (new_AGEMA_signal_31016), .Q (new_AGEMA_signal_31017) ) ;
    buf_clk new_AGEMA_reg_buffer_10064 ( .C (clk), .D (new_AGEMA_signal_31019), .Q (new_AGEMA_signal_31020) ) ;
    buf_clk new_AGEMA_reg_buffer_10067 ( .C (clk), .D (new_AGEMA_signal_31022), .Q (new_AGEMA_signal_31023) ) ;
    buf_clk new_AGEMA_reg_buffer_10070 ( .C (clk), .D (new_AGEMA_signal_31025), .Q (new_AGEMA_signal_31026) ) ;
    buf_clk new_AGEMA_reg_buffer_10073 ( .C (clk), .D (new_AGEMA_signal_31028), .Q (new_AGEMA_signal_31029) ) ;
    buf_clk new_AGEMA_reg_buffer_10076 ( .C (clk), .D (new_AGEMA_signal_31031), .Q (new_AGEMA_signal_31032) ) ;
    buf_clk new_AGEMA_reg_buffer_10079 ( .C (clk), .D (new_AGEMA_signal_31034), .Q (new_AGEMA_signal_31035) ) ;
    buf_clk new_AGEMA_reg_buffer_10082 ( .C (clk), .D (new_AGEMA_signal_31037), .Q (new_AGEMA_signal_31038) ) ;
    buf_clk new_AGEMA_reg_buffer_10085 ( .C (clk), .D (new_AGEMA_signal_31040), .Q (new_AGEMA_signal_31041) ) ;
    buf_clk new_AGEMA_reg_buffer_10088 ( .C (clk), .D (new_AGEMA_signal_31043), .Q (new_AGEMA_signal_31044) ) ;
    buf_clk new_AGEMA_reg_buffer_10091 ( .C (clk), .D (new_AGEMA_signal_31046), .Q (new_AGEMA_signal_31047) ) ;
    buf_clk new_AGEMA_reg_buffer_10094 ( .C (clk), .D (new_AGEMA_signal_31049), .Q (new_AGEMA_signal_31050) ) ;
    buf_clk new_AGEMA_reg_buffer_10097 ( .C (clk), .D (new_AGEMA_signal_31052), .Q (new_AGEMA_signal_31053) ) ;
    buf_clk new_AGEMA_reg_buffer_10100 ( .C (clk), .D (new_AGEMA_signal_31055), .Q (new_AGEMA_signal_31056) ) ;
    buf_clk new_AGEMA_reg_buffer_10103 ( .C (clk), .D (new_AGEMA_signal_31058), .Q (new_AGEMA_signal_31059) ) ;
    buf_clk new_AGEMA_reg_buffer_10106 ( .C (clk), .D (new_AGEMA_signal_31061), .Q (new_AGEMA_signal_31062) ) ;
    buf_clk new_AGEMA_reg_buffer_10109 ( .C (clk), .D (new_AGEMA_signal_31064), .Q (new_AGEMA_signal_31065) ) ;
    buf_clk new_AGEMA_reg_buffer_10112 ( .C (clk), .D (new_AGEMA_signal_31067), .Q (new_AGEMA_signal_31068) ) ;
    buf_clk new_AGEMA_reg_buffer_10115 ( .C (clk), .D (new_AGEMA_signal_31070), .Q (new_AGEMA_signal_31071) ) ;
    buf_clk new_AGEMA_reg_buffer_10118 ( .C (clk), .D (new_AGEMA_signal_31073), .Q (new_AGEMA_signal_31074) ) ;
    buf_clk new_AGEMA_reg_buffer_10121 ( .C (clk), .D (new_AGEMA_signal_31076), .Q (new_AGEMA_signal_31077) ) ;
    buf_clk new_AGEMA_reg_buffer_10124 ( .C (clk), .D (new_AGEMA_signal_31079), .Q (new_AGEMA_signal_31080) ) ;
    buf_clk new_AGEMA_reg_buffer_10127 ( .C (clk), .D (new_AGEMA_signal_31082), .Q (new_AGEMA_signal_31083) ) ;
    buf_clk new_AGEMA_reg_buffer_10130 ( .C (clk), .D (new_AGEMA_signal_31085), .Q (new_AGEMA_signal_31086) ) ;
    buf_clk new_AGEMA_reg_buffer_10133 ( .C (clk), .D (new_AGEMA_signal_31088), .Q (new_AGEMA_signal_31089) ) ;
    buf_clk new_AGEMA_reg_buffer_10136 ( .C (clk), .D (new_AGEMA_signal_31091), .Q (new_AGEMA_signal_31092) ) ;
    buf_clk new_AGEMA_reg_buffer_10139 ( .C (clk), .D (new_AGEMA_signal_31094), .Q (new_AGEMA_signal_31095) ) ;
    buf_clk new_AGEMA_reg_buffer_10142 ( .C (clk), .D (new_AGEMA_signal_31097), .Q (new_AGEMA_signal_31098) ) ;
    buf_clk new_AGEMA_reg_buffer_10145 ( .C (clk), .D (new_AGEMA_signal_31100), .Q (new_AGEMA_signal_31101) ) ;
    buf_clk new_AGEMA_reg_buffer_10148 ( .C (clk), .D (new_AGEMA_signal_31103), .Q (new_AGEMA_signal_31104) ) ;
    buf_clk new_AGEMA_reg_buffer_10151 ( .C (clk), .D (new_AGEMA_signal_31106), .Q (new_AGEMA_signal_31107) ) ;
    buf_clk new_AGEMA_reg_buffer_10154 ( .C (clk), .D (new_AGEMA_signal_31109), .Q (new_AGEMA_signal_31110) ) ;
    buf_clk new_AGEMA_reg_buffer_10157 ( .C (clk), .D (new_AGEMA_signal_31112), .Q (new_AGEMA_signal_31113) ) ;
    buf_clk new_AGEMA_reg_buffer_10160 ( .C (clk), .D (new_AGEMA_signal_31115), .Q (new_AGEMA_signal_31116) ) ;
    buf_clk new_AGEMA_reg_buffer_10163 ( .C (clk), .D (new_AGEMA_signal_31118), .Q (new_AGEMA_signal_31119) ) ;
    buf_clk new_AGEMA_reg_buffer_10166 ( .C (clk), .D (new_AGEMA_signal_31121), .Q (new_AGEMA_signal_31122) ) ;
    buf_clk new_AGEMA_reg_buffer_10169 ( .C (clk), .D (new_AGEMA_signal_31124), .Q (new_AGEMA_signal_31125) ) ;
    buf_clk new_AGEMA_reg_buffer_10172 ( .C (clk), .D (new_AGEMA_signal_31127), .Q (new_AGEMA_signal_31128) ) ;
    buf_clk new_AGEMA_reg_buffer_10175 ( .C (clk), .D (new_AGEMA_signal_31130), .Q (new_AGEMA_signal_31131) ) ;
    buf_clk new_AGEMA_reg_buffer_10178 ( .C (clk), .D (new_AGEMA_signal_31133), .Q (new_AGEMA_signal_31134) ) ;
    buf_clk new_AGEMA_reg_buffer_10181 ( .C (clk), .D (new_AGEMA_signal_31136), .Q (new_AGEMA_signal_31137) ) ;
    buf_clk new_AGEMA_reg_buffer_10184 ( .C (clk), .D (new_AGEMA_signal_31139), .Q (new_AGEMA_signal_31140) ) ;
    buf_clk new_AGEMA_reg_buffer_10187 ( .C (clk), .D (new_AGEMA_signal_31142), .Q (new_AGEMA_signal_31143) ) ;
    buf_clk new_AGEMA_reg_buffer_10190 ( .C (clk), .D (new_AGEMA_signal_31145), .Q (new_AGEMA_signal_31146) ) ;
    buf_clk new_AGEMA_reg_buffer_10193 ( .C (clk), .D (new_AGEMA_signal_31148), .Q (new_AGEMA_signal_31149) ) ;
    buf_clk new_AGEMA_reg_buffer_10196 ( .C (clk), .D (new_AGEMA_signal_31151), .Q (new_AGEMA_signal_31152) ) ;
    buf_clk new_AGEMA_reg_buffer_10199 ( .C (clk), .D (new_AGEMA_signal_31154), .Q (new_AGEMA_signal_31155) ) ;
    buf_clk new_AGEMA_reg_buffer_10202 ( .C (clk), .D (new_AGEMA_signal_31157), .Q (new_AGEMA_signal_31158) ) ;
    buf_clk new_AGEMA_reg_buffer_10205 ( .C (clk), .D (new_AGEMA_signal_31160), .Q (new_AGEMA_signal_31161) ) ;
    buf_clk new_AGEMA_reg_buffer_10208 ( .C (clk), .D (new_AGEMA_signal_31163), .Q (new_AGEMA_signal_31164) ) ;
    buf_clk new_AGEMA_reg_buffer_10211 ( .C (clk), .D (new_AGEMA_signal_31166), .Q (new_AGEMA_signal_31167) ) ;
    buf_clk new_AGEMA_reg_buffer_10214 ( .C (clk), .D (new_AGEMA_signal_31169), .Q (new_AGEMA_signal_31170) ) ;
    buf_clk new_AGEMA_reg_buffer_10217 ( .C (clk), .D (new_AGEMA_signal_31172), .Q (new_AGEMA_signal_31173) ) ;
    buf_clk new_AGEMA_reg_buffer_10220 ( .C (clk), .D (new_AGEMA_signal_31175), .Q (new_AGEMA_signal_31176) ) ;
    buf_clk new_AGEMA_reg_buffer_10223 ( .C (clk), .D (new_AGEMA_signal_31178), .Q (new_AGEMA_signal_31179) ) ;
    buf_clk new_AGEMA_reg_buffer_10226 ( .C (clk), .D (new_AGEMA_signal_31181), .Q (new_AGEMA_signal_31182) ) ;
    buf_clk new_AGEMA_reg_buffer_10229 ( .C (clk), .D (new_AGEMA_signal_31184), .Q (new_AGEMA_signal_31185) ) ;
    buf_clk new_AGEMA_reg_buffer_10232 ( .C (clk), .D (new_AGEMA_signal_31187), .Q (new_AGEMA_signal_31188) ) ;
    buf_clk new_AGEMA_reg_buffer_10235 ( .C (clk), .D (new_AGEMA_signal_31190), .Q (new_AGEMA_signal_31191) ) ;
    buf_clk new_AGEMA_reg_buffer_10238 ( .C (clk), .D (new_AGEMA_signal_31193), .Q (new_AGEMA_signal_31194) ) ;
    buf_clk new_AGEMA_reg_buffer_10241 ( .C (clk), .D (new_AGEMA_signal_31196), .Q (new_AGEMA_signal_31197) ) ;
    buf_clk new_AGEMA_reg_buffer_10244 ( .C (clk), .D (new_AGEMA_signal_31199), .Q (new_AGEMA_signal_31200) ) ;
    buf_clk new_AGEMA_reg_buffer_10247 ( .C (clk), .D (new_AGEMA_signal_31202), .Q (new_AGEMA_signal_31203) ) ;
    buf_clk new_AGEMA_reg_buffer_10250 ( .C (clk), .D (new_AGEMA_signal_31205), .Q (new_AGEMA_signal_31206) ) ;
    buf_clk new_AGEMA_reg_buffer_10253 ( .C (clk), .D (new_AGEMA_signal_31208), .Q (new_AGEMA_signal_31209) ) ;
    buf_clk new_AGEMA_reg_buffer_10256 ( .C (clk), .D (new_AGEMA_signal_31211), .Q (new_AGEMA_signal_31212) ) ;
    buf_clk new_AGEMA_reg_buffer_10259 ( .C (clk), .D (new_AGEMA_signal_31214), .Q (new_AGEMA_signal_31215) ) ;
    buf_clk new_AGEMA_reg_buffer_10262 ( .C (clk), .D (new_AGEMA_signal_31217), .Q (new_AGEMA_signal_31218) ) ;
    buf_clk new_AGEMA_reg_buffer_10265 ( .C (clk), .D (new_AGEMA_signal_31220), .Q (new_AGEMA_signal_31221) ) ;
    buf_clk new_AGEMA_reg_buffer_10268 ( .C (clk), .D (new_AGEMA_signal_31223), .Q (new_AGEMA_signal_31224) ) ;
    buf_clk new_AGEMA_reg_buffer_10271 ( .C (clk), .D (new_AGEMA_signal_31226), .Q (new_AGEMA_signal_31227) ) ;
    buf_clk new_AGEMA_reg_buffer_10274 ( .C (clk), .D (new_AGEMA_signal_31229), .Q (new_AGEMA_signal_31230) ) ;
    buf_clk new_AGEMA_reg_buffer_10277 ( .C (clk), .D (new_AGEMA_signal_31232), .Q (new_AGEMA_signal_31233) ) ;
    buf_clk new_AGEMA_reg_buffer_10280 ( .C (clk), .D (new_AGEMA_signal_31235), .Q (new_AGEMA_signal_31236) ) ;
    buf_clk new_AGEMA_reg_buffer_10283 ( .C (clk), .D (new_AGEMA_signal_31238), .Q (new_AGEMA_signal_31239) ) ;
    buf_clk new_AGEMA_reg_buffer_10286 ( .C (clk), .D (new_AGEMA_signal_31241), .Q (new_AGEMA_signal_31242) ) ;
    buf_clk new_AGEMA_reg_buffer_10289 ( .C (clk), .D (new_AGEMA_signal_31244), .Q (new_AGEMA_signal_31245) ) ;
    buf_clk new_AGEMA_reg_buffer_10292 ( .C (clk), .D (new_AGEMA_signal_31247), .Q (new_AGEMA_signal_31248) ) ;
    buf_clk new_AGEMA_reg_buffer_10295 ( .C (clk), .D (new_AGEMA_signal_31250), .Q (new_AGEMA_signal_31251) ) ;
    buf_clk new_AGEMA_reg_buffer_10298 ( .C (clk), .D (new_AGEMA_signal_31253), .Q (new_AGEMA_signal_31254) ) ;
    buf_clk new_AGEMA_reg_buffer_10301 ( .C (clk), .D (new_AGEMA_signal_31256), .Q (new_AGEMA_signal_31257) ) ;
    buf_clk new_AGEMA_reg_buffer_10304 ( .C (clk), .D (new_AGEMA_signal_31259), .Q (new_AGEMA_signal_31260) ) ;
    buf_clk new_AGEMA_reg_buffer_10307 ( .C (clk), .D (new_AGEMA_signal_31262), .Q (new_AGEMA_signal_31263) ) ;
    buf_clk new_AGEMA_reg_buffer_10310 ( .C (clk), .D (new_AGEMA_signal_31265), .Q (new_AGEMA_signal_31266) ) ;
    buf_clk new_AGEMA_reg_buffer_10313 ( .C (clk), .D (new_AGEMA_signal_31268), .Q (new_AGEMA_signal_31269) ) ;
    buf_clk new_AGEMA_reg_buffer_10316 ( .C (clk), .D (new_AGEMA_signal_31271), .Q (new_AGEMA_signal_31272) ) ;
    buf_clk new_AGEMA_reg_buffer_10319 ( .C (clk), .D (new_AGEMA_signal_31274), .Q (new_AGEMA_signal_31275) ) ;
    buf_clk new_AGEMA_reg_buffer_10322 ( .C (clk), .D (new_AGEMA_signal_31277), .Q (new_AGEMA_signal_31278) ) ;
    buf_clk new_AGEMA_reg_buffer_10325 ( .C (clk), .D (new_AGEMA_signal_31280), .Q (new_AGEMA_signal_31281) ) ;
    buf_clk new_AGEMA_reg_buffer_10328 ( .C (clk), .D (new_AGEMA_signal_31283), .Q (new_AGEMA_signal_31284) ) ;
    buf_clk new_AGEMA_reg_buffer_10331 ( .C (clk), .D (new_AGEMA_signal_31286), .Q (new_AGEMA_signal_31287) ) ;
    buf_clk new_AGEMA_reg_buffer_10334 ( .C (clk), .D (new_AGEMA_signal_31289), .Q (new_AGEMA_signal_31290) ) ;
    buf_clk new_AGEMA_reg_buffer_10337 ( .C (clk), .D (new_AGEMA_signal_31292), .Q (new_AGEMA_signal_31293) ) ;
    buf_clk new_AGEMA_reg_buffer_10340 ( .C (clk), .D (new_AGEMA_signal_31295), .Q (new_AGEMA_signal_31296) ) ;
    buf_clk new_AGEMA_reg_buffer_10343 ( .C (clk), .D (new_AGEMA_signal_31298), .Q (new_AGEMA_signal_31299) ) ;
    buf_clk new_AGEMA_reg_buffer_10346 ( .C (clk), .D (new_AGEMA_signal_31301), .Q (new_AGEMA_signal_31302) ) ;
    buf_clk new_AGEMA_reg_buffer_10349 ( .C (clk), .D (new_AGEMA_signal_31304), .Q (new_AGEMA_signal_31305) ) ;
    buf_clk new_AGEMA_reg_buffer_10352 ( .C (clk), .D (new_AGEMA_signal_31307), .Q (new_AGEMA_signal_31308) ) ;
    buf_clk new_AGEMA_reg_buffer_10355 ( .C (clk), .D (new_AGEMA_signal_31310), .Q (new_AGEMA_signal_31311) ) ;
    buf_clk new_AGEMA_reg_buffer_10358 ( .C (clk), .D (new_AGEMA_signal_31313), .Q (new_AGEMA_signal_31314) ) ;
    buf_clk new_AGEMA_reg_buffer_10361 ( .C (clk), .D (new_AGEMA_signal_31316), .Q (new_AGEMA_signal_31317) ) ;
    buf_clk new_AGEMA_reg_buffer_10364 ( .C (clk), .D (new_AGEMA_signal_31319), .Q (new_AGEMA_signal_31320) ) ;
    buf_clk new_AGEMA_reg_buffer_10367 ( .C (clk), .D (new_AGEMA_signal_31322), .Q (new_AGEMA_signal_31323) ) ;
    buf_clk new_AGEMA_reg_buffer_10370 ( .C (clk), .D (new_AGEMA_signal_31325), .Q (new_AGEMA_signal_31326) ) ;
    buf_clk new_AGEMA_reg_buffer_10373 ( .C (clk), .D (new_AGEMA_signal_31328), .Q (new_AGEMA_signal_31329) ) ;
    buf_clk new_AGEMA_reg_buffer_10376 ( .C (clk), .D (new_AGEMA_signal_31331), .Q (new_AGEMA_signal_31332) ) ;
    buf_clk new_AGEMA_reg_buffer_10379 ( .C (clk), .D (new_AGEMA_signal_31334), .Q (new_AGEMA_signal_31335) ) ;
    buf_clk new_AGEMA_reg_buffer_10382 ( .C (clk), .D (new_AGEMA_signal_31337), .Q (new_AGEMA_signal_31338) ) ;
    buf_clk new_AGEMA_reg_buffer_10385 ( .C (clk), .D (new_AGEMA_signal_31340), .Q (new_AGEMA_signal_31341) ) ;
    buf_clk new_AGEMA_reg_buffer_10388 ( .C (clk), .D (new_AGEMA_signal_31343), .Q (new_AGEMA_signal_31344) ) ;
    buf_clk new_AGEMA_reg_buffer_10391 ( .C (clk), .D (new_AGEMA_signal_31346), .Q (new_AGEMA_signal_31347) ) ;
    buf_clk new_AGEMA_reg_buffer_10394 ( .C (clk), .D (new_AGEMA_signal_31349), .Q (new_AGEMA_signal_31350) ) ;
    buf_clk new_AGEMA_reg_buffer_10397 ( .C (clk), .D (new_AGEMA_signal_31352), .Q (new_AGEMA_signal_31353) ) ;
    buf_clk new_AGEMA_reg_buffer_10400 ( .C (clk), .D (new_AGEMA_signal_31355), .Q (new_AGEMA_signal_31356) ) ;
    buf_clk new_AGEMA_reg_buffer_10403 ( .C (clk), .D (new_AGEMA_signal_31358), .Q (new_AGEMA_signal_31359) ) ;
    buf_clk new_AGEMA_reg_buffer_10406 ( .C (clk), .D (new_AGEMA_signal_31361), .Q (new_AGEMA_signal_31362) ) ;
    buf_clk new_AGEMA_reg_buffer_10409 ( .C (clk), .D (new_AGEMA_signal_31364), .Q (new_AGEMA_signal_31365) ) ;
    buf_clk new_AGEMA_reg_buffer_10412 ( .C (clk), .D (new_AGEMA_signal_31367), .Q (new_AGEMA_signal_31368) ) ;
    buf_clk new_AGEMA_reg_buffer_10415 ( .C (clk), .D (new_AGEMA_signal_31370), .Q (new_AGEMA_signal_31371) ) ;
    buf_clk new_AGEMA_reg_buffer_10418 ( .C (clk), .D (new_AGEMA_signal_31373), .Q (new_AGEMA_signal_31374) ) ;
    buf_clk new_AGEMA_reg_buffer_10421 ( .C (clk), .D (new_AGEMA_signal_31376), .Q (new_AGEMA_signal_31377) ) ;
    buf_clk new_AGEMA_reg_buffer_10424 ( .C (clk), .D (new_AGEMA_signal_31379), .Q (new_AGEMA_signal_31380) ) ;
    buf_clk new_AGEMA_reg_buffer_10427 ( .C (clk), .D (new_AGEMA_signal_31382), .Q (new_AGEMA_signal_31383) ) ;
    buf_clk new_AGEMA_reg_buffer_10430 ( .C (clk), .D (new_AGEMA_signal_31385), .Q (new_AGEMA_signal_31386) ) ;
    buf_clk new_AGEMA_reg_buffer_10433 ( .C (clk), .D (new_AGEMA_signal_31388), .Q (new_AGEMA_signal_31389) ) ;
    buf_clk new_AGEMA_reg_buffer_10436 ( .C (clk), .D (new_AGEMA_signal_31391), .Q (new_AGEMA_signal_31392) ) ;
    buf_clk new_AGEMA_reg_buffer_10439 ( .C (clk), .D (new_AGEMA_signal_31394), .Q (new_AGEMA_signal_31395) ) ;
    buf_clk new_AGEMA_reg_buffer_10442 ( .C (clk), .D (new_AGEMA_signal_31397), .Q (new_AGEMA_signal_31398) ) ;
    buf_clk new_AGEMA_reg_buffer_10445 ( .C (clk), .D (new_AGEMA_signal_31400), .Q (new_AGEMA_signal_31401) ) ;
    buf_clk new_AGEMA_reg_buffer_10448 ( .C (clk), .D (new_AGEMA_signal_31403), .Q (new_AGEMA_signal_31404) ) ;
    buf_clk new_AGEMA_reg_buffer_10451 ( .C (clk), .D (new_AGEMA_signal_31406), .Q (new_AGEMA_signal_31407) ) ;
    buf_clk new_AGEMA_reg_buffer_10454 ( .C (clk), .D (new_AGEMA_signal_31409), .Q (new_AGEMA_signal_31410) ) ;
    buf_clk new_AGEMA_reg_buffer_10457 ( .C (clk), .D (new_AGEMA_signal_31412), .Q (new_AGEMA_signal_31413) ) ;
    buf_clk new_AGEMA_reg_buffer_10460 ( .C (clk), .D (new_AGEMA_signal_31415), .Q (new_AGEMA_signal_31416) ) ;
    buf_clk new_AGEMA_reg_buffer_10463 ( .C (clk), .D (new_AGEMA_signal_31418), .Q (new_AGEMA_signal_31419) ) ;
    buf_clk new_AGEMA_reg_buffer_10466 ( .C (clk), .D (new_AGEMA_signal_31421), .Q (new_AGEMA_signal_31422) ) ;
    buf_clk new_AGEMA_reg_buffer_10469 ( .C (clk), .D (new_AGEMA_signal_31424), .Q (new_AGEMA_signal_31425) ) ;
    buf_clk new_AGEMA_reg_buffer_10472 ( .C (clk), .D (new_AGEMA_signal_31427), .Q (new_AGEMA_signal_31428) ) ;
    buf_clk new_AGEMA_reg_buffer_10475 ( .C (clk), .D (new_AGEMA_signal_31430), .Q (new_AGEMA_signal_31431) ) ;
    buf_clk new_AGEMA_reg_buffer_10478 ( .C (clk), .D (new_AGEMA_signal_31433), .Q (new_AGEMA_signal_31434) ) ;
    buf_clk new_AGEMA_reg_buffer_10481 ( .C (clk), .D (new_AGEMA_signal_31436), .Q (new_AGEMA_signal_31437) ) ;
    buf_clk new_AGEMA_reg_buffer_10484 ( .C (clk), .D (new_AGEMA_signal_31439), .Q (new_AGEMA_signal_31440) ) ;
    buf_clk new_AGEMA_reg_buffer_10487 ( .C (clk), .D (new_AGEMA_signal_31442), .Q (new_AGEMA_signal_31443) ) ;
    buf_clk new_AGEMA_reg_buffer_10490 ( .C (clk), .D (new_AGEMA_signal_31445), .Q (new_AGEMA_signal_31446) ) ;
    buf_clk new_AGEMA_reg_buffer_10493 ( .C (clk), .D (new_AGEMA_signal_31448), .Q (new_AGEMA_signal_31449) ) ;
    buf_clk new_AGEMA_reg_buffer_10496 ( .C (clk), .D (new_AGEMA_signal_31451), .Q (new_AGEMA_signal_31452) ) ;
    buf_clk new_AGEMA_reg_buffer_10499 ( .C (clk), .D (new_AGEMA_signal_31454), .Q (new_AGEMA_signal_31455) ) ;
    buf_clk new_AGEMA_reg_buffer_10502 ( .C (clk), .D (new_AGEMA_signal_31457), .Q (new_AGEMA_signal_31458) ) ;
    buf_clk new_AGEMA_reg_buffer_10505 ( .C (clk), .D (new_AGEMA_signal_31460), .Q (new_AGEMA_signal_31461) ) ;
    buf_clk new_AGEMA_reg_buffer_10508 ( .C (clk), .D (new_AGEMA_signal_31463), .Q (new_AGEMA_signal_31464) ) ;
    buf_clk new_AGEMA_reg_buffer_10511 ( .C (clk), .D (new_AGEMA_signal_31466), .Q (new_AGEMA_signal_31467) ) ;
    buf_clk new_AGEMA_reg_buffer_10514 ( .C (clk), .D (new_AGEMA_signal_31469), .Q (new_AGEMA_signal_31470) ) ;
    buf_clk new_AGEMA_reg_buffer_10517 ( .C (clk), .D (new_AGEMA_signal_31472), .Q (new_AGEMA_signal_31473) ) ;
    buf_clk new_AGEMA_reg_buffer_10520 ( .C (clk), .D (new_AGEMA_signal_31475), .Q (new_AGEMA_signal_31476) ) ;
    buf_clk new_AGEMA_reg_buffer_10523 ( .C (clk), .D (new_AGEMA_signal_31478), .Q (new_AGEMA_signal_31479) ) ;
    buf_clk new_AGEMA_reg_buffer_10526 ( .C (clk), .D (new_AGEMA_signal_31481), .Q (new_AGEMA_signal_31482) ) ;
    buf_clk new_AGEMA_reg_buffer_10529 ( .C (clk), .D (new_AGEMA_signal_31484), .Q (new_AGEMA_signal_31485) ) ;
    buf_clk new_AGEMA_reg_buffer_10532 ( .C (clk), .D (new_AGEMA_signal_31487), .Q (new_AGEMA_signal_31488) ) ;
    buf_clk new_AGEMA_reg_buffer_10535 ( .C (clk), .D (new_AGEMA_signal_31490), .Q (new_AGEMA_signal_31491) ) ;
    buf_clk new_AGEMA_reg_buffer_10538 ( .C (clk), .D (new_AGEMA_signal_31493), .Q (new_AGEMA_signal_31494) ) ;
    buf_clk new_AGEMA_reg_buffer_10541 ( .C (clk), .D (new_AGEMA_signal_31496), .Q (new_AGEMA_signal_31497) ) ;
    buf_clk new_AGEMA_reg_buffer_10544 ( .C (clk), .D (new_AGEMA_signal_31499), .Q (new_AGEMA_signal_31500) ) ;
    buf_clk new_AGEMA_reg_buffer_10547 ( .C (clk), .D (new_AGEMA_signal_31502), .Q (new_AGEMA_signal_31503) ) ;
    buf_clk new_AGEMA_reg_buffer_10550 ( .C (clk), .D (new_AGEMA_signal_31505), .Q (new_AGEMA_signal_31506) ) ;
    buf_clk new_AGEMA_reg_buffer_10553 ( .C (clk), .D (new_AGEMA_signal_31508), .Q (new_AGEMA_signal_31509) ) ;
    buf_clk new_AGEMA_reg_buffer_10556 ( .C (clk), .D (new_AGEMA_signal_31511), .Q (new_AGEMA_signal_31512) ) ;
    buf_clk new_AGEMA_reg_buffer_10559 ( .C (clk), .D (new_AGEMA_signal_31514), .Q (new_AGEMA_signal_31515) ) ;
    buf_clk new_AGEMA_reg_buffer_10562 ( .C (clk), .D (new_AGEMA_signal_31517), .Q (new_AGEMA_signal_31518) ) ;
    buf_clk new_AGEMA_reg_buffer_10565 ( .C (clk), .D (new_AGEMA_signal_31520), .Q (new_AGEMA_signal_31521) ) ;
    buf_clk new_AGEMA_reg_buffer_10568 ( .C (clk), .D (new_AGEMA_signal_31523), .Q (new_AGEMA_signal_31524) ) ;
    buf_clk new_AGEMA_reg_buffer_10571 ( .C (clk), .D (new_AGEMA_signal_31526), .Q (new_AGEMA_signal_31527) ) ;
    buf_clk new_AGEMA_reg_buffer_10574 ( .C (clk), .D (new_AGEMA_signal_31529), .Q (new_AGEMA_signal_31530) ) ;
    buf_clk new_AGEMA_reg_buffer_10577 ( .C (clk), .D (new_AGEMA_signal_31532), .Q (new_AGEMA_signal_31533) ) ;
    buf_clk new_AGEMA_reg_buffer_10580 ( .C (clk), .D (new_AGEMA_signal_31535), .Q (new_AGEMA_signal_31536) ) ;
    buf_clk new_AGEMA_reg_buffer_10583 ( .C (clk), .D (new_AGEMA_signal_31538), .Q (new_AGEMA_signal_31539) ) ;
    buf_clk new_AGEMA_reg_buffer_10586 ( .C (clk), .D (new_AGEMA_signal_31541), .Q (new_AGEMA_signal_31542) ) ;
    buf_clk new_AGEMA_reg_buffer_10589 ( .C (clk), .D (new_AGEMA_signal_31544), .Q (new_AGEMA_signal_31545) ) ;
    buf_clk new_AGEMA_reg_buffer_10592 ( .C (clk), .D (new_AGEMA_signal_31547), .Q (new_AGEMA_signal_31548) ) ;
    buf_clk new_AGEMA_reg_buffer_10595 ( .C (clk), .D (new_AGEMA_signal_31550), .Q (new_AGEMA_signal_31551) ) ;
    buf_clk new_AGEMA_reg_buffer_10598 ( .C (clk), .D (new_AGEMA_signal_31553), .Q (new_AGEMA_signal_31554) ) ;
    buf_clk new_AGEMA_reg_buffer_10601 ( .C (clk), .D (new_AGEMA_signal_31556), .Q (new_AGEMA_signal_31557) ) ;
    buf_clk new_AGEMA_reg_buffer_10604 ( .C (clk), .D (new_AGEMA_signal_31559), .Q (new_AGEMA_signal_31560) ) ;
    buf_clk new_AGEMA_reg_buffer_10607 ( .C (clk), .D (new_AGEMA_signal_31562), .Q (new_AGEMA_signal_31563) ) ;
    buf_clk new_AGEMA_reg_buffer_10610 ( .C (clk), .D (new_AGEMA_signal_31565), .Q (new_AGEMA_signal_31566) ) ;
    buf_clk new_AGEMA_reg_buffer_10613 ( .C (clk), .D (new_AGEMA_signal_31568), .Q (new_AGEMA_signal_31569) ) ;
    buf_clk new_AGEMA_reg_buffer_10616 ( .C (clk), .D (new_AGEMA_signal_31571), .Q (new_AGEMA_signal_31572) ) ;
    buf_clk new_AGEMA_reg_buffer_10619 ( .C (clk), .D (new_AGEMA_signal_31574), .Q (new_AGEMA_signal_31575) ) ;
    buf_clk new_AGEMA_reg_buffer_10622 ( .C (clk), .D (new_AGEMA_signal_31577), .Q (new_AGEMA_signal_31578) ) ;
    buf_clk new_AGEMA_reg_buffer_10625 ( .C (clk), .D (new_AGEMA_signal_31580), .Q (new_AGEMA_signal_31581) ) ;
    buf_clk new_AGEMA_reg_buffer_10628 ( .C (clk), .D (new_AGEMA_signal_31583), .Q (new_AGEMA_signal_31584) ) ;
    buf_clk new_AGEMA_reg_buffer_10631 ( .C (clk), .D (new_AGEMA_signal_31586), .Q (new_AGEMA_signal_31587) ) ;
    buf_clk new_AGEMA_reg_buffer_10634 ( .C (clk), .D (new_AGEMA_signal_31589), .Q (new_AGEMA_signal_31590) ) ;
    buf_clk new_AGEMA_reg_buffer_10637 ( .C (clk), .D (new_AGEMA_signal_31592), .Q (new_AGEMA_signal_31593) ) ;
    buf_clk new_AGEMA_reg_buffer_10640 ( .C (clk), .D (new_AGEMA_signal_31595), .Q (new_AGEMA_signal_31596) ) ;
    buf_clk new_AGEMA_reg_buffer_10643 ( .C (clk), .D (new_AGEMA_signal_31598), .Q (new_AGEMA_signal_31599) ) ;
    buf_clk new_AGEMA_reg_buffer_10646 ( .C (clk), .D (new_AGEMA_signal_31601), .Q (new_AGEMA_signal_31602) ) ;
    buf_clk new_AGEMA_reg_buffer_10649 ( .C (clk), .D (new_AGEMA_signal_31604), .Q (new_AGEMA_signal_31605) ) ;
    buf_clk new_AGEMA_reg_buffer_10652 ( .C (clk), .D (new_AGEMA_signal_31607), .Q (new_AGEMA_signal_31608) ) ;
    buf_clk new_AGEMA_reg_buffer_10655 ( .C (clk), .D (new_AGEMA_signal_31610), .Q (new_AGEMA_signal_31611) ) ;
    buf_clk new_AGEMA_reg_buffer_10658 ( .C (clk), .D (new_AGEMA_signal_31613), .Q (new_AGEMA_signal_31614) ) ;
    buf_clk new_AGEMA_reg_buffer_10661 ( .C (clk), .D (new_AGEMA_signal_31616), .Q (new_AGEMA_signal_31617) ) ;
    buf_clk new_AGEMA_reg_buffer_10664 ( .C (clk), .D (new_AGEMA_signal_31619), .Q (new_AGEMA_signal_31620) ) ;
    buf_clk new_AGEMA_reg_buffer_10667 ( .C (clk), .D (new_AGEMA_signal_31622), .Q (new_AGEMA_signal_31623) ) ;
    buf_clk new_AGEMA_reg_buffer_10670 ( .C (clk), .D (new_AGEMA_signal_31625), .Q (new_AGEMA_signal_31626) ) ;
    buf_clk new_AGEMA_reg_buffer_10673 ( .C (clk), .D (new_AGEMA_signal_31628), .Q (new_AGEMA_signal_31629) ) ;
    buf_clk new_AGEMA_reg_buffer_10676 ( .C (clk), .D (new_AGEMA_signal_31631), .Q (new_AGEMA_signal_31632) ) ;
    buf_clk new_AGEMA_reg_buffer_10679 ( .C (clk), .D (new_AGEMA_signal_31634), .Q (new_AGEMA_signal_31635) ) ;
    buf_clk new_AGEMA_reg_buffer_10682 ( .C (clk), .D (new_AGEMA_signal_31637), .Q (new_AGEMA_signal_31638) ) ;
    buf_clk new_AGEMA_reg_buffer_10685 ( .C (clk), .D (new_AGEMA_signal_31640), .Q (new_AGEMA_signal_31641) ) ;
    buf_clk new_AGEMA_reg_buffer_10688 ( .C (clk), .D (new_AGEMA_signal_31643), .Q (new_AGEMA_signal_31644) ) ;
    buf_clk new_AGEMA_reg_buffer_10691 ( .C (clk), .D (new_AGEMA_signal_31646), .Q (new_AGEMA_signal_31647) ) ;
    buf_clk new_AGEMA_reg_buffer_10694 ( .C (clk), .D (new_AGEMA_signal_31649), .Q (new_AGEMA_signal_31650) ) ;
    buf_clk new_AGEMA_reg_buffer_10697 ( .C (clk), .D (new_AGEMA_signal_31652), .Q (new_AGEMA_signal_31653) ) ;
    buf_clk new_AGEMA_reg_buffer_10700 ( .C (clk), .D (new_AGEMA_signal_31655), .Q (new_AGEMA_signal_31656) ) ;
    buf_clk new_AGEMA_reg_buffer_10703 ( .C (clk), .D (new_AGEMA_signal_31658), .Q (new_AGEMA_signal_31659) ) ;
    buf_clk new_AGEMA_reg_buffer_10706 ( .C (clk), .D (new_AGEMA_signal_31661), .Q (new_AGEMA_signal_31662) ) ;
    buf_clk new_AGEMA_reg_buffer_10710 ( .C (clk), .D (new_AGEMA_signal_31665), .Q (new_AGEMA_signal_31666) ) ;
    buf_clk new_AGEMA_reg_buffer_10714 ( .C (clk), .D (new_AGEMA_signal_31669), .Q (new_AGEMA_signal_31670) ) ;
    buf_clk new_AGEMA_reg_buffer_10718 ( .C (clk), .D (new_AGEMA_signal_31673), .Q (new_AGEMA_signal_31674) ) ;
    buf_clk new_AGEMA_reg_buffer_10722 ( .C (clk), .D (new_AGEMA_signal_31677), .Q (new_AGEMA_signal_31678) ) ;
    buf_clk new_AGEMA_reg_buffer_10726 ( .C (clk), .D (new_AGEMA_signal_31681), .Q (new_AGEMA_signal_31682) ) ;
    buf_clk new_AGEMA_reg_buffer_10730 ( .C (clk), .D (new_AGEMA_signal_31685), .Q (new_AGEMA_signal_31686) ) ;
    buf_clk new_AGEMA_reg_buffer_10734 ( .C (clk), .D (new_AGEMA_signal_31689), .Q (new_AGEMA_signal_31690) ) ;
    buf_clk new_AGEMA_reg_buffer_10738 ( .C (clk), .D (new_AGEMA_signal_31693), .Q (new_AGEMA_signal_31694) ) ;
    buf_clk new_AGEMA_reg_buffer_10742 ( .C (clk), .D (new_AGEMA_signal_31697), .Q (new_AGEMA_signal_31698) ) ;
    buf_clk new_AGEMA_reg_buffer_10746 ( .C (clk), .D (new_AGEMA_signal_31701), .Q (new_AGEMA_signal_31702) ) ;
    buf_clk new_AGEMA_reg_buffer_10750 ( .C (clk), .D (new_AGEMA_signal_31705), .Q (new_AGEMA_signal_31706) ) ;
    buf_clk new_AGEMA_reg_buffer_10754 ( .C (clk), .D (new_AGEMA_signal_31709), .Q (new_AGEMA_signal_31710) ) ;
    buf_clk new_AGEMA_reg_buffer_10758 ( .C (clk), .D (new_AGEMA_signal_31713), .Q (new_AGEMA_signal_31714) ) ;
    buf_clk new_AGEMA_reg_buffer_10762 ( .C (clk), .D (new_AGEMA_signal_31717), .Q (new_AGEMA_signal_31718) ) ;
    buf_clk new_AGEMA_reg_buffer_10766 ( .C (clk), .D (new_AGEMA_signal_31721), .Q (new_AGEMA_signal_31722) ) ;
    buf_clk new_AGEMA_reg_buffer_10770 ( .C (clk), .D (new_AGEMA_signal_31725), .Q (new_AGEMA_signal_31726) ) ;
    buf_clk new_AGEMA_reg_buffer_10774 ( .C (clk), .D (new_AGEMA_signal_31729), .Q (new_AGEMA_signal_31730) ) ;
    buf_clk new_AGEMA_reg_buffer_10778 ( .C (clk), .D (new_AGEMA_signal_31733), .Q (new_AGEMA_signal_31734) ) ;
    buf_clk new_AGEMA_reg_buffer_10782 ( .C (clk), .D (new_AGEMA_signal_31737), .Q (new_AGEMA_signal_31738) ) ;
    buf_clk new_AGEMA_reg_buffer_10786 ( .C (clk), .D (new_AGEMA_signal_31741), .Q (new_AGEMA_signal_31742) ) ;
    buf_clk new_AGEMA_reg_buffer_10790 ( .C (clk), .D (new_AGEMA_signal_31745), .Q (new_AGEMA_signal_31746) ) ;
    buf_clk new_AGEMA_reg_buffer_10794 ( .C (clk), .D (new_AGEMA_signal_31749), .Q (new_AGEMA_signal_31750) ) ;
    buf_clk new_AGEMA_reg_buffer_10798 ( .C (clk), .D (new_AGEMA_signal_31753), .Q (new_AGEMA_signal_31754) ) ;
    buf_clk new_AGEMA_reg_buffer_10802 ( .C (clk), .D (new_AGEMA_signal_31757), .Q (new_AGEMA_signal_31758) ) ;
    buf_clk new_AGEMA_reg_buffer_10806 ( .C (clk), .D (new_AGEMA_signal_31761), .Q (new_AGEMA_signal_31762) ) ;
    buf_clk new_AGEMA_reg_buffer_10810 ( .C (clk), .D (new_AGEMA_signal_31765), .Q (new_AGEMA_signal_31766) ) ;
    buf_clk new_AGEMA_reg_buffer_10814 ( .C (clk), .D (new_AGEMA_signal_31769), .Q (new_AGEMA_signal_31770) ) ;
    buf_clk new_AGEMA_reg_buffer_10818 ( .C (clk), .D (new_AGEMA_signal_31773), .Q (new_AGEMA_signal_31774) ) ;
    buf_clk new_AGEMA_reg_buffer_10822 ( .C (clk), .D (new_AGEMA_signal_31777), .Q (new_AGEMA_signal_31778) ) ;
    buf_clk new_AGEMA_reg_buffer_10826 ( .C (clk), .D (new_AGEMA_signal_31781), .Q (new_AGEMA_signal_31782) ) ;
    buf_clk new_AGEMA_reg_buffer_10830 ( .C (clk), .D (new_AGEMA_signal_31785), .Q (new_AGEMA_signal_31786) ) ;
    buf_clk new_AGEMA_reg_buffer_10834 ( .C (clk), .D (new_AGEMA_signal_31789), .Q (new_AGEMA_signal_31790) ) ;
    buf_clk new_AGEMA_reg_buffer_10838 ( .C (clk), .D (new_AGEMA_signal_31793), .Q (new_AGEMA_signal_31794) ) ;
    buf_clk new_AGEMA_reg_buffer_10842 ( .C (clk), .D (new_AGEMA_signal_31797), .Q (new_AGEMA_signal_31798) ) ;
    buf_clk new_AGEMA_reg_buffer_10846 ( .C (clk), .D (new_AGEMA_signal_31801), .Q (new_AGEMA_signal_31802) ) ;
    buf_clk new_AGEMA_reg_buffer_10850 ( .C (clk), .D (new_AGEMA_signal_31805), .Q (new_AGEMA_signal_31806) ) ;
    buf_clk new_AGEMA_reg_buffer_10854 ( .C (clk), .D (new_AGEMA_signal_31809), .Q (new_AGEMA_signal_31810) ) ;
    buf_clk new_AGEMA_reg_buffer_10858 ( .C (clk), .D (new_AGEMA_signal_31813), .Q (new_AGEMA_signal_31814) ) ;
    buf_clk new_AGEMA_reg_buffer_10862 ( .C (clk), .D (new_AGEMA_signal_31817), .Q (new_AGEMA_signal_31818) ) ;
    buf_clk new_AGEMA_reg_buffer_10866 ( .C (clk), .D (new_AGEMA_signal_31821), .Q (new_AGEMA_signal_31822) ) ;
    buf_clk new_AGEMA_reg_buffer_10870 ( .C (clk), .D (new_AGEMA_signal_31825), .Q (new_AGEMA_signal_31826) ) ;
    buf_clk new_AGEMA_reg_buffer_10874 ( .C (clk), .D (new_AGEMA_signal_31829), .Q (new_AGEMA_signal_31830) ) ;
    buf_clk new_AGEMA_reg_buffer_10878 ( .C (clk), .D (new_AGEMA_signal_31833), .Q (new_AGEMA_signal_31834) ) ;
    buf_clk new_AGEMA_reg_buffer_10882 ( .C (clk), .D (new_AGEMA_signal_31837), .Q (new_AGEMA_signal_31838) ) ;
    buf_clk new_AGEMA_reg_buffer_10886 ( .C (clk), .D (new_AGEMA_signal_31841), .Q (new_AGEMA_signal_31842) ) ;
    buf_clk new_AGEMA_reg_buffer_10890 ( .C (clk), .D (new_AGEMA_signal_31845), .Q (new_AGEMA_signal_31846) ) ;
    buf_clk new_AGEMA_reg_buffer_10894 ( .C (clk), .D (new_AGEMA_signal_31849), .Q (new_AGEMA_signal_31850) ) ;
    buf_clk new_AGEMA_reg_buffer_10898 ( .C (clk), .D (new_AGEMA_signal_31853), .Q (new_AGEMA_signal_31854) ) ;
    buf_clk new_AGEMA_reg_buffer_10902 ( .C (clk), .D (new_AGEMA_signal_31857), .Q (new_AGEMA_signal_31858) ) ;
    buf_clk new_AGEMA_reg_buffer_10906 ( .C (clk), .D (new_AGEMA_signal_31861), .Q (new_AGEMA_signal_31862) ) ;
    buf_clk new_AGEMA_reg_buffer_10910 ( .C (clk), .D (new_AGEMA_signal_31865), .Q (new_AGEMA_signal_31866) ) ;
    buf_clk new_AGEMA_reg_buffer_10914 ( .C (clk), .D (new_AGEMA_signal_31869), .Q (new_AGEMA_signal_31870) ) ;
    buf_clk new_AGEMA_reg_buffer_10918 ( .C (clk), .D (new_AGEMA_signal_31873), .Q (new_AGEMA_signal_31874) ) ;
    buf_clk new_AGEMA_reg_buffer_10922 ( .C (clk), .D (new_AGEMA_signal_31877), .Q (new_AGEMA_signal_31878) ) ;
    buf_clk new_AGEMA_reg_buffer_10926 ( .C (clk), .D (new_AGEMA_signal_31881), .Q (new_AGEMA_signal_31882) ) ;
    buf_clk new_AGEMA_reg_buffer_10930 ( .C (clk), .D (new_AGEMA_signal_31885), .Q (new_AGEMA_signal_31886) ) ;
    buf_clk new_AGEMA_reg_buffer_10934 ( .C (clk), .D (new_AGEMA_signal_31889), .Q (new_AGEMA_signal_31890) ) ;
    buf_clk new_AGEMA_reg_buffer_10938 ( .C (clk), .D (new_AGEMA_signal_31893), .Q (new_AGEMA_signal_31894) ) ;
    buf_clk new_AGEMA_reg_buffer_10942 ( .C (clk), .D (new_AGEMA_signal_31897), .Q (new_AGEMA_signal_31898) ) ;
    buf_clk new_AGEMA_reg_buffer_10946 ( .C (clk), .D (new_AGEMA_signal_31901), .Q (new_AGEMA_signal_31902) ) ;
    buf_clk new_AGEMA_reg_buffer_10950 ( .C (clk), .D (new_AGEMA_signal_31905), .Q (new_AGEMA_signal_31906) ) ;
    buf_clk new_AGEMA_reg_buffer_10954 ( .C (clk), .D (new_AGEMA_signal_31909), .Q (new_AGEMA_signal_31910) ) ;
    buf_clk new_AGEMA_reg_buffer_10958 ( .C (clk), .D (new_AGEMA_signal_31913), .Q (new_AGEMA_signal_31914) ) ;
    buf_clk new_AGEMA_reg_buffer_10962 ( .C (clk), .D (new_AGEMA_signal_31917), .Q (new_AGEMA_signal_31918) ) ;
    buf_clk new_AGEMA_reg_buffer_10966 ( .C (clk), .D (new_AGEMA_signal_31921), .Q (new_AGEMA_signal_31922) ) ;
    buf_clk new_AGEMA_reg_buffer_10970 ( .C (clk), .D (new_AGEMA_signal_31925), .Q (new_AGEMA_signal_31926) ) ;
    buf_clk new_AGEMA_reg_buffer_10974 ( .C (clk), .D (new_AGEMA_signal_31929), .Q (new_AGEMA_signal_31930) ) ;
    buf_clk new_AGEMA_reg_buffer_10978 ( .C (clk), .D (new_AGEMA_signal_31933), .Q (new_AGEMA_signal_31934) ) ;
    buf_clk new_AGEMA_reg_buffer_10982 ( .C (clk), .D (new_AGEMA_signal_31937), .Q (new_AGEMA_signal_31938) ) ;
    buf_clk new_AGEMA_reg_buffer_10986 ( .C (clk), .D (new_AGEMA_signal_31941), .Q (new_AGEMA_signal_31942) ) ;
    buf_clk new_AGEMA_reg_buffer_10990 ( .C (clk), .D (new_AGEMA_signal_31945), .Q (new_AGEMA_signal_31946) ) ;
    buf_clk new_AGEMA_reg_buffer_10994 ( .C (clk), .D (new_AGEMA_signal_31949), .Q (new_AGEMA_signal_31950) ) ;
    buf_clk new_AGEMA_reg_buffer_10998 ( .C (clk), .D (new_AGEMA_signal_31953), .Q (new_AGEMA_signal_31954) ) ;
    buf_clk new_AGEMA_reg_buffer_11002 ( .C (clk), .D (new_AGEMA_signal_31957), .Q (new_AGEMA_signal_31958) ) ;
    buf_clk new_AGEMA_reg_buffer_11006 ( .C (clk), .D (new_AGEMA_signal_31961), .Q (new_AGEMA_signal_31962) ) ;
    buf_clk new_AGEMA_reg_buffer_11010 ( .C (clk), .D (new_AGEMA_signal_31965), .Q (new_AGEMA_signal_31966) ) ;
    buf_clk new_AGEMA_reg_buffer_11014 ( .C (clk), .D (new_AGEMA_signal_31969), .Q (new_AGEMA_signal_31970) ) ;
    buf_clk new_AGEMA_reg_buffer_11018 ( .C (clk), .D (new_AGEMA_signal_31973), .Q (new_AGEMA_signal_31974) ) ;
    buf_clk new_AGEMA_reg_buffer_11022 ( .C (clk), .D (new_AGEMA_signal_31977), .Q (new_AGEMA_signal_31978) ) ;
    buf_clk new_AGEMA_reg_buffer_11026 ( .C (clk), .D (new_AGEMA_signal_31981), .Q (new_AGEMA_signal_31982) ) ;
    buf_clk new_AGEMA_reg_buffer_11030 ( .C (clk), .D (new_AGEMA_signal_31985), .Q (new_AGEMA_signal_31986) ) ;
    buf_clk new_AGEMA_reg_buffer_11034 ( .C (clk), .D (new_AGEMA_signal_31989), .Q (new_AGEMA_signal_31990) ) ;
    buf_clk new_AGEMA_reg_buffer_11038 ( .C (clk), .D (new_AGEMA_signal_31993), .Q (new_AGEMA_signal_31994) ) ;
    buf_clk new_AGEMA_reg_buffer_11042 ( .C (clk), .D (new_AGEMA_signal_31997), .Q (new_AGEMA_signal_31998) ) ;
    buf_clk new_AGEMA_reg_buffer_11046 ( .C (clk), .D (new_AGEMA_signal_32001), .Q (new_AGEMA_signal_32002) ) ;
    buf_clk new_AGEMA_reg_buffer_11050 ( .C (clk), .D (new_AGEMA_signal_32005), .Q (new_AGEMA_signal_32006) ) ;
    buf_clk new_AGEMA_reg_buffer_11054 ( .C (clk), .D (new_AGEMA_signal_32009), .Q (new_AGEMA_signal_32010) ) ;
    buf_clk new_AGEMA_reg_buffer_11058 ( .C (clk), .D (new_AGEMA_signal_32013), .Q (new_AGEMA_signal_32014) ) ;
    buf_clk new_AGEMA_reg_buffer_11062 ( .C (clk), .D (new_AGEMA_signal_32017), .Q (new_AGEMA_signal_32018) ) ;
    buf_clk new_AGEMA_reg_buffer_11066 ( .C (clk), .D (new_AGEMA_signal_32021), .Q (new_AGEMA_signal_32022) ) ;
    buf_clk new_AGEMA_reg_buffer_11070 ( .C (clk), .D (new_AGEMA_signal_32025), .Q (new_AGEMA_signal_32026) ) ;
    buf_clk new_AGEMA_reg_buffer_11074 ( .C (clk), .D (new_AGEMA_signal_32029), .Q (new_AGEMA_signal_32030) ) ;
    buf_clk new_AGEMA_reg_buffer_11078 ( .C (clk), .D (new_AGEMA_signal_32033), .Q (new_AGEMA_signal_32034) ) ;
    buf_clk new_AGEMA_reg_buffer_11082 ( .C (clk), .D (new_AGEMA_signal_32037), .Q (new_AGEMA_signal_32038) ) ;
    buf_clk new_AGEMA_reg_buffer_11086 ( .C (clk), .D (new_AGEMA_signal_32041), .Q (new_AGEMA_signal_32042) ) ;
    buf_clk new_AGEMA_reg_buffer_11090 ( .C (clk), .D (new_AGEMA_signal_32045), .Q (new_AGEMA_signal_32046) ) ;
    buf_clk new_AGEMA_reg_buffer_11094 ( .C (clk), .D (new_AGEMA_signal_32049), .Q (new_AGEMA_signal_32050) ) ;
    buf_clk new_AGEMA_reg_buffer_11098 ( .C (clk), .D (new_AGEMA_signal_32053), .Q (new_AGEMA_signal_32054) ) ;
    buf_clk new_AGEMA_reg_buffer_11102 ( .C (clk), .D (new_AGEMA_signal_32057), .Q (new_AGEMA_signal_32058) ) ;
    buf_clk new_AGEMA_reg_buffer_11106 ( .C (clk), .D (new_AGEMA_signal_32061), .Q (new_AGEMA_signal_32062) ) ;
    buf_clk new_AGEMA_reg_buffer_11110 ( .C (clk), .D (new_AGEMA_signal_32065), .Q (new_AGEMA_signal_32066) ) ;
    buf_clk new_AGEMA_reg_buffer_11114 ( .C (clk), .D (new_AGEMA_signal_32069), .Q (new_AGEMA_signal_32070) ) ;
    buf_clk new_AGEMA_reg_buffer_11118 ( .C (clk), .D (new_AGEMA_signal_32073), .Q (new_AGEMA_signal_32074) ) ;
    buf_clk new_AGEMA_reg_buffer_11122 ( .C (clk), .D (new_AGEMA_signal_32077), .Q (new_AGEMA_signal_32078) ) ;
    buf_clk new_AGEMA_reg_buffer_11126 ( .C (clk), .D (new_AGEMA_signal_32081), .Q (new_AGEMA_signal_32082) ) ;
    buf_clk new_AGEMA_reg_buffer_11130 ( .C (clk), .D (new_AGEMA_signal_32085), .Q (new_AGEMA_signal_32086) ) ;
    buf_clk new_AGEMA_reg_buffer_11134 ( .C (clk), .D (new_AGEMA_signal_32089), .Q (new_AGEMA_signal_32090) ) ;
    buf_clk new_AGEMA_reg_buffer_11138 ( .C (clk), .D (new_AGEMA_signal_32093), .Q (new_AGEMA_signal_32094) ) ;
    buf_clk new_AGEMA_reg_buffer_11142 ( .C (clk), .D (new_AGEMA_signal_32097), .Q (new_AGEMA_signal_32098) ) ;
    buf_clk new_AGEMA_reg_buffer_11146 ( .C (clk), .D (new_AGEMA_signal_32101), .Q (new_AGEMA_signal_32102) ) ;
    buf_clk new_AGEMA_reg_buffer_11150 ( .C (clk), .D (new_AGEMA_signal_32105), .Q (new_AGEMA_signal_32106) ) ;
    buf_clk new_AGEMA_reg_buffer_11154 ( .C (clk), .D (new_AGEMA_signal_32109), .Q (new_AGEMA_signal_32110) ) ;
    buf_clk new_AGEMA_reg_buffer_11158 ( .C (clk), .D (new_AGEMA_signal_32113), .Q (new_AGEMA_signal_32114) ) ;
    buf_clk new_AGEMA_reg_buffer_11162 ( .C (clk), .D (new_AGEMA_signal_32117), .Q (new_AGEMA_signal_32118) ) ;
    buf_clk new_AGEMA_reg_buffer_11166 ( .C (clk), .D (new_AGEMA_signal_32121), .Q (new_AGEMA_signal_32122) ) ;
    buf_clk new_AGEMA_reg_buffer_11170 ( .C (clk), .D (new_AGEMA_signal_32125), .Q (new_AGEMA_signal_32126) ) ;
    buf_clk new_AGEMA_reg_buffer_11174 ( .C (clk), .D (new_AGEMA_signal_32129), .Q (new_AGEMA_signal_32130) ) ;
    buf_clk new_AGEMA_reg_buffer_11178 ( .C (clk), .D (new_AGEMA_signal_32133), .Q (new_AGEMA_signal_32134) ) ;
    buf_clk new_AGEMA_reg_buffer_11182 ( .C (clk), .D (new_AGEMA_signal_32137), .Q (new_AGEMA_signal_32138) ) ;
    buf_clk new_AGEMA_reg_buffer_11186 ( .C (clk), .D (new_AGEMA_signal_32141), .Q (new_AGEMA_signal_32142) ) ;
    buf_clk new_AGEMA_reg_buffer_11190 ( .C (clk), .D (new_AGEMA_signal_32145), .Q (new_AGEMA_signal_32146) ) ;
    buf_clk new_AGEMA_reg_buffer_11194 ( .C (clk), .D (new_AGEMA_signal_32149), .Q (new_AGEMA_signal_32150) ) ;
    buf_clk new_AGEMA_reg_buffer_11198 ( .C (clk), .D (new_AGEMA_signal_32153), .Q (new_AGEMA_signal_32154) ) ;
    buf_clk new_AGEMA_reg_buffer_11202 ( .C (clk), .D (new_AGEMA_signal_32157), .Q (new_AGEMA_signal_32158) ) ;
    buf_clk new_AGEMA_reg_buffer_11206 ( .C (clk), .D (new_AGEMA_signal_32161), .Q (new_AGEMA_signal_32162) ) ;
    buf_clk new_AGEMA_reg_buffer_11210 ( .C (clk), .D (new_AGEMA_signal_32165), .Q (new_AGEMA_signal_32166) ) ;
    buf_clk new_AGEMA_reg_buffer_11214 ( .C (clk), .D (new_AGEMA_signal_32169), .Q (new_AGEMA_signal_32170) ) ;
    buf_clk new_AGEMA_reg_buffer_11218 ( .C (clk), .D (new_AGEMA_signal_32173), .Q (new_AGEMA_signal_32174) ) ;
    buf_clk new_AGEMA_reg_buffer_11222 ( .C (clk), .D (new_AGEMA_signal_32177), .Q (new_AGEMA_signal_32178) ) ;
    buf_clk new_AGEMA_reg_buffer_11226 ( .C (clk), .D (new_AGEMA_signal_32181), .Q (new_AGEMA_signal_32182) ) ;
    buf_clk new_AGEMA_reg_buffer_11230 ( .C (clk), .D (new_AGEMA_signal_32185), .Q (new_AGEMA_signal_32186) ) ;
    buf_clk new_AGEMA_reg_buffer_11234 ( .C (clk), .D (new_AGEMA_signal_32189), .Q (new_AGEMA_signal_32190) ) ;
    buf_clk new_AGEMA_reg_buffer_11238 ( .C (clk), .D (new_AGEMA_signal_32193), .Q (new_AGEMA_signal_32194) ) ;
    buf_clk new_AGEMA_reg_buffer_11242 ( .C (clk), .D (new_AGEMA_signal_32197), .Q (new_AGEMA_signal_32198) ) ;
    buf_clk new_AGEMA_reg_buffer_11246 ( .C (clk), .D (new_AGEMA_signal_32201), .Q (new_AGEMA_signal_32202) ) ;
    buf_clk new_AGEMA_reg_buffer_11250 ( .C (clk), .D (new_AGEMA_signal_32205), .Q (new_AGEMA_signal_32206) ) ;
    buf_clk new_AGEMA_reg_buffer_11254 ( .C (clk), .D (new_AGEMA_signal_32209), .Q (new_AGEMA_signal_32210) ) ;
    buf_clk new_AGEMA_reg_buffer_11258 ( .C (clk), .D (new_AGEMA_signal_32213), .Q (new_AGEMA_signal_32214) ) ;
    buf_clk new_AGEMA_reg_buffer_11262 ( .C (clk), .D (new_AGEMA_signal_32217), .Q (new_AGEMA_signal_32218) ) ;
    buf_clk new_AGEMA_reg_buffer_11266 ( .C (clk), .D (new_AGEMA_signal_32221), .Q (new_AGEMA_signal_32222) ) ;
    buf_clk new_AGEMA_reg_buffer_11270 ( .C (clk), .D (new_AGEMA_signal_32225), .Q (new_AGEMA_signal_32226) ) ;
    buf_clk new_AGEMA_reg_buffer_11274 ( .C (clk), .D (new_AGEMA_signal_32229), .Q (new_AGEMA_signal_32230) ) ;
    buf_clk new_AGEMA_reg_buffer_11278 ( .C (clk), .D (new_AGEMA_signal_32233), .Q (new_AGEMA_signal_32234) ) ;
    buf_clk new_AGEMA_reg_buffer_11282 ( .C (clk), .D (new_AGEMA_signal_32237), .Q (new_AGEMA_signal_32238) ) ;
    buf_clk new_AGEMA_reg_buffer_11286 ( .C (clk), .D (new_AGEMA_signal_32241), .Q (new_AGEMA_signal_32242) ) ;
    buf_clk new_AGEMA_reg_buffer_11290 ( .C (clk), .D (new_AGEMA_signal_32245), .Q (new_AGEMA_signal_32246) ) ;
    buf_clk new_AGEMA_reg_buffer_11294 ( .C (clk), .D (new_AGEMA_signal_32249), .Q (new_AGEMA_signal_32250) ) ;
    buf_clk new_AGEMA_reg_buffer_11298 ( .C (clk), .D (new_AGEMA_signal_32253), .Q (new_AGEMA_signal_32254) ) ;
    buf_clk new_AGEMA_reg_buffer_11302 ( .C (clk), .D (new_AGEMA_signal_32257), .Q (new_AGEMA_signal_32258) ) ;
    buf_clk new_AGEMA_reg_buffer_11306 ( .C (clk), .D (new_AGEMA_signal_32261), .Q (new_AGEMA_signal_32262) ) ;
    buf_clk new_AGEMA_reg_buffer_11310 ( .C (clk), .D (new_AGEMA_signal_32265), .Q (new_AGEMA_signal_32266) ) ;
    buf_clk new_AGEMA_reg_buffer_11314 ( .C (clk), .D (new_AGEMA_signal_32269), .Q (new_AGEMA_signal_32270) ) ;
    buf_clk new_AGEMA_reg_buffer_11318 ( .C (clk), .D (new_AGEMA_signal_32273), .Q (new_AGEMA_signal_32274) ) ;
    buf_clk new_AGEMA_reg_buffer_11322 ( .C (clk), .D (new_AGEMA_signal_32277), .Q (new_AGEMA_signal_32278) ) ;
    buf_clk new_AGEMA_reg_buffer_11326 ( .C (clk), .D (new_AGEMA_signal_32281), .Q (new_AGEMA_signal_32282) ) ;
    buf_clk new_AGEMA_reg_buffer_11330 ( .C (clk), .D (new_AGEMA_signal_32285), .Q (new_AGEMA_signal_32286) ) ;
    buf_clk new_AGEMA_reg_buffer_11334 ( .C (clk), .D (new_AGEMA_signal_32289), .Q (new_AGEMA_signal_32290) ) ;
    buf_clk new_AGEMA_reg_buffer_11338 ( .C (clk), .D (new_AGEMA_signal_32293), .Q (new_AGEMA_signal_32294) ) ;
    buf_clk new_AGEMA_reg_buffer_11342 ( .C (clk), .D (new_AGEMA_signal_32297), .Q (new_AGEMA_signal_32298) ) ;
    buf_clk new_AGEMA_reg_buffer_11346 ( .C (clk), .D (new_AGEMA_signal_32301), .Q (new_AGEMA_signal_32302) ) ;
    buf_clk new_AGEMA_reg_buffer_11350 ( .C (clk), .D (new_AGEMA_signal_32305), .Q (new_AGEMA_signal_32306) ) ;
    buf_clk new_AGEMA_reg_buffer_11354 ( .C (clk), .D (new_AGEMA_signal_32309), .Q (new_AGEMA_signal_32310) ) ;
    buf_clk new_AGEMA_reg_buffer_11358 ( .C (clk), .D (new_AGEMA_signal_32313), .Q (new_AGEMA_signal_32314) ) ;
    buf_clk new_AGEMA_reg_buffer_11362 ( .C (clk), .D (new_AGEMA_signal_32317), .Q (new_AGEMA_signal_32318) ) ;
    buf_clk new_AGEMA_reg_buffer_11366 ( .C (clk), .D (new_AGEMA_signal_32321), .Q (new_AGEMA_signal_32322) ) ;
    buf_clk new_AGEMA_reg_buffer_11370 ( .C (clk), .D (new_AGEMA_signal_32325), .Q (new_AGEMA_signal_32326) ) ;
    buf_clk new_AGEMA_reg_buffer_11374 ( .C (clk), .D (new_AGEMA_signal_32329), .Q (new_AGEMA_signal_32330) ) ;
    buf_clk new_AGEMA_reg_buffer_11378 ( .C (clk), .D (new_AGEMA_signal_32333), .Q (new_AGEMA_signal_32334) ) ;
    buf_clk new_AGEMA_reg_buffer_11382 ( .C (clk), .D (new_AGEMA_signal_32337), .Q (new_AGEMA_signal_32338) ) ;
    buf_clk new_AGEMA_reg_buffer_11386 ( .C (clk), .D (new_AGEMA_signal_32341), .Q (new_AGEMA_signal_32342) ) ;
    buf_clk new_AGEMA_reg_buffer_11390 ( .C (clk), .D (new_AGEMA_signal_32345), .Q (new_AGEMA_signal_32346) ) ;
    buf_clk new_AGEMA_reg_buffer_11394 ( .C (clk), .D (new_AGEMA_signal_32349), .Q (new_AGEMA_signal_32350) ) ;
    buf_clk new_AGEMA_reg_buffer_11398 ( .C (clk), .D (new_AGEMA_signal_32353), .Q (new_AGEMA_signal_32354) ) ;
    buf_clk new_AGEMA_reg_buffer_11402 ( .C (clk), .D (new_AGEMA_signal_32357), .Q (new_AGEMA_signal_32358) ) ;
    buf_clk new_AGEMA_reg_buffer_11406 ( .C (clk), .D (new_AGEMA_signal_32361), .Q (new_AGEMA_signal_32362) ) ;
    buf_clk new_AGEMA_reg_buffer_11410 ( .C (clk), .D (new_AGEMA_signal_32365), .Q (new_AGEMA_signal_32366) ) ;
    buf_clk new_AGEMA_reg_buffer_11414 ( .C (clk), .D (new_AGEMA_signal_32369), .Q (new_AGEMA_signal_32370) ) ;
    buf_clk new_AGEMA_reg_buffer_11418 ( .C (clk), .D (new_AGEMA_signal_32373), .Q (new_AGEMA_signal_32374) ) ;
    buf_clk new_AGEMA_reg_buffer_11422 ( .C (clk), .D (new_AGEMA_signal_32377), .Q (new_AGEMA_signal_32378) ) ;
    buf_clk new_AGEMA_reg_buffer_11426 ( .C (clk), .D (new_AGEMA_signal_32381), .Q (new_AGEMA_signal_32382) ) ;
    buf_clk new_AGEMA_reg_buffer_11430 ( .C (clk), .D (new_AGEMA_signal_32385), .Q (new_AGEMA_signal_32386) ) ;
    buf_clk new_AGEMA_reg_buffer_11434 ( .C (clk), .D (new_AGEMA_signal_32389), .Q (new_AGEMA_signal_32390) ) ;
    buf_clk new_AGEMA_reg_buffer_11438 ( .C (clk), .D (new_AGEMA_signal_32393), .Q (new_AGEMA_signal_32394) ) ;
    buf_clk new_AGEMA_reg_buffer_11442 ( .C (clk), .D (new_AGEMA_signal_32397), .Q (new_AGEMA_signal_32398) ) ;
    buf_clk new_AGEMA_reg_buffer_11446 ( .C (clk), .D (new_AGEMA_signal_32401), .Q (new_AGEMA_signal_32402) ) ;
    buf_clk new_AGEMA_reg_buffer_11450 ( .C (clk), .D (new_AGEMA_signal_32405), .Q (new_AGEMA_signal_32406) ) ;
    buf_clk new_AGEMA_reg_buffer_11454 ( .C (clk), .D (new_AGEMA_signal_32409), .Q (new_AGEMA_signal_32410) ) ;
    buf_clk new_AGEMA_reg_buffer_11458 ( .C (clk), .D (new_AGEMA_signal_32413), .Q (new_AGEMA_signal_32414) ) ;
    buf_clk new_AGEMA_reg_buffer_11462 ( .C (clk), .D (new_AGEMA_signal_32417), .Q (new_AGEMA_signal_32418) ) ;
    buf_clk new_AGEMA_reg_buffer_11466 ( .C (clk), .D (new_AGEMA_signal_32421), .Q (new_AGEMA_signal_32422) ) ;
    buf_clk new_AGEMA_reg_buffer_11470 ( .C (clk), .D (new_AGEMA_signal_32425), .Q (new_AGEMA_signal_32426) ) ;
    buf_clk new_AGEMA_reg_buffer_11474 ( .C (clk), .D (new_AGEMA_signal_32429), .Q (new_AGEMA_signal_32430) ) ;
    buf_clk new_AGEMA_reg_buffer_11478 ( .C (clk), .D (new_AGEMA_signal_32433), .Q (new_AGEMA_signal_32434) ) ;
    buf_clk new_AGEMA_reg_buffer_11482 ( .C (clk), .D (new_AGEMA_signal_32437), .Q (new_AGEMA_signal_32438) ) ;
    buf_clk new_AGEMA_reg_buffer_11486 ( .C (clk), .D (new_AGEMA_signal_32441), .Q (new_AGEMA_signal_32442) ) ;
    buf_clk new_AGEMA_reg_buffer_11490 ( .C (clk), .D (new_AGEMA_signal_32445), .Q (new_AGEMA_signal_32446) ) ;
    buf_clk new_AGEMA_reg_buffer_11494 ( .C (clk), .D (new_AGEMA_signal_32449), .Q (new_AGEMA_signal_32450) ) ;
    buf_clk new_AGEMA_reg_buffer_11498 ( .C (clk), .D (new_AGEMA_signal_32453), .Q (new_AGEMA_signal_32454) ) ;
    buf_clk new_AGEMA_reg_buffer_11502 ( .C (clk), .D (new_AGEMA_signal_32457), .Q (new_AGEMA_signal_32458) ) ;
    buf_clk new_AGEMA_reg_buffer_11506 ( .C (clk), .D (new_AGEMA_signal_32461), .Q (new_AGEMA_signal_32462) ) ;
    buf_clk new_AGEMA_reg_buffer_11510 ( .C (clk), .D (new_AGEMA_signal_32465), .Q (new_AGEMA_signal_32466) ) ;
    buf_clk new_AGEMA_reg_buffer_11514 ( .C (clk), .D (new_AGEMA_signal_32469), .Q (new_AGEMA_signal_32470) ) ;
    buf_clk new_AGEMA_reg_buffer_11518 ( .C (clk), .D (new_AGEMA_signal_32473), .Q (new_AGEMA_signal_32474) ) ;
    buf_clk new_AGEMA_reg_buffer_11522 ( .C (clk), .D (new_AGEMA_signal_32477), .Q (new_AGEMA_signal_32478) ) ;
    buf_clk new_AGEMA_reg_buffer_11526 ( .C (clk), .D (new_AGEMA_signal_32481), .Q (new_AGEMA_signal_32482) ) ;
    buf_clk new_AGEMA_reg_buffer_11530 ( .C (clk), .D (new_AGEMA_signal_32485), .Q (new_AGEMA_signal_32486) ) ;
    buf_clk new_AGEMA_reg_buffer_11534 ( .C (clk), .D (new_AGEMA_signal_32489), .Q (new_AGEMA_signal_32490) ) ;
    buf_clk new_AGEMA_reg_buffer_11538 ( .C (clk), .D (new_AGEMA_signal_32493), .Q (new_AGEMA_signal_32494) ) ;
    buf_clk new_AGEMA_reg_buffer_11542 ( .C (clk), .D (new_AGEMA_signal_32497), .Q (new_AGEMA_signal_32498) ) ;
    buf_clk new_AGEMA_reg_buffer_11546 ( .C (clk), .D (new_AGEMA_signal_32501), .Q (new_AGEMA_signal_32502) ) ;
    buf_clk new_AGEMA_reg_buffer_11550 ( .C (clk), .D (new_AGEMA_signal_32505), .Q (new_AGEMA_signal_32506) ) ;
    buf_clk new_AGEMA_reg_buffer_11554 ( .C (clk), .D (new_AGEMA_signal_32509), .Q (new_AGEMA_signal_32510) ) ;
    buf_clk new_AGEMA_reg_buffer_11558 ( .C (clk), .D (new_AGEMA_signal_32513), .Q (new_AGEMA_signal_32514) ) ;
    buf_clk new_AGEMA_reg_buffer_11562 ( .C (clk), .D (new_AGEMA_signal_32517), .Q (new_AGEMA_signal_32518) ) ;
    buf_clk new_AGEMA_reg_buffer_11566 ( .C (clk), .D (new_AGEMA_signal_32521), .Q (new_AGEMA_signal_32522) ) ;
    buf_clk new_AGEMA_reg_buffer_11570 ( .C (clk), .D (new_AGEMA_signal_32525), .Q (new_AGEMA_signal_32526) ) ;
    buf_clk new_AGEMA_reg_buffer_11574 ( .C (clk), .D (new_AGEMA_signal_32529), .Q (new_AGEMA_signal_32530) ) ;
    buf_clk new_AGEMA_reg_buffer_11578 ( .C (clk), .D (new_AGEMA_signal_32533), .Q (new_AGEMA_signal_32534) ) ;
    buf_clk new_AGEMA_reg_buffer_11582 ( .C (clk), .D (new_AGEMA_signal_32537), .Q (new_AGEMA_signal_32538) ) ;
    buf_clk new_AGEMA_reg_buffer_11586 ( .C (clk), .D (new_AGEMA_signal_32541), .Q (new_AGEMA_signal_32542) ) ;
    buf_clk new_AGEMA_reg_buffer_11590 ( .C (clk), .D (new_AGEMA_signal_32545), .Q (new_AGEMA_signal_32546) ) ;
    buf_clk new_AGEMA_reg_buffer_11594 ( .C (clk), .D (new_AGEMA_signal_32549), .Q (new_AGEMA_signal_32550) ) ;
    buf_clk new_AGEMA_reg_buffer_11598 ( .C (clk), .D (new_AGEMA_signal_32553), .Q (new_AGEMA_signal_32554) ) ;
    buf_clk new_AGEMA_reg_buffer_11602 ( .C (clk), .D (new_AGEMA_signal_32557), .Q (new_AGEMA_signal_32558) ) ;
    buf_clk new_AGEMA_reg_buffer_11606 ( .C (clk), .D (new_AGEMA_signal_32561), .Q (new_AGEMA_signal_32562) ) ;
    buf_clk new_AGEMA_reg_buffer_11610 ( .C (clk), .D (new_AGEMA_signal_32565), .Q (new_AGEMA_signal_32566) ) ;
    buf_clk new_AGEMA_reg_buffer_11614 ( .C (clk), .D (new_AGEMA_signal_32569), .Q (new_AGEMA_signal_32570) ) ;
    buf_clk new_AGEMA_reg_buffer_11618 ( .C (clk), .D (new_AGEMA_signal_32573), .Q (new_AGEMA_signal_32574) ) ;
    buf_clk new_AGEMA_reg_buffer_11622 ( .C (clk), .D (new_AGEMA_signal_32577), .Q (new_AGEMA_signal_32578) ) ;
    buf_clk new_AGEMA_reg_buffer_11626 ( .C (clk), .D (new_AGEMA_signal_32581), .Q (new_AGEMA_signal_32582) ) ;
    buf_clk new_AGEMA_reg_buffer_11630 ( .C (clk), .D (new_AGEMA_signal_32585), .Q (new_AGEMA_signal_32586) ) ;
    buf_clk new_AGEMA_reg_buffer_11634 ( .C (clk), .D (new_AGEMA_signal_32589), .Q (new_AGEMA_signal_32590) ) ;
    buf_clk new_AGEMA_reg_buffer_11638 ( .C (clk), .D (new_AGEMA_signal_32593), .Q (new_AGEMA_signal_32594) ) ;
    buf_clk new_AGEMA_reg_buffer_11642 ( .C (clk), .D (new_AGEMA_signal_32597), .Q (new_AGEMA_signal_32598) ) ;
    buf_clk new_AGEMA_reg_buffer_11646 ( .C (clk), .D (new_AGEMA_signal_32601), .Q (new_AGEMA_signal_32602) ) ;
    buf_clk new_AGEMA_reg_buffer_11650 ( .C (clk), .D (new_AGEMA_signal_32605), .Q (new_AGEMA_signal_32606) ) ;
    buf_clk new_AGEMA_reg_buffer_11654 ( .C (clk), .D (new_AGEMA_signal_32609), .Q (new_AGEMA_signal_32610) ) ;
    buf_clk new_AGEMA_reg_buffer_11658 ( .C (clk), .D (new_AGEMA_signal_32613), .Q (new_AGEMA_signal_32614) ) ;
    buf_clk new_AGEMA_reg_buffer_11662 ( .C (clk), .D (new_AGEMA_signal_32617), .Q (new_AGEMA_signal_32618) ) ;
    buf_clk new_AGEMA_reg_buffer_11666 ( .C (clk), .D (new_AGEMA_signal_32621), .Q (new_AGEMA_signal_32622) ) ;
    buf_clk new_AGEMA_reg_buffer_11670 ( .C (clk), .D (new_AGEMA_signal_32625), .Q (new_AGEMA_signal_32626) ) ;
    buf_clk new_AGEMA_reg_buffer_11674 ( .C (clk), .D (new_AGEMA_signal_32629), .Q (new_AGEMA_signal_32630) ) ;
    buf_clk new_AGEMA_reg_buffer_11678 ( .C (clk), .D (new_AGEMA_signal_32633), .Q (new_AGEMA_signal_32634) ) ;
    buf_clk new_AGEMA_reg_buffer_11682 ( .C (clk), .D (new_AGEMA_signal_32637), .Q (new_AGEMA_signal_32638) ) ;
    buf_clk new_AGEMA_reg_buffer_11686 ( .C (clk), .D (new_AGEMA_signal_32641), .Q (new_AGEMA_signal_32642) ) ;
    buf_clk new_AGEMA_reg_buffer_11690 ( .C (clk), .D (new_AGEMA_signal_32645), .Q (new_AGEMA_signal_32646) ) ;
    buf_clk new_AGEMA_reg_buffer_11694 ( .C (clk), .D (new_AGEMA_signal_32649), .Q (new_AGEMA_signal_32650) ) ;
    buf_clk new_AGEMA_reg_buffer_11698 ( .C (clk), .D (new_AGEMA_signal_32653), .Q (new_AGEMA_signal_32654) ) ;
    buf_clk new_AGEMA_reg_buffer_11702 ( .C (clk), .D (new_AGEMA_signal_32657), .Q (new_AGEMA_signal_32658) ) ;
    buf_clk new_AGEMA_reg_buffer_11706 ( .C (clk), .D (new_AGEMA_signal_32661), .Q (new_AGEMA_signal_32662) ) ;
    buf_clk new_AGEMA_reg_buffer_11710 ( .C (clk), .D (new_AGEMA_signal_32665), .Q (new_AGEMA_signal_32666) ) ;
    buf_clk new_AGEMA_reg_buffer_11714 ( .C (clk), .D (new_AGEMA_signal_32669), .Q (new_AGEMA_signal_32670) ) ;
    buf_clk new_AGEMA_reg_buffer_11718 ( .C (clk), .D (new_AGEMA_signal_32673), .Q (new_AGEMA_signal_32674) ) ;
    buf_clk new_AGEMA_reg_buffer_11722 ( .C (clk), .D (new_AGEMA_signal_32677), .Q (new_AGEMA_signal_32678) ) ;
    buf_clk new_AGEMA_reg_buffer_11726 ( .C (clk), .D (new_AGEMA_signal_32681), .Q (new_AGEMA_signal_32682) ) ;
    buf_clk new_AGEMA_reg_buffer_11730 ( .C (clk), .D (new_AGEMA_signal_32685), .Q (new_AGEMA_signal_32686) ) ;
    buf_clk new_AGEMA_reg_buffer_11734 ( .C (clk), .D (new_AGEMA_signal_32689), .Q (new_AGEMA_signal_32690) ) ;
    buf_clk new_AGEMA_reg_buffer_11738 ( .C (clk), .D (new_AGEMA_signal_32693), .Q (new_AGEMA_signal_32694) ) ;
    buf_clk new_AGEMA_reg_buffer_11742 ( .C (clk), .D (new_AGEMA_signal_32697), .Q (new_AGEMA_signal_32698) ) ;
    buf_clk new_AGEMA_reg_buffer_11746 ( .C (clk), .D (new_AGEMA_signal_32701), .Q (new_AGEMA_signal_32702) ) ;
    buf_clk new_AGEMA_reg_buffer_11750 ( .C (clk), .D (new_AGEMA_signal_32705), .Q (new_AGEMA_signal_32706) ) ;
    buf_clk new_AGEMA_reg_buffer_11754 ( .C (clk), .D (new_AGEMA_signal_32709), .Q (new_AGEMA_signal_32710) ) ;
    buf_clk new_AGEMA_reg_buffer_11758 ( .C (clk), .D (new_AGEMA_signal_32713), .Q (new_AGEMA_signal_32714) ) ;
    buf_clk new_AGEMA_reg_buffer_11762 ( .C (clk), .D (new_AGEMA_signal_32717), .Q (new_AGEMA_signal_32718) ) ;
    buf_clk new_AGEMA_reg_buffer_11766 ( .C (clk), .D (new_AGEMA_signal_32721), .Q (new_AGEMA_signal_32722) ) ;
    buf_clk new_AGEMA_reg_buffer_11770 ( .C (clk), .D (new_AGEMA_signal_32725), .Q (new_AGEMA_signal_32726) ) ;
    buf_clk new_AGEMA_reg_buffer_11774 ( .C (clk), .D (new_AGEMA_signal_32729), .Q (new_AGEMA_signal_32730) ) ;
    buf_clk new_AGEMA_reg_buffer_11778 ( .C (clk), .D (new_AGEMA_signal_32733), .Q (new_AGEMA_signal_32734) ) ;
    buf_clk new_AGEMA_reg_buffer_11782 ( .C (clk), .D (new_AGEMA_signal_32737), .Q (new_AGEMA_signal_32738) ) ;
    buf_clk new_AGEMA_reg_buffer_11786 ( .C (clk), .D (new_AGEMA_signal_32741), .Q (new_AGEMA_signal_32742) ) ;
    buf_clk new_AGEMA_reg_buffer_11790 ( .C (clk), .D (new_AGEMA_signal_32745), .Q (new_AGEMA_signal_32746) ) ;
    buf_clk new_AGEMA_reg_buffer_11794 ( .C (clk), .D (new_AGEMA_signal_32749), .Q (new_AGEMA_signal_32750) ) ;
    buf_clk new_AGEMA_reg_buffer_11798 ( .C (clk), .D (new_AGEMA_signal_32753), .Q (new_AGEMA_signal_32754) ) ;
    buf_clk new_AGEMA_reg_buffer_11802 ( .C (clk), .D (new_AGEMA_signal_32757), .Q (new_AGEMA_signal_32758) ) ;
    buf_clk new_AGEMA_reg_buffer_11806 ( .C (clk), .D (new_AGEMA_signal_32761), .Q (new_AGEMA_signal_32762) ) ;
    buf_clk new_AGEMA_reg_buffer_11810 ( .C (clk), .D (new_AGEMA_signal_32765), .Q (new_AGEMA_signal_32766) ) ;
    buf_clk new_AGEMA_reg_buffer_11814 ( .C (clk), .D (new_AGEMA_signal_32769), .Q (new_AGEMA_signal_32770) ) ;
    buf_clk new_AGEMA_reg_buffer_11818 ( .C (clk), .D (new_AGEMA_signal_32773), .Q (new_AGEMA_signal_32774) ) ;
    buf_clk new_AGEMA_reg_buffer_11822 ( .C (clk), .D (new_AGEMA_signal_32777), .Q (new_AGEMA_signal_32778) ) ;
    buf_clk new_AGEMA_reg_buffer_11826 ( .C (clk), .D (new_AGEMA_signal_32781), .Q (new_AGEMA_signal_32782) ) ;
    buf_clk new_AGEMA_reg_buffer_11830 ( .C (clk), .D (new_AGEMA_signal_32785), .Q (new_AGEMA_signal_32786) ) ;
    buf_clk new_AGEMA_reg_buffer_11834 ( .C (clk), .D (new_AGEMA_signal_32789), .Q (new_AGEMA_signal_32790) ) ;
    buf_clk new_AGEMA_reg_buffer_11838 ( .C (clk), .D (new_AGEMA_signal_32793), .Q (new_AGEMA_signal_32794) ) ;
    buf_clk new_AGEMA_reg_buffer_11842 ( .C (clk), .D (new_AGEMA_signal_32797), .Q (new_AGEMA_signal_32798) ) ;
    buf_clk new_AGEMA_reg_buffer_11846 ( .C (clk), .D (new_AGEMA_signal_32801), .Q (new_AGEMA_signal_32802) ) ;
    buf_clk new_AGEMA_reg_buffer_11850 ( .C (clk), .D (new_AGEMA_signal_32805), .Q (new_AGEMA_signal_32806) ) ;
    buf_clk new_AGEMA_reg_buffer_11854 ( .C (clk), .D (new_AGEMA_signal_32809), .Q (new_AGEMA_signal_32810) ) ;
    buf_clk new_AGEMA_reg_buffer_11858 ( .C (clk), .D (new_AGEMA_signal_32813), .Q (new_AGEMA_signal_32814) ) ;
    buf_clk new_AGEMA_reg_buffer_11862 ( .C (clk), .D (new_AGEMA_signal_32817), .Q (new_AGEMA_signal_32818) ) ;
    buf_clk new_AGEMA_reg_buffer_11866 ( .C (clk), .D (new_AGEMA_signal_32821), .Q (new_AGEMA_signal_32822) ) ;
    buf_clk new_AGEMA_reg_buffer_11870 ( .C (clk), .D (new_AGEMA_signal_32825), .Q (new_AGEMA_signal_32826) ) ;
    buf_clk new_AGEMA_reg_buffer_11874 ( .C (clk), .D (new_AGEMA_signal_32829), .Q (new_AGEMA_signal_32830) ) ;
    buf_clk new_AGEMA_reg_buffer_11878 ( .C (clk), .D (new_AGEMA_signal_32833), .Q (new_AGEMA_signal_32834) ) ;
    buf_clk new_AGEMA_reg_buffer_11882 ( .C (clk), .D (new_AGEMA_signal_32837), .Q (new_AGEMA_signal_32838) ) ;
    buf_clk new_AGEMA_reg_buffer_11886 ( .C (clk), .D (new_AGEMA_signal_32841), .Q (new_AGEMA_signal_32842) ) ;
    buf_clk new_AGEMA_reg_buffer_11890 ( .C (clk), .D (new_AGEMA_signal_32845), .Q (new_AGEMA_signal_32846) ) ;
    buf_clk new_AGEMA_reg_buffer_11894 ( .C (clk), .D (new_AGEMA_signal_32849), .Q (new_AGEMA_signal_32850) ) ;
    buf_clk new_AGEMA_reg_buffer_11898 ( .C (clk), .D (new_AGEMA_signal_32853), .Q (new_AGEMA_signal_32854) ) ;
    buf_clk new_AGEMA_reg_buffer_11902 ( .C (clk), .D (new_AGEMA_signal_32857), .Q (new_AGEMA_signal_32858) ) ;
    buf_clk new_AGEMA_reg_buffer_11906 ( .C (clk), .D (new_AGEMA_signal_32861), .Q (new_AGEMA_signal_32862) ) ;
    buf_clk new_AGEMA_reg_buffer_11910 ( .C (clk), .D (new_AGEMA_signal_32865), .Q (new_AGEMA_signal_32866) ) ;
    buf_clk new_AGEMA_reg_buffer_11914 ( .C (clk), .D (new_AGEMA_signal_32869), .Q (new_AGEMA_signal_32870) ) ;
    buf_clk new_AGEMA_reg_buffer_11918 ( .C (clk), .D (new_AGEMA_signal_32873), .Q (new_AGEMA_signal_32874) ) ;
    buf_clk new_AGEMA_reg_buffer_11922 ( .C (clk), .D (new_AGEMA_signal_32877), .Q (new_AGEMA_signal_32878) ) ;
    buf_clk new_AGEMA_reg_buffer_11926 ( .C (clk), .D (new_AGEMA_signal_32881), .Q (new_AGEMA_signal_32882) ) ;
    buf_clk new_AGEMA_reg_buffer_11930 ( .C (clk), .D (new_AGEMA_signal_32885), .Q (new_AGEMA_signal_32886) ) ;
    buf_clk new_AGEMA_reg_buffer_11934 ( .C (clk), .D (new_AGEMA_signal_32889), .Q (new_AGEMA_signal_32890) ) ;
    buf_clk new_AGEMA_reg_buffer_11938 ( .C (clk), .D (new_AGEMA_signal_32893), .Q (new_AGEMA_signal_32894) ) ;
    buf_clk new_AGEMA_reg_buffer_11942 ( .C (clk), .D (new_AGEMA_signal_32897), .Q (new_AGEMA_signal_32898) ) ;
    buf_clk new_AGEMA_reg_buffer_11946 ( .C (clk), .D (new_AGEMA_signal_32901), .Q (new_AGEMA_signal_32902) ) ;
    buf_clk new_AGEMA_reg_buffer_11950 ( .C (clk), .D (new_AGEMA_signal_32905), .Q (new_AGEMA_signal_32906) ) ;
    buf_clk new_AGEMA_reg_buffer_11954 ( .C (clk), .D (new_AGEMA_signal_32909), .Q (new_AGEMA_signal_32910) ) ;
    buf_clk new_AGEMA_reg_buffer_11958 ( .C (clk), .D (new_AGEMA_signal_32913), .Q (new_AGEMA_signal_32914) ) ;
    buf_clk new_AGEMA_reg_buffer_11962 ( .C (clk), .D (new_AGEMA_signal_32917), .Q (new_AGEMA_signal_32918) ) ;
    buf_clk new_AGEMA_reg_buffer_11966 ( .C (clk), .D (new_AGEMA_signal_32921), .Q (new_AGEMA_signal_32922) ) ;
    buf_clk new_AGEMA_reg_buffer_11970 ( .C (clk), .D (new_AGEMA_signal_32925), .Q (new_AGEMA_signal_32926) ) ;
    buf_clk new_AGEMA_reg_buffer_11974 ( .C (clk), .D (new_AGEMA_signal_32929), .Q (new_AGEMA_signal_32930) ) ;
    buf_clk new_AGEMA_reg_buffer_11978 ( .C (clk), .D (new_AGEMA_signal_32933), .Q (new_AGEMA_signal_32934) ) ;
    buf_clk new_AGEMA_reg_buffer_11982 ( .C (clk), .D (new_AGEMA_signal_32937), .Q (new_AGEMA_signal_32938) ) ;
    buf_clk new_AGEMA_reg_buffer_11986 ( .C (clk), .D (new_AGEMA_signal_32941), .Q (new_AGEMA_signal_32942) ) ;
    buf_clk new_AGEMA_reg_buffer_11990 ( .C (clk), .D (new_AGEMA_signal_32945), .Q (new_AGEMA_signal_32946) ) ;
    buf_clk new_AGEMA_reg_buffer_11994 ( .C (clk), .D (new_AGEMA_signal_32949), .Q (new_AGEMA_signal_32950) ) ;
    buf_clk new_AGEMA_reg_buffer_11998 ( .C (clk), .D (new_AGEMA_signal_32953), .Q (new_AGEMA_signal_32954) ) ;
    buf_clk new_AGEMA_reg_buffer_12002 ( .C (clk), .D (new_AGEMA_signal_32957), .Q (new_AGEMA_signal_32958) ) ;
    buf_clk new_AGEMA_reg_buffer_12006 ( .C (clk), .D (new_AGEMA_signal_32961), .Q (new_AGEMA_signal_32962) ) ;
    buf_clk new_AGEMA_reg_buffer_12010 ( .C (clk), .D (new_AGEMA_signal_32965), .Q (new_AGEMA_signal_32966) ) ;
    buf_clk new_AGEMA_reg_buffer_12014 ( .C (clk), .D (new_AGEMA_signal_32969), .Q (new_AGEMA_signal_32970) ) ;
    buf_clk new_AGEMA_reg_buffer_12018 ( .C (clk), .D (new_AGEMA_signal_32973), .Q (new_AGEMA_signal_32974) ) ;
    buf_clk new_AGEMA_reg_buffer_12022 ( .C (clk), .D (new_AGEMA_signal_32977), .Q (new_AGEMA_signal_32978) ) ;
    buf_clk new_AGEMA_reg_buffer_12026 ( .C (clk), .D (new_AGEMA_signal_32981), .Q (new_AGEMA_signal_32982) ) ;
    buf_clk new_AGEMA_reg_buffer_12030 ( .C (clk), .D (new_AGEMA_signal_32985), .Q (new_AGEMA_signal_32986) ) ;
    buf_clk new_AGEMA_reg_buffer_12034 ( .C (clk), .D (new_AGEMA_signal_32989), .Q (new_AGEMA_signal_32990) ) ;
    buf_clk new_AGEMA_reg_buffer_12038 ( .C (clk), .D (new_AGEMA_signal_32993), .Q (new_AGEMA_signal_32994) ) ;
    buf_clk new_AGEMA_reg_buffer_12042 ( .C (clk), .D (new_AGEMA_signal_32997), .Q (new_AGEMA_signal_32998) ) ;
    buf_clk new_AGEMA_reg_buffer_12046 ( .C (clk), .D (new_AGEMA_signal_33001), .Q (new_AGEMA_signal_33002) ) ;
    buf_clk new_AGEMA_reg_buffer_12050 ( .C (clk), .D (new_AGEMA_signal_33005), .Q (new_AGEMA_signal_33006) ) ;
    buf_clk new_AGEMA_reg_buffer_12054 ( .C (clk), .D (new_AGEMA_signal_33009), .Q (new_AGEMA_signal_33010) ) ;
    buf_clk new_AGEMA_reg_buffer_12058 ( .C (clk), .D (new_AGEMA_signal_33013), .Q (new_AGEMA_signal_33014) ) ;
    buf_clk new_AGEMA_reg_buffer_12062 ( .C (clk), .D (new_AGEMA_signal_33017), .Q (new_AGEMA_signal_33018) ) ;
    buf_clk new_AGEMA_reg_buffer_12066 ( .C (clk), .D (new_AGEMA_signal_33021), .Q (new_AGEMA_signal_33022) ) ;
    buf_clk new_AGEMA_reg_buffer_12070 ( .C (clk), .D (new_AGEMA_signal_33025), .Q (new_AGEMA_signal_33026) ) ;
    buf_clk new_AGEMA_reg_buffer_12074 ( .C (clk), .D (new_AGEMA_signal_33029), .Q (new_AGEMA_signal_33030) ) ;
    buf_clk new_AGEMA_reg_buffer_12078 ( .C (clk), .D (new_AGEMA_signal_33033), .Q (new_AGEMA_signal_33034) ) ;
    buf_clk new_AGEMA_reg_buffer_12082 ( .C (clk), .D (new_AGEMA_signal_33037), .Q (new_AGEMA_signal_33038) ) ;
    buf_clk new_AGEMA_reg_buffer_12086 ( .C (clk), .D (new_AGEMA_signal_33041), .Q (new_AGEMA_signal_33042) ) ;
    buf_clk new_AGEMA_reg_buffer_12090 ( .C (clk), .D (new_AGEMA_signal_33045), .Q (new_AGEMA_signal_33046) ) ;
    buf_clk new_AGEMA_reg_buffer_12094 ( .C (clk), .D (new_AGEMA_signal_33049), .Q (new_AGEMA_signal_33050) ) ;
    buf_clk new_AGEMA_reg_buffer_12098 ( .C (clk), .D (new_AGEMA_signal_33053), .Q (new_AGEMA_signal_33054) ) ;
    buf_clk new_AGEMA_reg_buffer_12102 ( .C (clk), .D (new_AGEMA_signal_33057), .Q (new_AGEMA_signal_33058) ) ;
    buf_clk new_AGEMA_reg_buffer_12106 ( .C (clk), .D (new_AGEMA_signal_33061), .Q (new_AGEMA_signal_33062) ) ;
    buf_clk new_AGEMA_reg_buffer_12110 ( .C (clk), .D (new_AGEMA_signal_33065), .Q (new_AGEMA_signal_33066) ) ;
    buf_clk new_AGEMA_reg_buffer_12114 ( .C (clk), .D (new_AGEMA_signal_33069), .Q (new_AGEMA_signal_33070) ) ;
    buf_clk new_AGEMA_reg_buffer_12118 ( .C (clk), .D (new_AGEMA_signal_33073), .Q (new_AGEMA_signal_33074) ) ;
    buf_clk new_AGEMA_reg_buffer_12122 ( .C (clk), .D (new_AGEMA_signal_33077), .Q (new_AGEMA_signal_33078) ) ;
    buf_clk new_AGEMA_reg_buffer_12126 ( .C (clk), .D (new_AGEMA_signal_33081), .Q (new_AGEMA_signal_33082) ) ;
    buf_clk new_AGEMA_reg_buffer_12130 ( .C (clk), .D (new_AGEMA_signal_33085), .Q (new_AGEMA_signal_33086) ) ;
    buf_clk new_AGEMA_reg_buffer_12134 ( .C (clk), .D (new_AGEMA_signal_33089), .Q (new_AGEMA_signal_33090) ) ;
    buf_clk new_AGEMA_reg_buffer_12138 ( .C (clk), .D (new_AGEMA_signal_33093), .Q (new_AGEMA_signal_33094) ) ;
    buf_clk new_AGEMA_reg_buffer_12142 ( .C (clk), .D (new_AGEMA_signal_33097), .Q (new_AGEMA_signal_33098) ) ;
    buf_clk new_AGEMA_reg_buffer_12146 ( .C (clk), .D (new_AGEMA_signal_33101), .Q (new_AGEMA_signal_33102) ) ;
    buf_clk new_AGEMA_reg_buffer_12150 ( .C (clk), .D (new_AGEMA_signal_33105), .Q (new_AGEMA_signal_33106) ) ;
    buf_clk new_AGEMA_reg_buffer_12154 ( .C (clk), .D (new_AGEMA_signal_33109), .Q (new_AGEMA_signal_33110) ) ;
    buf_clk new_AGEMA_reg_buffer_12158 ( .C (clk), .D (new_AGEMA_signal_33113), .Q (new_AGEMA_signal_33114) ) ;
    buf_clk new_AGEMA_reg_buffer_12162 ( .C (clk), .D (new_AGEMA_signal_33117), .Q (new_AGEMA_signal_33118) ) ;
    buf_clk new_AGEMA_reg_buffer_12166 ( .C (clk), .D (new_AGEMA_signal_33121), .Q (new_AGEMA_signal_33122) ) ;
    buf_clk new_AGEMA_reg_buffer_12170 ( .C (clk), .D (new_AGEMA_signal_33125), .Q (new_AGEMA_signal_33126) ) ;
    buf_clk new_AGEMA_reg_buffer_12174 ( .C (clk), .D (new_AGEMA_signal_33129), .Q (new_AGEMA_signal_33130) ) ;
    buf_clk new_AGEMA_reg_buffer_12178 ( .C (clk), .D (new_AGEMA_signal_33133), .Q (new_AGEMA_signal_33134) ) ;
    buf_clk new_AGEMA_reg_buffer_12182 ( .C (clk), .D (new_AGEMA_signal_33137), .Q (new_AGEMA_signal_33138) ) ;
    buf_clk new_AGEMA_reg_buffer_12186 ( .C (clk), .D (new_AGEMA_signal_33141), .Q (new_AGEMA_signal_33142) ) ;
    buf_clk new_AGEMA_reg_buffer_12190 ( .C (clk), .D (new_AGEMA_signal_33145), .Q (new_AGEMA_signal_33146) ) ;
    buf_clk new_AGEMA_reg_buffer_12194 ( .C (clk), .D (new_AGEMA_signal_33149), .Q (new_AGEMA_signal_33150) ) ;
    buf_clk new_AGEMA_reg_buffer_12198 ( .C (clk), .D (new_AGEMA_signal_33153), .Q (new_AGEMA_signal_33154) ) ;
    buf_clk new_AGEMA_reg_buffer_12202 ( .C (clk), .D (new_AGEMA_signal_33157), .Q (new_AGEMA_signal_33158) ) ;
    buf_clk new_AGEMA_reg_buffer_12206 ( .C (clk), .D (new_AGEMA_signal_33161), .Q (new_AGEMA_signal_33162) ) ;
    buf_clk new_AGEMA_reg_buffer_12210 ( .C (clk), .D (new_AGEMA_signal_33165), .Q (new_AGEMA_signal_33166) ) ;
    buf_clk new_AGEMA_reg_buffer_12214 ( .C (clk), .D (new_AGEMA_signal_33169), .Q (new_AGEMA_signal_33170) ) ;
    buf_clk new_AGEMA_reg_buffer_12218 ( .C (clk), .D (new_AGEMA_signal_33173), .Q (new_AGEMA_signal_33174) ) ;
    buf_clk new_AGEMA_reg_buffer_12222 ( .C (clk), .D (new_AGEMA_signal_33177), .Q (new_AGEMA_signal_33178) ) ;
    buf_clk new_AGEMA_reg_buffer_12226 ( .C (clk), .D (new_AGEMA_signal_33181), .Q (new_AGEMA_signal_33182) ) ;
    buf_clk new_AGEMA_reg_buffer_12230 ( .C (clk), .D (new_AGEMA_signal_33185), .Q (new_AGEMA_signal_33186) ) ;
    buf_clk new_AGEMA_reg_buffer_12234 ( .C (clk), .D (new_AGEMA_signal_33189), .Q (new_AGEMA_signal_33190) ) ;
    buf_clk new_AGEMA_reg_buffer_12238 ( .C (clk), .D (new_AGEMA_signal_33193), .Q (new_AGEMA_signal_33194) ) ;
    buf_clk new_AGEMA_reg_buffer_12242 ( .C (clk), .D (new_AGEMA_signal_33197), .Q (new_AGEMA_signal_33198) ) ;
    buf_clk new_AGEMA_reg_buffer_12246 ( .C (clk), .D (new_AGEMA_signal_33201), .Q (new_AGEMA_signal_33202) ) ;
    buf_clk new_AGEMA_reg_buffer_12250 ( .C (clk), .D (new_AGEMA_signal_33205), .Q (new_AGEMA_signal_33206) ) ;
    buf_clk new_AGEMA_reg_buffer_12254 ( .C (clk), .D (new_AGEMA_signal_33209), .Q (new_AGEMA_signal_33210) ) ;
    buf_clk new_AGEMA_reg_buffer_12258 ( .C (clk), .D (new_AGEMA_signal_33213), .Q (new_AGEMA_signal_33214) ) ;
    buf_clk new_AGEMA_reg_buffer_12262 ( .C (clk), .D (new_AGEMA_signal_33217), .Q (new_AGEMA_signal_33218) ) ;
    buf_clk new_AGEMA_reg_buffer_12266 ( .C (clk), .D (new_AGEMA_signal_33221), .Q (new_AGEMA_signal_33222) ) ;
    buf_clk new_AGEMA_reg_buffer_12270 ( .C (clk), .D (new_AGEMA_signal_33225), .Q (new_AGEMA_signal_33226) ) ;
    buf_clk new_AGEMA_reg_buffer_12274 ( .C (clk), .D (new_AGEMA_signal_33229), .Q (new_AGEMA_signal_33230) ) ;
    buf_clk new_AGEMA_reg_buffer_12278 ( .C (clk), .D (new_AGEMA_signal_33233), .Q (new_AGEMA_signal_33234) ) ;
    buf_clk new_AGEMA_reg_buffer_12282 ( .C (clk), .D (new_AGEMA_signal_33237), .Q (new_AGEMA_signal_33238) ) ;
    buf_clk new_AGEMA_reg_buffer_12286 ( .C (clk), .D (new_AGEMA_signal_33241), .Q (new_AGEMA_signal_33242) ) ;
    buf_clk new_AGEMA_reg_buffer_12290 ( .C (clk), .D (new_AGEMA_signal_33245), .Q (new_AGEMA_signal_33246) ) ;
    buf_clk new_AGEMA_reg_buffer_12294 ( .C (clk), .D (new_AGEMA_signal_33249), .Q (new_AGEMA_signal_33250) ) ;
    buf_clk new_AGEMA_reg_buffer_12298 ( .C (clk), .D (new_AGEMA_signal_33253), .Q (new_AGEMA_signal_33254) ) ;
    buf_clk new_AGEMA_reg_buffer_12302 ( .C (clk), .D (new_AGEMA_signal_33257), .Q (new_AGEMA_signal_33258) ) ;
    buf_clk new_AGEMA_reg_buffer_12306 ( .C (clk), .D (new_AGEMA_signal_33261), .Q (new_AGEMA_signal_33262) ) ;
    buf_clk new_AGEMA_reg_buffer_12310 ( .C (clk), .D (new_AGEMA_signal_33265), .Q (new_AGEMA_signal_33266) ) ;
    buf_clk new_AGEMA_reg_buffer_12314 ( .C (clk), .D (new_AGEMA_signal_33269), .Q (new_AGEMA_signal_33270) ) ;
    buf_clk new_AGEMA_reg_buffer_12318 ( .C (clk), .D (new_AGEMA_signal_33273), .Q (new_AGEMA_signal_33274) ) ;
    buf_clk new_AGEMA_reg_buffer_12322 ( .C (clk), .D (new_AGEMA_signal_33277), .Q (new_AGEMA_signal_33278) ) ;
    buf_clk new_AGEMA_reg_buffer_12326 ( .C (clk), .D (new_AGEMA_signal_33281), .Q (new_AGEMA_signal_33282) ) ;
    buf_clk new_AGEMA_reg_buffer_12330 ( .C (clk), .D (new_AGEMA_signal_33285), .Q (new_AGEMA_signal_33286) ) ;
    buf_clk new_AGEMA_reg_buffer_12334 ( .C (clk), .D (new_AGEMA_signal_33289), .Q (new_AGEMA_signal_33290) ) ;
    buf_clk new_AGEMA_reg_buffer_12338 ( .C (clk), .D (new_AGEMA_signal_33293), .Q (new_AGEMA_signal_33294) ) ;
    buf_clk new_AGEMA_reg_buffer_12342 ( .C (clk), .D (new_AGEMA_signal_33297), .Q (new_AGEMA_signal_33298) ) ;
    buf_clk new_AGEMA_reg_buffer_12346 ( .C (clk), .D (new_AGEMA_signal_33301), .Q (new_AGEMA_signal_33302) ) ;
    buf_clk new_AGEMA_reg_buffer_12350 ( .C (clk), .D (new_AGEMA_signal_33305), .Q (new_AGEMA_signal_33306) ) ;
    buf_clk new_AGEMA_reg_buffer_12354 ( .C (clk), .D (new_AGEMA_signal_33309), .Q (new_AGEMA_signal_33310) ) ;
    buf_clk new_AGEMA_reg_buffer_12358 ( .C (clk), .D (new_AGEMA_signal_33313), .Q (new_AGEMA_signal_33314) ) ;
    buf_clk new_AGEMA_reg_buffer_12362 ( .C (clk), .D (new_AGEMA_signal_33317), .Q (new_AGEMA_signal_33318) ) ;
    buf_clk new_AGEMA_reg_buffer_12366 ( .C (clk), .D (new_AGEMA_signal_33321), .Q (new_AGEMA_signal_33322) ) ;
    buf_clk new_AGEMA_reg_buffer_12370 ( .C (clk), .D (new_AGEMA_signal_33325), .Q (new_AGEMA_signal_33326) ) ;
    buf_clk new_AGEMA_reg_buffer_12374 ( .C (clk), .D (new_AGEMA_signal_33329), .Q (new_AGEMA_signal_33330) ) ;
    buf_clk new_AGEMA_reg_buffer_12378 ( .C (clk), .D (new_AGEMA_signal_33333), .Q (new_AGEMA_signal_33334) ) ;
    buf_clk new_AGEMA_reg_buffer_12382 ( .C (clk), .D (new_AGEMA_signal_33337), .Q (new_AGEMA_signal_33338) ) ;
    buf_clk new_AGEMA_reg_buffer_12386 ( .C (clk), .D (new_AGEMA_signal_33341), .Q (new_AGEMA_signal_33342) ) ;
    buf_clk new_AGEMA_reg_buffer_12390 ( .C (clk), .D (new_AGEMA_signal_33345), .Q (new_AGEMA_signal_33346) ) ;
    buf_clk new_AGEMA_reg_buffer_12394 ( .C (clk), .D (new_AGEMA_signal_33349), .Q (new_AGEMA_signal_33350) ) ;
    buf_clk new_AGEMA_reg_buffer_12398 ( .C (clk), .D (new_AGEMA_signal_33353), .Q (new_AGEMA_signal_33354) ) ;
    buf_clk new_AGEMA_reg_buffer_12402 ( .C (clk), .D (new_AGEMA_signal_33357), .Q (new_AGEMA_signal_33358) ) ;
    buf_clk new_AGEMA_reg_buffer_12406 ( .C (clk), .D (new_AGEMA_signal_33361), .Q (new_AGEMA_signal_33362) ) ;
    buf_clk new_AGEMA_reg_buffer_12410 ( .C (clk), .D (new_AGEMA_signal_33365), .Q (new_AGEMA_signal_33366) ) ;
    buf_clk new_AGEMA_reg_buffer_12414 ( .C (clk), .D (new_AGEMA_signal_33369), .Q (new_AGEMA_signal_33370) ) ;
    buf_clk new_AGEMA_reg_buffer_12418 ( .C (clk), .D (new_AGEMA_signal_33373), .Q (new_AGEMA_signal_33374) ) ;
    buf_clk new_AGEMA_reg_buffer_12422 ( .C (clk), .D (new_AGEMA_signal_33377), .Q (new_AGEMA_signal_33378) ) ;
    buf_clk new_AGEMA_reg_buffer_12426 ( .C (clk), .D (new_AGEMA_signal_33381), .Q (new_AGEMA_signal_33382) ) ;
    buf_clk new_AGEMA_reg_buffer_12430 ( .C (clk), .D (new_AGEMA_signal_33385), .Q (new_AGEMA_signal_33386) ) ;
    buf_clk new_AGEMA_reg_buffer_12434 ( .C (clk), .D (new_AGEMA_signal_33389), .Q (new_AGEMA_signal_33390) ) ;
    buf_clk new_AGEMA_reg_buffer_12438 ( .C (clk), .D (new_AGEMA_signal_33393), .Q (new_AGEMA_signal_33394) ) ;
    buf_clk new_AGEMA_reg_buffer_12442 ( .C (clk), .D (new_AGEMA_signal_33397), .Q (new_AGEMA_signal_33398) ) ;
    buf_clk new_AGEMA_reg_buffer_12446 ( .C (clk), .D (new_AGEMA_signal_33401), .Q (new_AGEMA_signal_33402) ) ;
    buf_clk new_AGEMA_reg_buffer_12450 ( .C (clk), .D (new_AGEMA_signal_33405), .Q (new_AGEMA_signal_33406) ) ;
    buf_clk new_AGEMA_reg_buffer_12454 ( .C (clk), .D (new_AGEMA_signal_33409), .Q (new_AGEMA_signal_33410) ) ;
    buf_clk new_AGEMA_reg_buffer_12458 ( .C (clk), .D (new_AGEMA_signal_33413), .Q (new_AGEMA_signal_33414) ) ;
    buf_clk new_AGEMA_reg_buffer_12462 ( .C (clk), .D (new_AGEMA_signal_33417), .Q (new_AGEMA_signal_33418) ) ;
    buf_clk new_AGEMA_reg_buffer_12466 ( .C (clk), .D (new_AGEMA_signal_33421), .Q (new_AGEMA_signal_33422) ) ;
    buf_clk new_AGEMA_reg_buffer_12470 ( .C (clk), .D (new_AGEMA_signal_33425), .Q (new_AGEMA_signal_33426) ) ;
    buf_clk new_AGEMA_reg_buffer_12474 ( .C (clk), .D (new_AGEMA_signal_33429), .Q (new_AGEMA_signal_33430) ) ;
    buf_clk new_AGEMA_reg_buffer_12478 ( .C (clk), .D (new_AGEMA_signal_33433), .Q (new_AGEMA_signal_33434) ) ;
    buf_clk new_AGEMA_reg_buffer_12482 ( .C (clk), .D (new_AGEMA_signal_33437), .Q (new_AGEMA_signal_33438) ) ;
    buf_clk new_AGEMA_reg_buffer_12486 ( .C (clk), .D (new_AGEMA_signal_33441), .Q (new_AGEMA_signal_33442) ) ;
    buf_clk new_AGEMA_reg_buffer_12490 ( .C (clk), .D (new_AGEMA_signal_33445), .Q (new_AGEMA_signal_33446) ) ;
    buf_clk new_AGEMA_reg_buffer_12494 ( .C (clk), .D (new_AGEMA_signal_33449), .Q (new_AGEMA_signal_33450) ) ;
    buf_clk new_AGEMA_reg_buffer_12498 ( .C (clk), .D (new_AGEMA_signal_33453), .Q (new_AGEMA_signal_33454) ) ;
    buf_clk new_AGEMA_reg_buffer_12502 ( .C (clk), .D (new_AGEMA_signal_33457), .Q (new_AGEMA_signal_33458) ) ;
    buf_clk new_AGEMA_reg_buffer_12506 ( .C (clk), .D (new_AGEMA_signal_33461), .Q (new_AGEMA_signal_33462) ) ;
    buf_clk new_AGEMA_reg_buffer_12510 ( .C (clk), .D (new_AGEMA_signal_33465), .Q (new_AGEMA_signal_33466) ) ;
    buf_clk new_AGEMA_reg_buffer_12514 ( .C (clk), .D (new_AGEMA_signal_33469), .Q (new_AGEMA_signal_33470) ) ;
    buf_clk new_AGEMA_reg_buffer_12518 ( .C (clk), .D (new_AGEMA_signal_33473), .Q (new_AGEMA_signal_33474) ) ;
    buf_clk new_AGEMA_reg_buffer_12522 ( .C (clk), .D (new_AGEMA_signal_33477), .Q (new_AGEMA_signal_33478) ) ;
    buf_clk new_AGEMA_reg_buffer_12526 ( .C (clk), .D (new_AGEMA_signal_33481), .Q (new_AGEMA_signal_33482) ) ;
    buf_clk new_AGEMA_reg_buffer_12530 ( .C (clk), .D (new_AGEMA_signal_33485), .Q (new_AGEMA_signal_33486) ) ;
    buf_clk new_AGEMA_reg_buffer_12534 ( .C (clk), .D (new_AGEMA_signal_33489), .Q (new_AGEMA_signal_33490) ) ;
    buf_clk new_AGEMA_reg_buffer_12538 ( .C (clk), .D (new_AGEMA_signal_33493), .Q (new_AGEMA_signal_33494) ) ;
    buf_clk new_AGEMA_reg_buffer_12542 ( .C (clk), .D (new_AGEMA_signal_33497), .Q (new_AGEMA_signal_33498) ) ;
    buf_clk new_AGEMA_reg_buffer_12546 ( .C (clk), .D (new_AGEMA_signal_33501), .Q (new_AGEMA_signal_33502) ) ;
    buf_clk new_AGEMA_reg_buffer_12550 ( .C (clk), .D (new_AGEMA_signal_33505), .Q (new_AGEMA_signal_33506) ) ;
    buf_clk new_AGEMA_reg_buffer_12554 ( .C (clk), .D (new_AGEMA_signal_33509), .Q (new_AGEMA_signal_33510) ) ;
    buf_clk new_AGEMA_reg_buffer_12558 ( .C (clk), .D (new_AGEMA_signal_33513), .Q (new_AGEMA_signal_33514) ) ;
    buf_clk new_AGEMA_reg_buffer_12562 ( .C (clk), .D (new_AGEMA_signal_33517), .Q (new_AGEMA_signal_33518) ) ;
    buf_clk new_AGEMA_reg_buffer_12566 ( .C (clk), .D (new_AGEMA_signal_33521), .Q (new_AGEMA_signal_33522) ) ;
    buf_clk new_AGEMA_reg_buffer_12570 ( .C (clk), .D (new_AGEMA_signal_33525), .Q (new_AGEMA_signal_33526) ) ;
    buf_clk new_AGEMA_reg_buffer_12574 ( .C (clk), .D (new_AGEMA_signal_33529), .Q (new_AGEMA_signal_33530) ) ;
    buf_clk new_AGEMA_reg_buffer_12578 ( .C (clk), .D (new_AGEMA_signal_33533), .Q (new_AGEMA_signal_33534) ) ;
    buf_clk new_AGEMA_reg_buffer_12582 ( .C (clk), .D (new_AGEMA_signal_33537), .Q (new_AGEMA_signal_33538) ) ;
    buf_clk new_AGEMA_reg_buffer_12586 ( .C (clk), .D (new_AGEMA_signal_33541), .Q (new_AGEMA_signal_33542) ) ;
    buf_clk new_AGEMA_reg_buffer_12590 ( .C (clk), .D (new_AGEMA_signal_33545), .Q (new_AGEMA_signal_33546) ) ;
    buf_clk new_AGEMA_reg_buffer_12594 ( .C (clk), .D (new_AGEMA_signal_33549), .Q (new_AGEMA_signal_33550) ) ;
    buf_clk new_AGEMA_reg_buffer_12598 ( .C (clk), .D (new_AGEMA_signal_33553), .Q (new_AGEMA_signal_33554) ) ;
    buf_clk new_AGEMA_reg_buffer_12602 ( .C (clk), .D (new_AGEMA_signal_33557), .Q (new_AGEMA_signal_33558) ) ;
    buf_clk new_AGEMA_reg_buffer_12606 ( .C (clk), .D (new_AGEMA_signal_33561), .Q (new_AGEMA_signal_33562) ) ;
    buf_clk new_AGEMA_reg_buffer_12610 ( .C (clk), .D (new_AGEMA_signal_33565), .Q (new_AGEMA_signal_33566) ) ;
    buf_clk new_AGEMA_reg_buffer_12614 ( .C (clk), .D (new_AGEMA_signal_33569), .Q (new_AGEMA_signal_33570) ) ;
    buf_clk new_AGEMA_reg_buffer_12618 ( .C (clk), .D (new_AGEMA_signal_33573), .Q (new_AGEMA_signal_33574) ) ;
    buf_clk new_AGEMA_reg_buffer_12622 ( .C (clk), .D (new_AGEMA_signal_33577), .Q (new_AGEMA_signal_33578) ) ;
    buf_clk new_AGEMA_reg_buffer_12626 ( .C (clk), .D (new_AGEMA_signal_33581), .Q (new_AGEMA_signal_33582) ) ;
    buf_clk new_AGEMA_reg_buffer_12630 ( .C (clk), .D (new_AGEMA_signal_33585), .Q (new_AGEMA_signal_33586) ) ;
    buf_clk new_AGEMA_reg_buffer_12634 ( .C (clk), .D (new_AGEMA_signal_33589), .Q (new_AGEMA_signal_33590) ) ;
    buf_clk new_AGEMA_reg_buffer_12638 ( .C (clk), .D (new_AGEMA_signal_33593), .Q (new_AGEMA_signal_33594) ) ;
    buf_clk new_AGEMA_reg_buffer_12642 ( .C (clk), .D (new_AGEMA_signal_33597), .Q (new_AGEMA_signal_33598) ) ;
    buf_clk new_AGEMA_reg_buffer_12646 ( .C (clk), .D (new_AGEMA_signal_33601), .Q (new_AGEMA_signal_33602) ) ;
    buf_clk new_AGEMA_reg_buffer_12650 ( .C (clk), .D (new_AGEMA_signal_33605), .Q (new_AGEMA_signal_33606) ) ;
    buf_clk new_AGEMA_reg_buffer_12654 ( .C (clk), .D (new_AGEMA_signal_33609), .Q (new_AGEMA_signal_33610) ) ;
    buf_clk new_AGEMA_reg_buffer_12658 ( .C (clk), .D (new_AGEMA_signal_33613), .Q (new_AGEMA_signal_33614) ) ;
    buf_clk new_AGEMA_reg_buffer_12662 ( .C (clk), .D (new_AGEMA_signal_33617), .Q (new_AGEMA_signal_33618) ) ;
    buf_clk new_AGEMA_reg_buffer_12666 ( .C (clk), .D (new_AGEMA_signal_33621), .Q (new_AGEMA_signal_33622) ) ;
    buf_clk new_AGEMA_reg_buffer_12670 ( .C (clk), .D (new_AGEMA_signal_33625), .Q (new_AGEMA_signal_33626) ) ;
    buf_clk new_AGEMA_reg_buffer_12674 ( .C (clk), .D (new_AGEMA_signal_33629), .Q (new_AGEMA_signal_33630) ) ;
    buf_clk new_AGEMA_reg_buffer_12678 ( .C (clk), .D (new_AGEMA_signal_33633), .Q (new_AGEMA_signal_33634) ) ;
    buf_clk new_AGEMA_reg_buffer_12682 ( .C (clk), .D (new_AGEMA_signal_33637), .Q (new_AGEMA_signal_33638) ) ;
    buf_clk new_AGEMA_reg_buffer_12686 ( .C (clk), .D (new_AGEMA_signal_33641), .Q (new_AGEMA_signal_33642) ) ;
    buf_clk new_AGEMA_reg_buffer_12690 ( .C (clk), .D (new_AGEMA_signal_33645), .Q (new_AGEMA_signal_33646) ) ;
    buf_clk new_AGEMA_reg_buffer_12694 ( .C (clk), .D (new_AGEMA_signal_33649), .Q (new_AGEMA_signal_33650) ) ;
    buf_clk new_AGEMA_reg_buffer_12698 ( .C (clk), .D (new_AGEMA_signal_33653), .Q (new_AGEMA_signal_33654) ) ;
    buf_clk new_AGEMA_reg_buffer_12702 ( .C (clk), .D (new_AGEMA_signal_33657), .Q (new_AGEMA_signal_33658) ) ;
    buf_clk new_AGEMA_reg_buffer_12706 ( .C (clk), .D (new_AGEMA_signal_33661), .Q (new_AGEMA_signal_33662) ) ;
    buf_clk new_AGEMA_reg_buffer_12710 ( .C (clk), .D (new_AGEMA_signal_33665), .Q (new_AGEMA_signal_33666) ) ;
    buf_clk new_AGEMA_reg_buffer_12714 ( .C (clk), .D (new_AGEMA_signal_33669), .Q (new_AGEMA_signal_33670) ) ;
    buf_clk new_AGEMA_reg_buffer_12718 ( .C (clk), .D (new_AGEMA_signal_33673), .Q (new_AGEMA_signal_33674) ) ;
    buf_clk new_AGEMA_reg_buffer_12722 ( .C (clk), .D (new_AGEMA_signal_33677), .Q (new_AGEMA_signal_33678) ) ;
    buf_clk new_AGEMA_reg_buffer_12726 ( .C (clk), .D (new_AGEMA_signal_33681), .Q (new_AGEMA_signal_33682) ) ;
    buf_clk new_AGEMA_reg_buffer_12730 ( .C (clk), .D (new_AGEMA_signal_33685), .Q (new_AGEMA_signal_33686) ) ;
    buf_clk new_AGEMA_reg_buffer_12734 ( .C (clk), .D (new_AGEMA_signal_33689), .Q (new_AGEMA_signal_33690) ) ;
    buf_clk new_AGEMA_reg_buffer_12738 ( .C (clk), .D (new_AGEMA_signal_33693), .Q (new_AGEMA_signal_33694) ) ;
    buf_clk new_AGEMA_reg_buffer_12742 ( .C (clk), .D (new_AGEMA_signal_33697), .Q (new_AGEMA_signal_33698) ) ;
    buf_clk new_AGEMA_reg_buffer_12746 ( .C (clk), .D (new_AGEMA_signal_33701), .Q (new_AGEMA_signal_33702) ) ;
    buf_clk new_AGEMA_reg_buffer_12750 ( .C (clk), .D (new_AGEMA_signal_33705), .Q (new_AGEMA_signal_33706) ) ;
    buf_clk new_AGEMA_reg_buffer_12754 ( .C (clk), .D (new_AGEMA_signal_33709), .Q (new_AGEMA_signal_33710) ) ;
    buf_clk new_AGEMA_reg_buffer_12758 ( .C (clk), .D (new_AGEMA_signal_33713), .Q (new_AGEMA_signal_33714) ) ;
    buf_clk new_AGEMA_reg_buffer_12762 ( .C (clk), .D (new_AGEMA_signal_33717), .Q (new_AGEMA_signal_33718) ) ;
    buf_clk new_AGEMA_reg_buffer_12766 ( .C (clk), .D (new_AGEMA_signal_33721), .Q (new_AGEMA_signal_33722) ) ;
    buf_clk new_AGEMA_reg_buffer_12770 ( .C (clk), .D (new_AGEMA_signal_33725), .Q (new_AGEMA_signal_33726) ) ;
    buf_clk new_AGEMA_reg_buffer_12774 ( .C (clk), .D (new_AGEMA_signal_33729), .Q (new_AGEMA_signal_33730) ) ;
    buf_clk new_AGEMA_reg_buffer_12778 ( .C (clk), .D (new_AGEMA_signal_33733), .Q (new_AGEMA_signal_33734) ) ;
    buf_clk new_AGEMA_reg_buffer_12782 ( .C (clk), .D (new_AGEMA_signal_33737), .Q (new_AGEMA_signal_33738) ) ;
    buf_clk new_AGEMA_reg_buffer_12786 ( .C (clk), .D (new_AGEMA_signal_33741), .Q (new_AGEMA_signal_33742) ) ;
    buf_clk new_AGEMA_reg_buffer_12790 ( .C (clk), .D (new_AGEMA_signal_33745), .Q (new_AGEMA_signal_33746) ) ;
    buf_clk new_AGEMA_reg_buffer_12794 ( .C (clk), .D (new_AGEMA_signal_33749), .Q (new_AGEMA_signal_33750) ) ;
    buf_clk new_AGEMA_reg_buffer_12798 ( .C (clk), .D (new_AGEMA_signal_33753), .Q (new_AGEMA_signal_33754) ) ;
    buf_clk new_AGEMA_reg_buffer_12802 ( .C (clk), .D (new_AGEMA_signal_33757), .Q (new_AGEMA_signal_33758) ) ;
    buf_clk new_AGEMA_reg_buffer_12806 ( .C (clk), .D (new_AGEMA_signal_33761), .Q (new_AGEMA_signal_33762) ) ;
    buf_clk new_AGEMA_reg_buffer_12810 ( .C (clk), .D (new_AGEMA_signal_33765), .Q (new_AGEMA_signal_33766) ) ;
    buf_clk new_AGEMA_reg_buffer_12814 ( .C (clk), .D (new_AGEMA_signal_33769), .Q (new_AGEMA_signal_33770) ) ;
    buf_clk new_AGEMA_reg_buffer_12818 ( .C (clk), .D (new_AGEMA_signal_33773), .Q (new_AGEMA_signal_33774) ) ;
    buf_clk new_AGEMA_reg_buffer_12822 ( .C (clk), .D (new_AGEMA_signal_33777), .Q (new_AGEMA_signal_33778) ) ;
    buf_clk new_AGEMA_reg_buffer_12826 ( .C (clk), .D (new_AGEMA_signal_33781), .Q (new_AGEMA_signal_33782) ) ;
    buf_clk new_AGEMA_reg_buffer_12830 ( .C (clk), .D (new_AGEMA_signal_33785), .Q (new_AGEMA_signal_33786) ) ;
    buf_clk new_AGEMA_reg_buffer_12834 ( .C (clk), .D (new_AGEMA_signal_33789), .Q (new_AGEMA_signal_33790) ) ;
    buf_clk new_AGEMA_reg_buffer_12838 ( .C (clk), .D (new_AGEMA_signal_33793), .Q (new_AGEMA_signal_33794) ) ;
    buf_clk new_AGEMA_reg_buffer_12842 ( .C (clk), .D (new_AGEMA_signal_33797), .Q (new_AGEMA_signal_33798) ) ;
    buf_clk new_AGEMA_reg_buffer_12846 ( .C (clk), .D (new_AGEMA_signal_33801), .Q (new_AGEMA_signal_33802) ) ;
    buf_clk new_AGEMA_reg_buffer_12850 ( .C (clk), .D (new_AGEMA_signal_33805), .Q (new_AGEMA_signal_33806) ) ;
    buf_clk new_AGEMA_reg_buffer_12854 ( .C (clk), .D (new_AGEMA_signal_33809), .Q (new_AGEMA_signal_33810) ) ;
    buf_clk new_AGEMA_reg_buffer_12858 ( .C (clk), .D (new_AGEMA_signal_33813), .Q (new_AGEMA_signal_33814) ) ;
    buf_clk new_AGEMA_reg_buffer_12862 ( .C (clk), .D (new_AGEMA_signal_33817), .Q (new_AGEMA_signal_33818) ) ;
    buf_clk new_AGEMA_reg_buffer_12866 ( .C (clk), .D (new_AGEMA_signal_33821), .Q (new_AGEMA_signal_33822) ) ;
    buf_clk new_AGEMA_reg_buffer_12870 ( .C (clk), .D (new_AGEMA_signal_33825), .Q (new_AGEMA_signal_33826) ) ;
    buf_clk new_AGEMA_reg_buffer_12874 ( .C (clk), .D (new_AGEMA_signal_33829), .Q (new_AGEMA_signal_33830) ) ;
    buf_clk new_AGEMA_reg_buffer_12878 ( .C (clk), .D (new_AGEMA_signal_33833), .Q (new_AGEMA_signal_33834) ) ;
    buf_clk new_AGEMA_reg_buffer_12882 ( .C (clk), .D (new_AGEMA_signal_33837), .Q (new_AGEMA_signal_33838) ) ;
    buf_clk new_AGEMA_reg_buffer_12886 ( .C (clk), .D (new_AGEMA_signal_33841), .Q (new_AGEMA_signal_33842) ) ;
    buf_clk new_AGEMA_reg_buffer_12890 ( .C (clk), .D (new_AGEMA_signal_33845), .Q (new_AGEMA_signal_33846) ) ;
    buf_clk new_AGEMA_reg_buffer_12894 ( .C (clk), .D (new_AGEMA_signal_33849), .Q (new_AGEMA_signal_33850) ) ;
    buf_clk new_AGEMA_reg_buffer_12898 ( .C (clk), .D (new_AGEMA_signal_33853), .Q (new_AGEMA_signal_33854) ) ;
    buf_clk new_AGEMA_reg_buffer_12902 ( .C (clk), .D (new_AGEMA_signal_33857), .Q (new_AGEMA_signal_33858) ) ;
    buf_clk new_AGEMA_reg_buffer_12906 ( .C (clk), .D (new_AGEMA_signal_33861), .Q (new_AGEMA_signal_33862) ) ;
    buf_clk new_AGEMA_reg_buffer_12910 ( .C (clk), .D (new_AGEMA_signal_33865), .Q (new_AGEMA_signal_33866) ) ;
    buf_clk new_AGEMA_reg_buffer_12914 ( .C (clk), .D (new_AGEMA_signal_33869), .Q (new_AGEMA_signal_33870) ) ;
    buf_clk new_AGEMA_reg_buffer_12918 ( .C (clk), .D (new_AGEMA_signal_33873), .Q (new_AGEMA_signal_33874) ) ;
    buf_clk new_AGEMA_reg_buffer_12922 ( .C (clk), .D (new_AGEMA_signal_33877), .Q (new_AGEMA_signal_33878) ) ;
    buf_clk new_AGEMA_reg_buffer_12926 ( .C (clk), .D (new_AGEMA_signal_33881), .Q (new_AGEMA_signal_33882) ) ;
    buf_clk new_AGEMA_reg_buffer_12930 ( .C (clk), .D (new_AGEMA_signal_33885), .Q (new_AGEMA_signal_33886) ) ;
    buf_clk new_AGEMA_reg_buffer_12934 ( .C (clk), .D (new_AGEMA_signal_33889), .Q (new_AGEMA_signal_33890) ) ;
    buf_clk new_AGEMA_reg_buffer_12938 ( .C (clk), .D (new_AGEMA_signal_33893), .Q (new_AGEMA_signal_33894) ) ;
    buf_clk new_AGEMA_reg_buffer_12942 ( .C (clk), .D (new_AGEMA_signal_33897), .Q (new_AGEMA_signal_33898) ) ;
    buf_clk new_AGEMA_reg_buffer_12946 ( .C (clk), .D (new_AGEMA_signal_33901), .Q (new_AGEMA_signal_33902) ) ;
    buf_clk new_AGEMA_reg_buffer_12950 ( .C (clk), .D (new_AGEMA_signal_33905), .Q (new_AGEMA_signal_33906) ) ;
    buf_clk new_AGEMA_reg_buffer_12954 ( .C (clk), .D (new_AGEMA_signal_33909), .Q (new_AGEMA_signal_33910) ) ;
    buf_clk new_AGEMA_reg_buffer_12958 ( .C (clk), .D (new_AGEMA_signal_33913), .Q (new_AGEMA_signal_33914) ) ;
    buf_clk new_AGEMA_reg_buffer_12962 ( .C (clk), .D (new_AGEMA_signal_33917), .Q (new_AGEMA_signal_33918) ) ;
    buf_clk new_AGEMA_reg_buffer_12966 ( .C (clk), .D (new_AGEMA_signal_33921), .Q (new_AGEMA_signal_33922) ) ;
    buf_clk new_AGEMA_reg_buffer_12970 ( .C (clk), .D (new_AGEMA_signal_33925), .Q (new_AGEMA_signal_33926) ) ;
    buf_clk new_AGEMA_reg_buffer_12974 ( .C (clk), .D (new_AGEMA_signal_33929), .Q (new_AGEMA_signal_33930) ) ;
    buf_clk new_AGEMA_reg_buffer_12978 ( .C (clk), .D (new_AGEMA_signal_33933), .Q (new_AGEMA_signal_33934) ) ;
    buf_clk new_AGEMA_reg_buffer_12982 ( .C (clk), .D (new_AGEMA_signal_33937), .Q (new_AGEMA_signal_33938) ) ;
    buf_clk new_AGEMA_reg_buffer_12986 ( .C (clk), .D (new_AGEMA_signal_33941), .Q (new_AGEMA_signal_33942) ) ;
    buf_clk new_AGEMA_reg_buffer_12990 ( .C (clk), .D (new_AGEMA_signal_33945), .Q (new_AGEMA_signal_33946) ) ;
    buf_clk new_AGEMA_reg_buffer_12994 ( .C (clk), .D (new_AGEMA_signal_33949), .Q (new_AGEMA_signal_33950) ) ;
    buf_clk new_AGEMA_reg_buffer_12998 ( .C (clk), .D (new_AGEMA_signal_33953), .Q (new_AGEMA_signal_33954) ) ;
    buf_clk new_AGEMA_reg_buffer_13002 ( .C (clk), .D (new_AGEMA_signal_33957), .Q (new_AGEMA_signal_33958) ) ;
    buf_clk new_AGEMA_reg_buffer_13006 ( .C (clk), .D (new_AGEMA_signal_33961), .Q (new_AGEMA_signal_33962) ) ;
    buf_clk new_AGEMA_reg_buffer_13010 ( .C (clk), .D (new_AGEMA_signal_33965), .Q (new_AGEMA_signal_33966) ) ;
    buf_clk new_AGEMA_reg_buffer_13014 ( .C (clk), .D (new_AGEMA_signal_33969), .Q (new_AGEMA_signal_33970) ) ;
    buf_clk new_AGEMA_reg_buffer_13018 ( .C (clk), .D (new_AGEMA_signal_33973), .Q (new_AGEMA_signal_33974) ) ;
    buf_clk new_AGEMA_reg_buffer_13022 ( .C (clk), .D (new_AGEMA_signal_33977), .Q (new_AGEMA_signal_33978) ) ;
    buf_clk new_AGEMA_reg_buffer_13026 ( .C (clk), .D (new_AGEMA_signal_33981), .Q (new_AGEMA_signal_33982) ) ;
    buf_clk new_AGEMA_reg_buffer_13030 ( .C (clk), .D (new_AGEMA_signal_33985), .Q (new_AGEMA_signal_33986) ) ;
    buf_clk new_AGEMA_reg_buffer_13034 ( .C (clk), .D (new_AGEMA_signal_33989), .Q (new_AGEMA_signal_33990) ) ;
    buf_clk new_AGEMA_reg_buffer_13038 ( .C (clk), .D (new_AGEMA_signal_33993), .Q (new_AGEMA_signal_33994) ) ;
    buf_clk new_AGEMA_reg_buffer_13042 ( .C (clk), .D (new_AGEMA_signal_33997), .Q (new_AGEMA_signal_33998) ) ;
    buf_clk new_AGEMA_reg_buffer_13046 ( .C (clk), .D (new_AGEMA_signal_34001), .Q (new_AGEMA_signal_34002) ) ;
    buf_clk new_AGEMA_reg_buffer_13050 ( .C (clk), .D (new_AGEMA_signal_34005), .Q (new_AGEMA_signal_34006) ) ;
    buf_clk new_AGEMA_reg_buffer_13054 ( .C (clk), .D (new_AGEMA_signal_34009), .Q (new_AGEMA_signal_34010) ) ;
    buf_clk new_AGEMA_reg_buffer_13058 ( .C (clk), .D (new_AGEMA_signal_34013), .Q (new_AGEMA_signal_34014) ) ;
    buf_clk new_AGEMA_reg_buffer_13062 ( .C (clk), .D (new_AGEMA_signal_34017), .Q (new_AGEMA_signal_34018) ) ;
    buf_clk new_AGEMA_reg_buffer_13066 ( .C (clk), .D (new_AGEMA_signal_34021), .Q (new_AGEMA_signal_34022) ) ;
    buf_clk new_AGEMA_reg_buffer_13070 ( .C (clk), .D (new_AGEMA_signal_34025), .Q (new_AGEMA_signal_34026) ) ;
    buf_clk new_AGEMA_reg_buffer_13074 ( .C (clk), .D (new_AGEMA_signal_34029), .Q (new_AGEMA_signal_34030) ) ;
    buf_clk new_AGEMA_reg_buffer_13078 ( .C (clk), .D (new_AGEMA_signal_34033), .Q (new_AGEMA_signal_34034) ) ;
    buf_clk new_AGEMA_reg_buffer_13082 ( .C (clk), .D (new_AGEMA_signal_34037), .Q (new_AGEMA_signal_34038) ) ;
    buf_clk new_AGEMA_reg_buffer_13086 ( .C (clk), .D (new_AGEMA_signal_34041), .Q (new_AGEMA_signal_34042) ) ;
    buf_clk new_AGEMA_reg_buffer_13090 ( .C (clk), .D (new_AGEMA_signal_34045), .Q (new_AGEMA_signal_34046) ) ;
    buf_clk new_AGEMA_reg_buffer_13094 ( .C (clk), .D (new_AGEMA_signal_34049), .Q (new_AGEMA_signal_34050) ) ;
    buf_clk new_AGEMA_reg_buffer_13098 ( .C (clk), .D (new_AGEMA_signal_34053), .Q (new_AGEMA_signal_34054) ) ;
    buf_clk new_AGEMA_reg_buffer_13102 ( .C (clk), .D (new_AGEMA_signal_34057), .Q (new_AGEMA_signal_34058) ) ;
    buf_clk new_AGEMA_reg_buffer_13106 ( .C (clk), .D (new_AGEMA_signal_34061), .Q (new_AGEMA_signal_34062) ) ;
    buf_clk new_AGEMA_reg_buffer_13110 ( .C (clk), .D (new_AGEMA_signal_34065), .Q (new_AGEMA_signal_34066) ) ;
    buf_clk new_AGEMA_reg_buffer_13114 ( .C (clk), .D (new_AGEMA_signal_34069), .Q (new_AGEMA_signal_34070) ) ;
    buf_clk new_AGEMA_reg_buffer_13118 ( .C (clk), .D (new_AGEMA_signal_34073), .Q (new_AGEMA_signal_34074) ) ;
    buf_clk new_AGEMA_reg_buffer_13122 ( .C (clk), .D (new_AGEMA_signal_34077), .Q (new_AGEMA_signal_34078) ) ;
    buf_clk new_AGEMA_reg_buffer_13126 ( .C (clk), .D (new_AGEMA_signal_34081), .Q (new_AGEMA_signal_34082) ) ;
    buf_clk new_AGEMA_reg_buffer_13130 ( .C (clk), .D (new_AGEMA_signal_34085), .Q (new_AGEMA_signal_34086) ) ;
    buf_clk new_AGEMA_reg_buffer_13134 ( .C (clk), .D (new_AGEMA_signal_34089), .Q (new_AGEMA_signal_34090) ) ;
    buf_clk new_AGEMA_reg_buffer_13138 ( .C (clk), .D (new_AGEMA_signal_34093), .Q (new_AGEMA_signal_34094) ) ;
    buf_clk new_AGEMA_reg_buffer_13142 ( .C (clk), .D (new_AGEMA_signal_34097), .Q (new_AGEMA_signal_34098) ) ;
    buf_clk new_AGEMA_reg_buffer_13146 ( .C (clk), .D (new_AGEMA_signal_34101), .Q (new_AGEMA_signal_34102) ) ;
    buf_clk new_AGEMA_reg_buffer_13150 ( .C (clk), .D (new_AGEMA_signal_34105), .Q (new_AGEMA_signal_34106) ) ;
    buf_clk new_AGEMA_reg_buffer_13154 ( .C (clk), .D (new_AGEMA_signal_34109), .Q (new_AGEMA_signal_34110) ) ;
    buf_clk new_AGEMA_reg_buffer_13158 ( .C (clk), .D (new_AGEMA_signal_34113), .Q (new_AGEMA_signal_34114) ) ;
    buf_clk new_AGEMA_reg_buffer_13162 ( .C (clk), .D (new_AGEMA_signal_34117), .Q (new_AGEMA_signal_34118) ) ;
    buf_clk new_AGEMA_reg_buffer_13166 ( .C (clk), .D (new_AGEMA_signal_34121), .Q (new_AGEMA_signal_34122) ) ;
    buf_clk new_AGEMA_reg_buffer_13170 ( .C (clk), .D (new_AGEMA_signal_34125), .Q (new_AGEMA_signal_34126) ) ;
    buf_clk new_AGEMA_reg_buffer_13174 ( .C (clk), .D (new_AGEMA_signal_34129), .Q (new_AGEMA_signal_34130) ) ;
    buf_clk new_AGEMA_reg_buffer_13178 ( .C (clk), .D (new_AGEMA_signal_34133), .Q (new_AGEMA_signal_34134) ) ;
    buf_clk new_AGEMA_reg_buffer_13182 ( .C (clk), .D (new_AGEMA_signal_34137), .Q (new_AGEMA_signal_34138) ) ;
    buf_clk new_AGEMA_reg_buffer_13186 ( .C (clk), .D (new_AGEMA_signal_34141), .Q (new_AGEMA_signal_34142) ) ;
    buf_clk new_AGEMA_reg_buffer_13190 ( .C (clk), .D (new_AGEMA_signal_34145), .Q (new_AGEMA_signal_34146) ) ;
    buf_clk new_AGEMA_reg_buffer_13194 ( .C (clk), .D (new_AGEMA_signal_34149), .Q (new_AGEMA_signal_34150) ) ;
    buf_clk new_AGEMA_reg_buffer_13198 ( .C (clk), .D (new_AGEMA_signal_34153), .Q (new_AGEMA_signal_34154) ) ;
    buf_clk new_AGEMA_reg_buffer_13202 ( .C (clk), .D (new_AGEMA_signal_34157), .Q (new_AGEMA_signal_34158) ) ;
    buf_clk new_AGEMA_reg_buffer_13206 ( .C (clk), .D (new_AGEMA_signal_34161), .Q (new_AGEMA_signal_34162) ) ;
    buf_clk new_AGEMA_reg_buffer_13210 ( .C (clk), .D (new_AGEMA_signal_34165), .Q (new_AGEMA_signal_34166) ) ;
    buf_clk new_AGEMA_reg_buffer_13214 ( .C (clk), .D (new_AGEMA_signal_34169), .Q (new_AGEMA_signal_34170) ) ;
    buf_clk new_AGEMA_reg_buffer_13218 ( .C (clk), .D (new_AGEMA_signal_34173), .Q (new_AGEMA_signal_34174) ) ;
    buf_clk new_AGEMA_reg_buffer_13222 ( .C (clk), .D (new_AGEMA_signal_34177), .Q (new_AGEMA_signal_34178) ) ;
    buf_clk new_AGEMA_reg_buffer_13226 ( .C (clk), .D (new_AGEMA_signal_34181), .Q (new_AGEMA_signal_34182) ) ;
    buf_clk new_AGEMA_reg_buffer_13230 ( .C (clk), .D (new_AGEMA_signal_34185), .Q (new_AGEMA_signal_34186) ) ;
    buf_clk new_AGEMA_reg_buffer_13234 ( .C (clk), .D (new_AGEMA_signal_34189), .Q (new_AGEMA_signal_34190) ) ;
    buf_clk new_AGEMA_reg_buffer_13238 ( .C (clk), .D (new_AGEMA_signal_34193), .Q (new_AGEMA_signal_34194) ) ;
    buf_clk new_AGEMA_reg_buffer_13242 ( .C (clk), .D (new_AGEMA_signal_34197), .Q (new_AGEMA_signal_34198) ) ;
    buf_clk new_AGEMA_reg_buffer_13246 ( .C (clk), .D (new_AGEMA_signal_34201), .Q (new_AGEMA_signal_34202) ) ;
    buf_clk new_AGEMA_reg_buffer_13250 ( .C (clk), .D (new_AGEMA_signal_34205), .Q (new_AGEMA_signal_34206) ) ;
    buf_clk new_AGEMA_reg_buffer_13254 ( .C (clk), .D (new_AGEMA_signal_34209), .Q (new_AGEMA_signal_34210) ) ;
    buf_clk new_AGEMA_reg_buffer_13258 ( .C (clk), .D (new_AGEMA_signal_34213), .Q (new_AGEMA_signal_34214) ) ;
    buf_clk new_AGEMA_reg_buffer_13262 ( .C (clk), .D (new_AGEMA_signal_34217), .Q (new_AGEMA_signal_34218) ) ;
    buf_clk new_AGEMA_reg_buffer_13266 ( .C (clk), .D (new_AGEMA_signal_34221), .Q (new_AGEMA_signal_34222) ) ;
    buf_clk new_AGEMA_reg_buffer_13270 ( .C (clk), .D (new_AGEMA_signal_34225), .Q (new_AGEMA_signal_34226) ) ;
    buf_clk new_AGEMA_reg_buffer_13274 ( .C (clk), .D (new_AGEMA_signal_34229), .Q (new_AGEMA_signal_34230) ) ;
    buf_clk new_AGEMA_reg_buffer_13278 ( .C (clk), .D (new_AGEMA_signal_34233), .Q (new_AGEMA_signal_34234) ) ;
    buf_clk new_AGEMA_reg_buffer_13282 ( .C (clk), .D (new_AGEMA_signal_34237), .Q (new_AGEMA_signal_34238) ) ;
    buf_clk new_AGEMA_reg_buffer_13286 ( .C (clk), .D (new_AGEMA_signal_34241), .Q (new_AGEMA_signal_34242) ) ;
    buf_clk new_AGEMA_reg_buffer_13290 ( .C (clk), .D (new_AGEMA_signal_34245), .Q (new_AGEMA_signal_34246) ) ;
    buf_clk new_AGEMA_reg_buffer_13294 ( .C (clk), .D (new_AGEMA_signal_34249), .Q (new_AGEMA_signal_34250) ) ;
    buf_clk new_AGEMA_reg_buffer_13298 ( .C (clk), .D (new_AGEMA_signal_34253), .Q (new_AGEMA_signal_34254) ) ;
    buf_clk new_AGEMA_reg_buffer_13302 ( .C (clk), .D (new_AGEMA_signal_34257), .Q (new_AGEMA_signal_34258) ) ;
    buf_clk new_AGEMA_reg_buffer_13306 ( .C (clk), .D (new_AGEMA_signal_34261), .Q (new_AGEMA_signal_34262) ) ;
    buf_clk new_AGEMA_reg_buffer_13310 ( .C (clk), .D (new_AGEMA_signal_34265), .Q (new_AGEMA_signal_34266) ) ;
    buf_clk new_AGEMA_reg_buffer_13314 ( .C (clk), .D (new_AGEMA_signal_34269), .Q (new_AGEMA_signal_34270) ) ;
    buf_clk new_AGEMA_reg_buffer_13318 ( .C (clk), .D (new_AGEMA_signal_34273), .Q (new_AGEMA_signal_34274) ) ;
    buf_clk new_AGEMA_reg_buffer_13322 ( .C (clk), .D (new_AGEMA_signal_34277), .Q (new_AGEMA_signal_34278) ) ;
    buf_clk new_AGEMA_reg_buffer_13326 ( .C (clk), .D (new_AGEMA_signal_34281), .Q (new_AGEMA_signal_34282) ) ;
    buf_clk new_AGEMA_reg_buffer_13330 ( .C (clk), .D (new_AGEMA_signal_34285), .Q (new_AGEMA_signal_34286) ) ;
    buf_clk new_AGEMA_reg_buffer_13334 ( .C (clk), .D (new_AGEMA_signal_34289), .Q (new_AGEMA_signal_34290) ) ;
    buf_clk new_AGEMA_reg_buffer_13338 ( .C (clk), .D (new_AGEMA_signal_34293), .Q (new_AGEMA_signal_34294) ) ;
    buf_clk new_AGEMA_reg_buffer_13342 ( .C (clk), .D (new_AGEMA_signal_34297), .Q (new_AGEMA_signal_34298) ) ;
    buf_clk new_AGEMA_reg_buffer_13346 ( .C (clk), .D (new_AGEMA_signal_34301), .Q (new_AGEMA_signal_34302) ) ;
    buf_clk new_AGEMA_reg_buffer_13350 ( .C (clk), .D (new_AGEMA_signal_34305), .Q (new_AGEMA_signal_34306) ) ;
    buf_clk new_AGEMA_reg_buffer_13354 ( .C (clk), .D (new_AGEMA_signal_34309), .Q (new_AGEMA_signal_34310) ) ;
    buf_clk new_AGEMA_reg_buffer_13358 ( .C (clk), .D (new_AGEMA_signal_34313), .Q (new_AGEMA_signal_34314) ) ;
    buf_clk new_AGEMA_reg_buffer_13362 ( .C (clk), .D (new_AGEMA_signal_34317), .Q (new_AGEMA_signal_34318) ) ;
    buf_clk new_AGEMA_reg_buffer_13366 ( .C (clk), .D (new_AGEMA_signal_34321), .Q (new_AGEMA_signal_34322) ) ;
    buf_clk new_AGEMA_reg_buffer_13370 ( .C (clk), .D (new_AGEMA_signal_34325), .Q (new_AGEMA_signal_34326) ) ;
    buf_clk new_AGEMA_reg_buffer_13374 ( .C (clk), .D (new_AGEMA_signal_34329), .Q (new_AGEMA_signal_34330) ) ;
    buf_clk new_AGEMA_reg_buffer_13378 ( .C (clk), .D (new_AGEMA_signal_34333), .Q (new_AGEMA_signal_34334) ) ;
    buf_clk new_AGEMA_reg_buffer_13382 ( .C (clk), .D (new_AGEMA_signal_34337), .Q (new_AGEMA_signal_34338) ) ;
    buf_clk new_AGEMA_reg_buffer_13386 ( .C (clk), .D (new_AGEMA_signal_34341), .Q (new_AGEMA_signal_34342) ) ;
    buf_clk new_AGEMA_reg_buffer_13390 ( .C (clk), .D (new_AGEMA_signal_34345), .Q (new_AGEMA_signal_34346) ) ;
    buf_clk new_AGEMA_reg_buffer_13394 ( .C (clk), .D (new_AGEMA_signal_34349), .Q (new_AGEMA_signal_34350) ) ;
    buf_clk new_AGEMA_reg_buffer_13398 ( .C (clk), .D (new_AGEMA_signal_34353), .Q (new_AGEMA_signal_34354) ) ;
    buf_clk new_AGEMA_reg_buffer_13402 ( .C (clk), .D (new_AGEMA_signal_34357), .Q (new_AGEMA_signal_34358) ) ;
    buf_clk new_AGEMA_reg_buffer_13406 ( .C (clk), .D (new_AGEMA_signal_34361), .Q (new_AGEMA_signal_34362) ) ;
    buf_clk new_AGEMA_reg_buffer_13410 ( .C (clk), .D (new_AGEMA_signal_34365), .Q (new_AGEMA_signal_34366) ) ;
    buf_clk new_AGEMA_reg_buffer_13414 ( .C (clk), .D (new_AGEMA_signal_34369), .Q (new_AGEMA_signal_34370) ) ;
    buf_clk new_AGEMA_reg_buffer_13418 ( .C (clk), .D (new_AGEMA_signal_34373), .Q (new_AGEMA_signal_34374) ) ;
    buf_clk new_AGEMA_reg_buffer_13422 ( .C (clk), .D (new_AGEMA_signal_34377), .Q (new_AGEMA_signal_34378) ) ;
    buf_clk new_AGEMA_reg_buffer_13426 ( .C (clk), .D (new_AGEMA_signal_34381), .Q (new_AGEMA_signal_34382) ) ;
    buf_clk new_AGEMA_reg_buffer_13430 ( .C (clk), .D (new_AGEMA_signal_34385), .Q (new_AGEMA_signal_34386) ) ;
    buf_clk new_AGEMA_reg_buffer_13434 ( .C (clk), .D (new_AGEMA_signal_34389), .Q (new_AGEMA_signal_34390) ) ;
    buf_clk new_AGEMA_reg_buffer_13438 ( .C (clk), .D (new_AGEMA_signal_34393), .Q (new_AGEMA_signal_34394) ) ;
    buf_clk new_AGEMA_reg_buffer_13442 ( .C (clk), .D (new_AGEMA_signal_34397), .Q (new_AGEMA_signal_34398) ) ;
    buf_clk new_AGEMA_reg_buffer_13446 ( .C (clk), .D (new_AGEMA_signal_34401), .Q (new_AGEMA_signal_34402) ) ;
    buf_clk new_AGEMA_reg_buffer_13450 ( .C (clk), .D (new_AGEMA_signal_34405), .Q (new_AGEMA_signal_34406) ) ;
    buf_clk new_AGEMA_reg_buffer_13454 ( .C (clk), .D (new_AGEMA_signal_34409), .Q (new_AGEMA_signal_34410) ) ;
    buf_clk new_AGEMA_reg_buffer_13458 ( .C (clk), .D (new_AGEMA_signal_34413), .Q (new_AGEMA_signal_34414) ) ;
    buf_clk new_AGEMA_reg_buffer_13462 ( .C (clk), .D (new_AGEMA_signal_34417), .Q (new_AGEMA_signal_34418) ) ;
    buf_clk new_AGEMA_reg_buffer_13466 ( .C (clk), .D (new_AGEMA_signal_34421), .Q (new_AGEMA_signal_34422) ) ;
    buf_clk new_AGEMA_reg_buffer_13470 ( .C (clk), .D (new_AGEMA_signal_34425), .Q (new_AGEMA_signal_34426) ) ;
    buf_clk new_AGEMA_reg_buffer_13474 ( .C (clk), .D (new_AGEMA_signal_34429), .Q (new_AGEMA_signal_34430) ) ;
    buf_clk new_AGEMA_reg_buffer_13478 ( .C (clk), .D (new_AGEMA_signal_34433), .Q (new_AGEMA_signal_34434) ) ;
    buf_clk new_AGEMA_reg_buffer_13482 ( .C (clk), .D (new_AGEMA_signal_34437), .Q (new_AGEMA_signal_34438) ) ;
    buf_clk new_AGEMA_reg_buffer_13486 ( .C (clk), .D (new_AGEMA_signal_34441), .Q (new_AGEMA_signal_34442) ) ;
    buf_clk new_AGEMA_reg_buffer_13490 ( .C (clk), .D (new_AGEMA_signal_34445), .Q (new_AGEMA_signal_34446) ) ;
    buf_clk new_AGEMA_reg_buffer_13494 ( .C (clk), .D (new_AGEMA_signal_34449), .Q (new_AGEMA_signal_34450) ) ;
    buf_clk new_AGEMA_reg_buffer_13498 ( .C (clk), .D (new_AGEMA_signal_34453), .Q (new_AGEMA_signal_34454) ) ;
    buf_clk new_AGEMA_reg_buffer_13502 ( .C (clk), .D (new_AGEMA_signal_34457), .Q (new_AGEMA_signal_34458) ) ;
    buf_clk new_AGEMA_reg_buffer_13506 ( .C (clk), .D (new_AGEMA_signal_34461), .Q (new_AGEMA_signal_34462) ) ;
    buf_clk new_AGEMA_reg_buffer_13510 ( .C (clk), .D (new_AGEMA_signal_34465), .Q (new_AGEMA_signal_34466) ) ;
    buf_clk new_AGEMA_reg_buffer_13514 ( .C (clk), .D (new_AGEMA_signal_34469), .Q (new_AGEMA_signal_34470) ) ;
    buf_clk new_AGEMA_reg_buffer_13518 ( .C (clk), .D (new_AGEMA_signal_34473), .Q (new_AGEMA_signal_34474) ) ;
    buf_clk new_AGEMA_reg_buffer_13522 ( .C (clk), .D (new_AGEMA_signal_34477), .Q (new_AGEMA_signal_34478) ) ;
    buf_clk new_AGEMA_reg_buffer_13526 ( .C (clk), .D (new_AGEMA_signal_34481), .Q (new_AGEMA_signal_34482) ) ;
    buf_clk new_AGEMA_reg_buffer_13530 ( .C (clk), .D (new_AGEMA_signal_34485), .Q (new_AGEMA_signal_34486) ) ;
    buf_clk new_AGEMA_reg_buffer_13534 ( .C (clk), .D (new_AGEMA_signal_34489), .Q (new_AGEMA_signal_34490) ) ;
    buf_clk new_AGEMA_reg_buffer_13538 ( .C (clk), .D (new_AGEMA_signal_34493), .Q (new_AGEMA_signal_34494) ) ;
    buf_clk new_AGEMA_reg_buffer_13542 ( .C (clk), .D (new_AGEMA_signal_34497), .Q (new_AGEMA_signal_34498) ) ;
    buf_clk new_AGEMA_reg_buffer_13546 ( .C (clk), .D (new_AGEMA_signal_34501), .Q (new_AGEMA_signal_34502) ) ;
    buf_clk new_AGEMA_reg_buffer_13550 ( .C (clk), .D (new_AGEMA_signal_34505), .Q (new_AGEMA_signal_34506) ) ;
    buf_clk new_AGEMA_reg_buffer_13554 ( .C (clk), .D (new_AGEMA_signal_34509), .Q (new_AGEMA_signal_34510) ) ;
    buf_clk new_AGEMA_reg_buffer_13558 ( .C (clk), .D (new_AGEMA_signal_34513), .Q (new_AGEMA_signal_34514) ) ;
    buf_clk new_AGEMA_reg_buffer_13562 ( .C (clk), .D (new_AGEMA_signal_34517), .Q (new_AGEMA_signal_34518) ) ;
    buf_clk new_AGEMA_reg_buffer_13566 ( .C (clk), .D (new_AGEMA_signal_34521), .Q (new_AGEMA_signal_34522) ) ;
    buf_clk new_AGEMA_reg_buffer_13570 ( .C (clk), .D (new_AGEMA_signal_34525), .Q (new_AGEMA_signal_34526) ) ;
    buf_clk new_AGEMA_reg_buffer_13574 ( .C (clk), .D (new_AGEMA_signal_34529), .Q (new_AGEMA_signal_34530) ) ;
    buf_clk new_AGEMA_reg_buffer_13578 ( .C (clk), .D (new_AGEMA_signal_34533), .Q (new_AGEMA_signal_34534) ) ;
    buf_clk new_AGEMA_reg_buffer_13582 ( .C (clk), .D (new_AGEMA_signal_34537), .Q (new_AGEMA_signal_34538) ) ;
    buf_clk new_AGEMA_reg_buffer_13586 ( .C (clk), .D (new_AGEMA_signal_34541), .Q (new_AGEMA_signal_34542) ) ;
    buf_clk new_AGEMA_reg_buffer_13590 ( .C (clk), .D (new_AGEMA_signal_34545), .Q (new_AGEMA_signal_34546) ) ;
    buf_clk new_AGEMA_reg_buffer_13594 ( .C (clk), .D (new_AGEMA_signal_34549), .Q (new_AGEMA_signal_34550) ) ;
    buf_clk new_AGEMA_reg_buffer_13598 ( .C (clk), .D (new_AGEMA_signal_34553), .Q (new_AGEMA_signal_34554) ) ;
    buf_clk new_AGEMA_reg_buffer_13602 ( .C (clk), .D (new_AGEMA_signal_34557), .Q (new_AGEMA_signal_34558) ) ;
    buf_clk new_AGEMA_reg_buffer_13606 ( .C (clk), .D (new_AGEMA_signal_34561), .Q (new_AGEMA_signal_34562) ) ;
    buf_clk new_AGEMA_reg_buffer_13610 ( .C (clk), .D (new_AGEMA_signal_34565), .Q (new_AGEMA_signal_34566) ) ;
    buf_clk new_AGEMA_reg_buffer_13614 ( .C (clk), .D (new_AGEMA_signal_34569), .Q (new_AGEMA_signal_34570) ) ;
    buf_clk new_AGEMA_reg_buffer_13618 ( .C (clk), .D (new_AGEMA_signal_34573), .Q (new_AGEMA_signal_34574) ) ;
    buf_clk new_AGEMA_reg_buffer_13622 ( .C (clk), .D (new_AGEMA_signal_34577), .Q (new_AGEMA_signal_34578) ) ;
    buf_clk new_AGEMA_reg_buffer_13626 ( .C (clk), .D (new_AGEMA_signal_34581), .Q (new_AGEMA_signal_34582) ) ;
    buf_clk new_AGEMA_reg_buffer_13630 ( .C (clk), .D (new_AGEMA_signal_34585), .Q (new_AGEMA_signal_34586) ) ;
    buf_clk new_AGEMA_reg_buffer_13634 ( .C (clk), .D (new_AGEMA_signal_34589), .Q (new_AGEMA_signal_34590) ) ;
    buf_clk new_AGEMA_reg_buffer_13638 ( .C (clk), .D (new_AGEMA_signal_34593), .Q (new_AGEMA_signal_34594) ) ;
    buf_clk new_AGEMA_reg_buffer_13642 ( .C (clk), .D (new_AGEMA_signal_34597), .Q (new_AGEMA_signal_34598) ) ;
    buf_clk new_AGEMA_reg_buffer_13646 ( .C (clk), .D (new_AGEMA_signal_34601), .Q (new_AGEMA_signal_34602) ) ;
    buf_clk new_AGEMA_reg_buffer_13650 ( .C (clk), .D (new_AGEMA_signal_34605), .Q (new_AGEMA_signal_34606) ) ;
    buf_clk new_AGEMA_reg_buffer_13654 ( .C (clk), .D (new_AGEMA_signal_34609), .Q (new_AGEMA_signal_34610) ) ;
    buf_clk new_AGEMA_reg_buffer_13658 ( .C (clk), .D (new_AGEMA_signal_34613), .Q (new_AGEMA_signal_34614) ) ;
    buf_clk new_AGEMA_reg_buffer_13662 ( .C (clk), .D (new_AGEMA_signal_34617), .Q (new_AGEMA_signal_34618) ) ;
    buf_clk new_AGEMA_reg_buffer_13666 ( .C (clk), .D (new_AGEMA_signal_34621), .Q (new_AGEMA_signal_34622) ) ;
    buf_clk new_AGEMA_reg_buffer_13670 ( .C (clk), .D (new_AGEMA_signal_34625), .Q (new_AGEMA_signal_34626) ) ;
    buf_clk new_AGEMA_reg_buffer_13674 ( .C (clk), .D (new_AGEMA_signal_34629), .Q (new_AGEMA_signal_34630) ) ;
    buf_clk new_AGEMA_reg_buffer_13678 ( .C (clk), .D (new_AGEMA_signal_34633), .Q (new_AGEMA_signal_34634) ) ;
    buf_clk new_AGEMA_reg_buffer_13682 ( .C (clk), .D (new_AGEMA_signal_34637), .Q (new_AGEMA_signal_34638) ) ;
    buf_clk new_AGEMA_reg_buffer_13686 ( .C (clk), .D (new_AGEMA_signal_34641), .Q (new_AGEMA_signal_34642) ) ;
    buf_clk new_AGEMA_reg_buffer_13690 ( .C (clk), .D (new_AGEMA_signal_34645), .Q (new_AGEMA_signal_34646) ) ;
    buf_clk new_AGEMA_reg_buffer_13694 ( .C (clk), .D (new_AGEMA_signal_34649), .Q (new_AGEMA_signal_34650) ) ;
    buf_clk new_AGEMA_reg_buffer_13698 ( .C (clk), .D (new_AGEMA_signal_34653), .Q (new_AGEMA_signal_34654) ) ;
    buf_clk new_AGEMA_reg_buffer_13702 ( .C (clk), .D (new_AGEMA_signal_34657), .Q (new_AGEMA_signal_34658) ) ;
    buf_clk new_AGEMA_reg_buffer_13706 ( .C (clk), .D (new_AGEMA_signal_34661), .Q (new_AGEMA_signal_34662) ) ;
    buf_clk new_AGEMA_reg_buffer_13710 ( .C (clk), .D (new_AGEMA_signal_34665), .Q (new_AGEMA_signal_34666) ) ;
    buf_clk new_AGEMA_reg_buffer_13714 ( .C (clk), .D (new_AGEMA_signal_34669), .Q (new_AGEMA_signal_34670) ) ;
    buf_clk new_AGEMA_reg_buffer_13718 ( .C (clk), .D (new_AGEMA_signal_34673), .Q (new_AGEMA_signal_34674) ) ;
    buf_clk new_AGEMA_reg_buffer_13722 ( .C (clk), .D (new_AGEMA_signal_34677), .Q (new_AGEMA_signal_34678) ) ;
    buf_clk new_AGEMA_reg_buffer_13726 ( .C (clk), .D (new_AGEMA_signal_34681), .Q (new_AGEMA_signal_34682) ) ;
    buf_clk new_AGEMA_reg_buffer_13730 ( .C (clk), .D (new_AGEMA_signal_34685), .Q (new_AGEMA_signal_34686) ) ;
    buf_clk new_AGEMA_reg_buffer_13734 ( .C (clk), .D (new_AGEMA_signal_34689), .Q (new_AGEMA_signal_34690) ) ;
    buf_clk new_AGEMA_reg_buffer_13738 ( .C (clk), .D (new_AGEMA_signal_34693), .Q (new_AGEMA_signal_34694) ) ;
    buf_clk new_AGEMA_reg_buffer_13742 ( .C (clk), .D (new_AGEMA_signal_34697), .Q (new_AGEMA_signal_34698) ) ;
    buf_clk new_AGEMA_reg_buffer_13746 ( .C (clk), .D (new_AGEMA_signal_34701), .Q (new_AGEMA_signal_34702) ) ;
    buf_clk new_AGEMA_reg_buffer_13750 ( .C (clk), .D (new_AGEMA_signal_34705), .Q (new_AGEMA_signal_34706) ) ;
    buf_clk new_AGEMA_reg_buffer_13754 ( .C (clk), .D (new_AGEMA_signal_34709), .Q (new_AGEMA_signal_34710) ) ;
    buf_clk new_AGEMA_reg_buffer_13758 ( .C (clk), .D (new_AGEMA_signal_34713), .Q (new_AGEMA_signal_34714) ) ;
    buf_clk new_AGEMA_reg_buffer_13762 ( .C (clk), .D (new_AGEMA_signal_34717), .Q (new_AGEMA_signal_34718) ) ;
    buf_clk new_AGEMA_reg_buffer_13766 ( .C (clk), .D (new_AGEMA_signal_34721), .Q (new_AGEMA_signal_34722) ) ;
    buf_clk new_AGEMA_reg_buffer_13770 ( .C (clk), .D (new_AGEMA_signal_34725), .Q (new_AGEMA_signal_34726) ) ;
    buf_clk new_AGEMA_reg_buffer_13774 ( .C (clk), .D (new_AGEMA_signal_34729), .Q (new_AGEMA_signal_34730) ) ;
    buf_clk new_AGEMA_reg_buffer_13778 ( .C (clk), .D (new_AGEMA_signal_34733), .Q (new_AGEMA_signal_34734) ) ;
    buf_clk new_AGEMA_reg_buffer_13782 ( .C (clk), .D (new_AGEMA_signal_34737), .Q (new_AGEMA_signal_34738) ) ;
    buf_clk new_AGEMA_reg_buffer_13786 ( .C (clk), .D (new_AGEMA_signal_34741), .Q (new_AGEMA_signal_34742) ) ;
    buf_clk new_AGEMA_reg_buffer_13790 ( .C (clk), .D (new_AGEMA_signal_34745), .Q (new_AGEMA_signal_34746) ) ;
    buf_clk new_AGEMA_reg_buffer_13794 ( .C (clk), .D (new_AGEMA_signal_34749), .Q (new_AGEMA_signal_34750) ) ;
    buf_clk new_AGEMA_reg_buffer_13798 ( .C (clk), .D (new_AGEMA_signal_34753), .Q (new_AGEMA_signal_34754) ) ;
    buf_clk new_AGEMA_reg_buffer_13802 ( .C (clk), .D (new_AGEMA_signal_34757), .Q (new_AGEMA_signal_34758) ) ;
    buf_clk new_AGEMA_reg_buffer_13806 ( .C (clk), .D (new_AGEMA_signal_34761), .Q (new_AGEMA_signal_34762) ) ;
    buf_clk new_AGEMA_reg_buffer_13810 ( .C (clk), .D (new_AGEMA_signal_34765), .Q (new_AGEMA_signal_34766) ) ;
    buf_clk new_AGEMA_reg_buffer_13814 ( .C (clk), .D (new_AGEMA_signal_34769), .Q (new_AGEMA_signal_34770) ) ;
    buf_clk new_AGEMA_reg_buffer_13818 ( .C (clk), .D (new_AGEMA_signal_34773), .Q (new_AGEMA_signal_34774) ) ;
    buf_clk new_AGEMA_reg_buffer_13822 ( .C (clk), .D (new_AGEMA_signal_34777), .Q (new_AGEMA_signal_34778) ) ;
    buf_clk new_AGEMA_reg_buffer_13826 ( .C (clk), .D (new_AGEMA_signal_34781), .Q (new_AGEMA_signal_34782) ) ;
    buf_clk new_AGEMA_reg_buffer_13830 ( .C (clk), .D (new_AGEMA_signal_34785), .Q (new_AGEMA_signal_34786) ) ;
    buf_clk new_AGEMA_reg_buffer_13834 ( .C (clk), .D (new_AGEMA_signal_34789), .Q (new_AGEMA_signal_34790) ) ;
    buf_clk new_AGEMA_reg_buffer_13838 ( .C (clk), .D (new_AGEMA_signal_34793), .Q (new_AGEMA_signal_34794) ) ;
    buf_clk new_AGEMA_reg_buffer_13842 ( .C (clk), .D (new_AGEMA_signal_34797), .Q (new_AGEMA_signal_34798) ) ;
    buf_clk new_AGEMA_reg_buffer_13846 ( .C (clk), .D (new_AGEMA_signal_34801), .Q (new_AGEMA_signal_34802) ) ;
    buf_clk new_AGEMA_reg_buffer_13850 ( .C (clk), .D (new_AGEMA_signal_34805), .Q (new_AGEMA_signal_34806) ) ;
    buf_clk new_AGEMA_reg_buffer_13854 ( .C (clk), .D (new_AGEMA_signal_34809), .Q (new_AGEMA_signal_34810) ) ;
    buf_clk new_AGEMA_reg_buffer_13858 ( .C (clk), .D (new_AGEMA_signal_34813), .Q (new_AGEMA_signal_34814) ) ;
    buf_clk new_AGEMA_reg_buffer_13862 ( .C (clk), .D (new_AGEMA_signal_34817), .Q (new_AGEMA_signal_34818) ) ;
    buf_clk new_AGEMA_reg_buffer_13866 ( .C (clk), .D (new_AGEMA_signal_34821), .Q (new_AGEMA_signal_34822) ) ;
    buf_clk new_AGEMA_reg_buffer_13870 ( .C (clk), .D (new_AGEMA_signal_34825), .Q (new_AGEMA_signal_34826) ) ;
    buf_clk new_AGEMA_reg_buffer_13874 ( .C (clk), .D (new_AGEMA_signal_34829), .Q (new_AGEMA_signal_34830) ) ;
    buf_clk new_AGEMA_reg_buffer_13878 ( .C (clk), .D (new_AGEMA_signal_34833), .Q (new_AGEMA_signal_34834) ) ;
    buf_clk new_AGEMA_reg_buffer_13882 ( .C (clk), .D (new_AGEMA_signal_34837), .Q (new_AGEMA_signal_34838) ) ;
    buf_clk new_AGEMA_reg_buffer_13886 ( .C (clk), .D (new_AGEMA_signal_34841), .Q (new_AGEMA_signal_34842) ) ;
    buf_clk new_AGEMA_reg_buffer_13890 ( .C (clk), .D (new_AGEMA_signal_34845), .Q (new_AGEMA_signal_34846) ) ;
    buf_clk new_AGEMA_reg_buffer_13894 ( .C (clk), .D (new_AGEMA_signal_34849), .Q (new_AGEMA_signal_34850) ) ;
    buf_clk new_AGEMA_reg_buffer_13898 ( .C (clk), .D (new_AGEMA_signal_34853), .Q (new_AGEMA_signal_34854) ) ;
    buf_clk new_AGEMA_reg_buffer_13902 ( .C (clk), .D (new_AGEMA_signal_34857), .Q (new_AGEMA_signal_34858) ) ;
    buf_clk new_AGEMA_reg_buffer_13906 ( .C (clk), .D (new_AGEMA_signal_34861), .Q (new_AGEMA_signal_34862) ) ;
    buf_clk new_AGEMA_reg_buffer_13910 ( .C (clk), .D (new_AGEMA_signal_34865), .Q (new_AGEMA_signal_34866) ) ;
    buf_clk new_AGEMA_reg_buffer_13914 ( .C (clk), .D (new_AGEMA_signal_34869), .Q (new_AGEMA_signal_34870) ) ;
    buf_clk new_AGEMA_reg_buffer_13918 ( .C (clk), .D (new_AGEMA_signal_34873), .Q (new_AGEMA_signal_34874) ) ;
    buf_clk new_AGEMA_reg_buffer_13922 ( .C (clk), .D (new_AGEMA_signal_34877), .Q (new_AGEMA_signal_34878) ) ;
    buf_clk new_AGEMA_reg_buffer_13926 ( .C (clk), .D (new_AGEMA_signal_34881), .Q (new_AGEMA_signal_34882) ) ;
    buf_clk new_AGEMA_reg_buffer_13930 ( .C (clk), .D (new_AGEMA_signal_34885), .Q (new_AGEMA_signal_34886) ) ;
    buf_clk new_AGEMA_reg_buffer_13934 ( .C (clk), .D (new_AGEMA_signal_34889), .Q (new_AGEMA_signal_34890) ) ;
    buf_clk new_AGEMA_reg_buffer_13938 ( .C (clk), .D (new_AGEMA_signal_34893), .Q (new_AGEMA_signal_34894) ) ;
    buf_clk new_AGEMA_reg_buffer_13942 ( .C (clk), .D (new_AGEMA_signal_34897), .Q (new_AGEMA_signal_34898) ) ;
    buf_clk new_AGEMA_reg_buffer_13946 ( .C (clk), .D (new_AGEMA_signal_34901), .Q (new_AGEMA_signal_34902) ) ;
    buf_clk new_AGEMA_reg_buffer_13950 ( .C (clk), .D (new_AGEMA_signal_34905), .Q (new_AGEMA_signal_34906) ) ;
    buf_clk new_AGEMA_reg_buffer_13954 ( .C (clk), .D (new_AGEMA_signal_34909), .Q (new_AGEMA_signal_34910) ) ;
    buf_clk new_AGEMA_reg_buffer_13958 ( .C (clk), .D (new_AGEMA_signal_34913), .Q (new_AGEMA_signal_34914) ) ;
    buf_clk new_AGEMA_reg_buffer_13962 ( .C (clk), .D (new_AGEMA_signal_34917), .Q (new_AGEMA_signal_34918) ) ;
    buf_clk new_AGEMA_reg_buffer_13966 ( .C (clk), .D (new_AGEMA_signal_34921), .Q (new_AGEMA_signal_34922) ) ;
    buf_clk new_AGEMA_reg_buffer_13970 ( .C (clk), .D (new_AGEMA_signal_34925), .Q (new_AGEMA_signal_34926) ) ;
    buf_clk new_AGEMA_reg_buffer_13974 ( .C (clk), .D (new_AGEMA_signal_34929), .Q (new_AGEMA_signal_34930) ) ;
    buf_clk new_AGEMA_reg_buffer_13978 ( .C (clk), .D (new_AGEMA_signal_34933), .Q (new_AGEMA_signal_34934) ) ;
    buf_clk new_AGEMA_reg_buffer_13982 ( .C (clk), .D (new_AGEMA_signal_34937), .Q (new_AGEMA_signal_34938) ) ;
    buf_clk new_AGEMA_reg_buffer_13986 ( .C (clk), .D (new_AGEMA_signal_34941), .Q (new_AGEMA_signal_34942) ) ;
    buf_clk new_AGEMA_reg_buffer_13990 ( .C (clk), .D (new_AGEMA_signal_34945), .Q (new_AGEMA_signal_34946) ) ;
    buf_clk new_AGEMA_reg_buffer_13994 ( .C (clk), .D (new_AGEMA_signal_34949), .Q (new_AGEMA_signal_34950) ) ;
    buf_clk new_AGEMA_reg_buffer_13998 ( .C (clk), .D (new_AGEMA_signal_34953), .Q (new_AGEMA_signal_34954) ) ;
    buf_clk new_AGEMA_reg_buffer_14002 ( .C (clk), .D (new_AGEMA_signal_34957), .Q (new_AGEMA_signal_34958) ) ;
    buf_clk new_AGEMA_reg_buffer_14006 ( .C (clk), .D (new_AGEMA_signal_34961), .Q (new_AGEMA_signal_34962) ) ;
    buf_clk new_AGEMA_reg_buffer_14010 ( .C (clk), .D (new_AGEMA_signal_34965), .Q (new_AGEMA_signal_34966) ) ;
    buf_clk new_AGEMA_reg_buffer_14014 ( .C (clk), .D (new_AGEMA_signal_34969), .Q (new_AGEMA_signal_34970) ) ;
    buf_clk new_AGEMA_reg_buffer_14018 ( .C (clk), .D (new_AGEMA_signal_34973), .Q (new_AGEMA_signal_34974) ) ;
    buf_clk new_AGEMA_reg_buffer_14022 ( .C (clk), .D (new_AGEMA_signal_34977), .Q (new_AGEMA_signal_34978) ) ;
    buf_clk new_AGEMA_reg_buffer_14026 ( .C (clk), .D (new_AGEMA_signal_34981), .Q (new_AGEMA_signal_34982) ) ;
    buf_clk new_AGEMA_reg_buffer_14030 ( .C (clk), .D (new_AGEMA_signal_34985), .Q (new_AGEMA_signal_34986) ) ;
    buf_clk new_AGEMA_reg_buffer_14034 ( .C (clk), .D (new_AGEMA_signal_34989), .Q (new_AGEMA_signal_34990) ) ;
    buf_clk new_AGEMA_reg_buffer_14038 ( .C (clk), .D (new_AGEMA_signal_34993), .Q (new_AGEMA_signal_34994) ) ;
    buf_clk new_AGEMA_reg_buffer_14042 ( .C (clk), .D (new_AGEMA_signal_34997), .Q (new_AGEMA_signal_34998) ) ;
    buf_clk new_AGEMA_reg_buffer_14046 ( .C (clk), .D (new_AGEMA_signal_35001), .Q (new_AGEMA_signal_35002) ) ;
    buf_clk new_AGEMA_reg_buffer_14050 ( .C (clk), .D (new_AGEMA_signal_35005), .Q (new_AGEMA_signal_35006) ) ;
    buf_clk new_AGEMA_reg_buffer_14054 ( .C (clk), .D (new_AGEMA_signal_35009), .Q (new_AGEMA_signal_35010) ) ;
    buf_clk new_AGEMA_reg_buffer_14058 ( .C (clk), .D (new_AGEMA_signal_35013), .Q (new_AGEMA_signal_35014) ) ;
    buf_clk new_AGEMA_reg_buffer_14062 ( .C (clk), .D (new_AGEMA_signal_35017), .Q (new_AGEMA_signal_35018) ) ;
    buf_clk new_AGEMA_reg_buffer_14066 ( .C (clk), .D (new_AGEMA_signal_35021), .Q (new_AGEMA_signal_35022) ) ;
    buf_clk new_AGEMA_reg_buffer_14070 ( .C (clk), .D (new_AGEMA_signal_35025), .Q (new_AGEMA_signal_35026) ) ;
    buf_clk new_AGEMA_reg_buffer_14074 ( .C (clk), .D (new_AGEMA_signal_35029), .Q (new_AGEMA_signal_35030) ) ;
    buf_clk new_AGEMA_reg_buffer_14078 ( .C (clk), .D (new_AGEMA_signal_35033), .Q (new_AGEMA_signal_35034) ) ;
    buf_clk new_AGEMA_reg_buffer_14082 ( .C (clk), .D (new_AGEMA_signal_35037), .Q (new_AGEMA_signal_35038) ) ;
    buf_clk new_AGEMA_reg_buffer_14086 ( .C (clk), .D (new_AGEMA_signal_35041), .Q (new_AGEMA_signal_35042) ) ;
    buf_clk new_AGEMA_reg_buffer_14090 ( .C (clk), .D (new_AGEMA_signal_35045), .Q (new_AGEMA_signal_35046) ) ;
    buf_clk new_AGEMA_reg_buffer_14094 ( .C (clk), .D (new_AGEMA_signal_35049), .Q (new_AGEMA_signal_35050) ) ;
    buf_clk new_AGEMA_reg_buffer_14098 ( .C (clk), .D (new_AGEMA_signal_35053), .Q (new_AGEMA_signal_35054) ) ;
    buf_clk new_AGEMA_reg_buffer_14102 ( .C (clk), .D (new_AGEMA_signal_35057), .Q (new_AGEMA_signal_35058) ) ;
    buf_clk new_AGEMA_reg_buffer_14106 ( .C (clk), .D (new_AGEMA_signal_35061), .Q (new_AGEMA_signal_35062) ) ;
    buf_clk new_AGEMA_reg_buffer_14110 ( .C (clk), .D (new_AGEMA_signal_35065), .Q (new_AGEMA_signal_35066) ) ;
    buf_clk new_AGEMA_reg_buffer_14114 ( .C (clk), .D (new_AGEMA_signal_35069), .Q (new_AGEMA_signal_35070) ) ;
    buf_clk new_AGEMA_reg_buffer_14118 ( .C (clk), .D (new_AGEMA_signal_35073), .Q (new_AGEMA_signal_35074) ) ;
    buf_clk new_AGEMA_reg_buffer_14122 ( .C (clk), .D (new_AGEMA_signal_35077), .Q (new_AGEMA_signal_35078) ) ;
    buf_clk new_AGEMA_reg_buffer_14126 ( .C (clk), .D (new_AGEMA_signal_35081), .Q (new_AGEMA_signal_35082) ) ;
    buf_clk new_AGEMA_reg_buffer_14130 ( .C (clk), .D (new_AGEMA_signal_35085), .Q (new_AGEMA_signal_35086) ) ;
    buf_clk new_AGEMA_reg_buffer_14134 ( .C (clk), .D (new_AGEMA_signal_35089), .Q (new_AGEMA_signal_35090) ) ;
    buf_clk new_AGEMA_reg_buffer_14138 ( .C (clk), .D (new_AGEMA_signal_35093), .Q (new_AGEMA_signal_35094) ) ;
    buf_clk new_AGEMA_reg_buffer_14142 ( .C (clk), .D (new_AGEMA_signal_35097), .Q (new_AGEMA_signal_35098) ) ;
    buf_clk new_AGEMA_reg_buffer_14146 ( .C (clk), .D (new_AGEMA_signal_35101), .Q (new_AGEMA_signal_35102) ) ;
    buf_clk new_AGEMA_reg_buffer_14150 ( .C (clk), .D (new_AGEMA_signal_35105), .Q (new_AGEMA_signal_35106) ) ;
    buf_clk new_AGEMA_reg_buffer_14154 ( .C (clk), .D (new_AGEMA_signal_35109), .Q (new_AGEMA_signal_35110) ) ;
    buf_clk new_AGEMA_reg_buffer_14158 ( .C (clk), .D (new_AGEMA_signal_35113), .Q (new_AGEMA_signal_35114) ) ;
    buf_clk new_AGEMA_reg_buffer_14162 ( .C (clk), .D (new_AGEMA_signal_35117), .Q (new_AGEMA_signal_35118) ) ;
    buf_clk new_AGEMA_reg_buffer_14166 ( .C (clk), .D (new_AGEMA_signal_35121), .Q (new_AGEMA_signal_35122) ) ;
    buf_clk new_AGEMA_reg_buffer_14170 ( .C (clk), .D (new_AGEMA_signal_35125), .Q (new_AGEMA_signal_35126) ) ;
    buf_clk new_AGEMA_reg_buffer_14174 ( .C (clk), .D (new_AGEMA_signal_35129), .Q (new_AGEMA_signal_35130) ) ;
    buf_clk new_AGEMA_reg_buffer_14178 ( .C (clk), .D (new_AGEMA_signal_35133), .Q (new_AGEMA_signal_35134) ) ;
    buf_clk new_AGEMA_reg_buffer_14182 ( .C (clk), .D (new_AGEMA_signal_35137), .Q (new_AGEMA_signal_35138) ) ;
    buf_clk new_AGEMA_reg_buffer_14186 ( .C (clk), .D (new_AGEMA_signal_35141), .Q (new_AGEMA_signal_35142) ) ;
    buf_clk new_AGEMA_reg_buffer_14190 ( .C (clk), .D (new_AGEMA_signal_35145), .Q (new_AGEMA_signal_35146) ) ;
    buf_clk new_AGEMA_reg_buffer_14194 ( .C (clk), .D (new_AGEMA_signal_35149), .Q (new_AGEMA_signal_35150) ) ;
    buf_clk new_AGEMA_reg_buffer_14198 ( .C (clk), .D (new_AGEMA_signal_35153), .Q (new_AGEMA_signal_35154) ) ;
    buf_clk new_AGEMA_reg_buffer_14202 ( .C (clk), .D (new_AGEMA_signal_35157), .Q (new_AGEMA_signal_35158) ) ;
    buf_clk new_AGEMA_reg_buffer_14206 ( .C (clk), .D (new_AGEMA_signal_35161), .Q (new_AGEMA_signal_35162) ) ;
    buf_clk new_AGEMA_reg_buffer_14210 ( .C (clk), .D (new_AGEMA_signal_35165), .Q (new_AGEMA_signal_35166) ) ;
    buf_clk new_AGEMA_reg_buffer_14214 ( .C (clk), .D (new_AGEMA_signal_35169), .Q (new_AGEMA_signal_35170) ) ;
    buf_clk new_AGEMA_reg_buffer_14218 ( .C (clk), .D (new_AGEMA_signal_35173), .Q (new_AGEMA_signal_35174) ) ;
    buf_clk new_AGEMA_reg_buffer_14222 ( .C (clk), .D (new_AGEMA_signal_35177), .Q (new_AGEMA_signal_35178) ) ;
    buf_clk new_AGEMA_reg_buffer_14226 ( .C (clk), .D (new_AGEMA_signal_35181), .Q (new_AGEMA_signal_35182) ) ;
    buf_clk new_AGEMA_reg_buffer_14230 ( .C (clk), .D (new_AGEMA_signal_35185), .Q (new_AGEMA_signal_35186) ) ;
    buf_clk new_AGEMA_reg_buffer_14234 ( .C (clk), .D (new_AGEMA_signal_35189), .Q (new_AGEMA_signal_35190) ) ;
    buf_clk new_AGEMA_reg_buffer_14238 ( .C (clk), .D (new_AGEMA_signal_35193), .Q (new_AGEMA_signal_35194) ) ;
    buf_clk new_AGEMA_reg_buffer_14242 ( .C (clk), .D (new_AGEMA_signal_35197), .Q (new_AGEMA_signal_35198) ) ;
    buf_clk new_AGEMA_reg_buffer_14246 ( .C (clk), .D (new_AGEMA_signal_35201), .Q (new_AGEMA_signal_35202) ) ;
    buf_clk new_AGEMA_reg_buffer_14250 ( .C (clk), .D (new_AGEMA_signal_35205), .Q (new_AGEMA_signal_35206) ) ;
    buf_clk new_AGEMA_reg_buffer_14254 ( .C (clk), .D (new_AGEMA_signal_35209), .Q (new_AGEMA_signal_35210) ) ;
    buf_clk new_AGEMA_reg_buffer_14258 ( .C (clk), .D (new_AGEMA_signal_35213), .Q (new_AGEMA_signal_35214) ) ;
    buf_clk new_AGEMA_reg_buffer_14262 ( .C (clk), .D (new_AGEMA_signal_35217), .Q (new_AGEMA_signal_35218) ) ;
    buf_clk new_AGEMA_reg_buffer_14266 ( .C (clk), .D (new_AGEMA_signal_35221), .Q (new_AGEMA_signal_35222) ) ;
    buf_clk new_AGEMA_reg_buffer_14270 ( .C (clk), .D (new_AGEMA_signal_35225), .Q (new_AGEMA_signal_35226) ) ;
    buf_clk new_AGEMA_reg_buffer_14274 ( .C (clk), .D (new_AGEMA_signal_35229), .Q (new_AGEMA_signal_35230) ) ;
    buf_clk new_AGEMA_reg_buffer_14278 ( .C (clk), .D (new_AGEMA_signal_35233), .Q (new_AGEMA_signal_35234) ) ;
    buf_clk new_AGEMA_reg_buffer_14282 ( .C (clk), .D (new_AGEMA_signal_35237), .Q (new_AGEMA_signal_35238) ) ;
    buf_clk new_AGEMA_reg_buffer_14286 ( .C (clk), .D (new_AGEMA_signal_35241), .Q (new_AGEMA_signal_35242) ) ;
    buf_clk new_AGEMA_reg_buffer_14290 ( .C (clk), .D (new_AGEMA_signal_35245), .Q (new_AGEMA_signal_35246) ) ;
    buf_clk new_AGEMA_reg_buffer_14294 ( .C (clk), .D (new_AGEMA_signal_35249), .Q (new_AGEMA_signal_35250) ) ;
    buf_clk new_AGEMA_reg_buffer_14298 ( .C (clk), .D (new_AGEMA_signal_35253), .Q (new_AGEMA_signal_35254) ) ;
    buf_clk new_AGEMA_reg_buffer_14302 ( .C (clk), .D (new_AGEMA_signal_35257), .Q (new_AGEMA_signal_35258) ) ;
    buf_clk new_AGEMA_reg_buffer_14306 ( .C (clk), .D (new_AGEMA_signal_35261), .Q (new_AGEMA_signal_35262) ) ;
    buf_clk new_AGEMA_reg_buffer_14310 ( .C (clk), .D (new_AGEMA_signal_35265), .Q (new_AGEMA_signal_35266) ) ;
    buf_clk new_AGEMA_reg_buffer_14314 ( .C (clk), .D (new_AGEMA_signal_35269), .Q (new_AGEMA_signal_35270) ) ;
    buf_clk new_AGEMA_reg_buffer_14318 ( .C (clk), .D (new_AGEMA_signal_35273), .Q (new_AGEMA_signal_35274) ) ;
    buf_clk new_AGEMA_reg_buffer_14322 ( .C (clk), .D (new_AGEMA_signal_35277), .Q (new_AGEMA_signal_35278) ) ;
    buf_clk new_AGEMA_reg_buffer_14326 ( .C (clk), .D (new_AGEMA_signal_35281), .Q (new_AGEMA_signal_35282) ) ;
    buf_clk new_AGEMA_reg_buffer_14330 ( .C (clk), .D (new_AGEMA_signal_35285), .Q (new_AGEMA_signal_35286) ) ;
    buf_clk new_AGEMA_reg_buffer_14334 ( .C (clk), .D (new_AGEMA_signal_35289), .Q (new_AGEMA_signal_35290) ) ;
    buf_clk new_AGEMA_reg_buffer_14338 ( .C (clk), .D (new_AGEMA_signal_35293), .Q (new_AGEMA_signal_35294) ) ;
    buf_clk new_AGEMA_reg_buffer_14342 ( .C (clk), .D (new_AGEMA_signal_35297), .Q (new_AGEMA_signal_35298) ) ;
    buf_clk new_AGEMA_reg_buffer_14346 ( .C (clk), .D (new_AGEMA_signal_35301), .Q (new_AGEMA_signal_35302) ) ;
    buf_clk new_AGEMA_reg_buffer_14350 ( .C (clk), .D (new_AGEMA_signal_35305), .Q (new_AGEMA_signal_35306) ) ;
    buf_clk new_AGEMA_reg_buffer_14354 ( .C (clk), .D (new_AGEMA_signal_35309), .Q (new_AGEMA_signal_35310) ) ;
    buf_clk new_AGEMA_reg_buffer_14358 ( .C (clk), .D (new_AGEMA_signal_35313), .Q (new_AGEMA_signal_35314) ) ;
    buf_clk new_AGEMA_reg_buffer_14362 ( .C (clk), .D (new_AGEMA_signal_35317), .Q (new_AGEMA_signal_35318) ) ;
    buf_clk new_AGEMA_reg_buffer_14366 ( .C (clk), .D (new_AGEMA_signal_35321), .Q (new_AGEMA_signal_35322) ) ;
    buf_clk new_AGEMA_reg_buffer_14370 ( .C (clk), .D (new_AGEMA_signal_35325), .Q (new_AGEMA_signal_35326) ) ;
    buf_clk new_AGEMA_reg_buffer_14374 ( .C (clk), .D (new_AGEMA_signal_35329), .Q (new_AGEMA_signal_35330) ) ;
    buf_clk new_AGEMA_reg_buffer_14378 ( .C (clk), .D (new_AGEMA_signal_35333), .Q (new_AGEMA_signal_35334) ) ;
    buf_clk new_AGEMA_reg_buffer_14382 ( .C (clk), .D (new_AGEMA_signal_35337), .Q (new_AGEMA_signal_35338) ) ;
    buf_clk new_AGEMA_reg_buffer_14386 ( .C (clk), .D (new_AGEMA_signal_35341), .Q (new_AGEMA_signal_35342) ) ;
    buf_clk new_AGEMA_reg_buffer_14390 ( .C (clk), .D (new_AGEMA_signal_35345), .Q (new_AGEMA_signal_35346) ) ;
    buf_clk new_AGEMA_reg_buffer_14394 ( .C (clk), .D (new_AGEMA_signal_35349), .Q (new_AGEMA_signal_35350) ) ;
    buf_clk new_AGEMA_reg_buffer_14398 ( .C (clk), .D (new_AGEMA_signal_35353), .Q (new_AGEMA_signal_35354) ) ;
    buf_clk new_AGEMA_reg_buffer_14402 ( .C (clk), .D (new_AGEMA_signal_35357), .Q (new_AGEMA_signal_35358) ) ;
    buf_clk new_AGEMA_reg_buffer_14406 ( .C (clk), .D (new_AGEMA_signal_35361), .Q (new_AGEMA_signal_35362) ) ;
    buf_clk new_AGEMA_reg_buffer_14410 ( .C (clk), .D (new_AGEMA_signal_35365), .Q (new_AGEMA_signal_35366) ) ;
    buf_clk new_AGEMA_reg_buffer_14414 ( .C (clk), .D (new_AGEMA_signal_35369), .Q (new_AGEMA_signal_35370) ) ;
    buf_clk new_AGEMA_reg_buffer_14418 ( .C (clk), .D (new_AGEMA_signal_35373), .Q (new_AGEMA_signal_35374) ) ;
    buf_clk new_AGEMA_reg_buffer_14422 ( .C (clk), .D (new_AGEMA_signal_35377), .Q (new_AGEMA_signal_35378) ) ;
    buf_clk new_AGEMA_reg_buffer_14426 ( .C (clk), .D (new_AGEMA_signal_35381), .Q (new_AGEMA_signal_35382) ) ;
    buf_clk new_AGEMA_reg_buffer_14430 ( .C (clk), .D (new_AGEMA_signal_35385), .Q (new_AGEMA_signal_35386) ) ;
    buf_clk new_AGEMA_reg_buffer_14434 ( .C (clk), .D (new_AGEMA_signal_35389), .Q (new_AGEMA_signal_35390) ) ;
    buf_clk new_AGEMA_reg_buffer_14438 ( .C (clk), .D (new_AGEMA_signal_35393), .Q (new_AGEMA_signal_35394) ) ;
    buf_clk new_AGEMA_reg_buffer_14442 ( .C (clk), .D (new_AGEMA_signal_35397), .Q (new_AGEMA_signal_35398) ) ;
    buf_clk new_AGEMA_reg_buffer_14446 ( .C (clk), .D (new_AGEMA_signal_35401), .Q (new_AGEMA_signal_35402) ) ;
    buf_clk new_AGEMA_reg_buffer_14450 ( .C (clk), .D (new_AGEMA_signal_35405), .Q (new_AGEMA_signal_35406) ) ;
    buf_clk new_AGEMA_reg_buffer_14454 ( .C (clk), .D (new_AGEMA_signal_35409), .Q (new_AGEMA_signal_35410) ) ;
    buf_clk new_AGEMA_reg_buffer_14458 ( .C (clk), .D (new_AGEMA_signal_35413), .Q (new_AGEMA_signal_35414) ) ;
    buf_clk new_AGEMA_reg_buffer_14462 ( .C (clk), .D (new_AGEMA_signal_35417), .Q (new_AGEMA_signal_35418) ) ;
    buf_clk new_AGEMA_reg_buffer_14466 ( .C (clk), .D (new_AGEMA_signal_35421), .Q (new_AGEMA_signal_35422) ) ;
    buf_clk new_AGEMA_reg_buffer_14470 ( .C (clk), .D (new_AGEMA_signal_35425), .Q (new_AGEMA_signal_35426) ) ;
    buf_clk new_AGEMA_reg_buffer_14474 ( .C (clk), .D (new_AGEMA_signal_35429), .Q (new_AGEMA_signal_35430) ) ;
    buf_clk new_AGEMA_reg_buffer_14478 ( .C (clk), .D (new_AGEMA_signal_35433), .Q (new_AGEMA_signal_35434) ) ;
    buf_clk new_AGEMA_reg_buffer_14482 ( .C (clk), .D (new_AGEMA_signal_35437), .Q (new_AGEMA_signal_35438) ) ;
    buf_clk new_AGEMA_reg_buffer_14486 ( .C (clk), .D (new_AGEMA_signal_35441), .Q (new_AGEMA_signal_35442) ) ;
    buf_clk new_AGEMA_reg_buffer_14490 ( .C (clk), .D (new_AGEMA_signal_35445), .Q (new_AGEMA_signal_35446) ) ;
    buf_clk new_AGEMA_reg_buffer_14494 ( .C (clk), .D (new_AGEMA_signal_35449), .Q (new_AGEMA_signal_35450) ) ;
    buf_clk new_AGEMA_reg_buffer_14498 ( .C (clk), .D (new_AGEMA_signal_35453), .Q (new_AGEMA_signal_35454) ) ;
    buf_clk new_AGEMA_reg_buffer_14502 ( .C (clk), .D (new_AGEMA_signal_35457), .Q (new_AGEMA_signal_35458) ) ;
    buf_clk new_AGEMA_reg_buffer_14506 ( .C (clk), .D (new_AGEMA_signal_35461), .Q (new_AGEMA_signal_35462) ) ;
    buf_clk new_AGEMA_reg_buffer_14510 ( .C (clk), .D (new_AGEMA_signal_35465), .Q (new_AGEMA_signal_35466) ) ;
    buf_clk new_AGEMA_reg_buffer_14514 ( .C (clk), .D (new_AGEMA_signal_35469), .Q (new_AGEMA_signal_35470) ) ;
    buf_clk new_AGEMA_reg_buffer_14518 ( .C (clk), .D (new_AGEMA_signal_35473), .Q (new_AGEMA_signal_35474) ) ;
    buf_clk new_AGEMA_reg_buffer_14522 ( .C (clk), .D (new_AGEMA_signal_35477), .Q (new_AGEMA_signal_35478) ) ;
    buf_clk new_AGEMA_reg_buffer_14526 ( .C (clk), .D (new_AGEMA_signal_35481), .Q (new_AGEMA_signal_35482) ) ;
    buf_clk new_AGEMA_reg_buffer_14530 ( .C (clk), .D (new_AGEMA_signal_35485), .Q (new_AGEMA_signal_35486) ) ;
    buf_clk new_AGEMA_reg_buffer_14534 ( .C (clk), .D (new_AGEMA_signal_35489), .Q (new_AGEMA_signal_35490) ) ;
    buf_clk new_AGEMA_reg_buffer_14538 ( .C (clk), .D (new_AGEMA_signal_35493), .Q (new_AGEMA_signal_35494) ) ;
    buf_clk new_AGEMA_reg_buffer_14542 ( .C (clk), .D (new_AGEMA_signal_35497), .Q (new_AGEMA_signal_35498) ) ;
    buf_clk new_AGEMA_reg_buffer_14546 ( .C (clk), .D (new_AGEMA_signal_35501), .Q (new_AGEMA_signal_35502) ) ;
    buf_clk new_AGEMA_reg_buffer_14550 ( .C (clk), .D (new_AGEMA_signal_35505), .Q (new_AGEMA_signal_35506) ) ;
    buf_clk new_AGEMA_reg_buffer_14554 ( .C (clk), .D (new_AGEMA_signal_35509), .Q (new_AGEMA_signal_35510) ) ;
    buf_clk new_AGEMA_reg_buffer_14558 ( .C (clk), .D (new_AGEMA_signal_35513), .Q (new_AGEMA_signal_35514) ) ;
    buf_clk new_AGEMA_reg_buffer_14562 ( .C (clk), .D (new_AGEMA_signal_35517), .Q (new_AGEMA_signal_35518) ) ;
    buf_clk new_AGEMA_reg_buffer_14566 ( .C (clk), .D (new_AGEMA_signal_35521), .Q (new_AGEMA_signal_35522) ) ;
    buf_clk new_AGEMA_reg_buffer_14570 ( .C (clk), .D (new_AGEMA_signal_35525), .Q (new_AGEMA_signal_35526) ) ;
    buf_clk new_AGEMA_reg_buffer_14574 ( .C (clk), .D (new_AGEMA_signal_35529), .Q (new_AGEMA_signal_35530) ) ;
    buf_clk new_AGEMA_reg_buffer_14578 ( .C (clk), .D (new_AGEMA_signal_35533), .Q (new_AGEMA_signal_35534) ) ;
    buf_clk new_AGEMA_reg_buffer_14582 ( .C (clk), .D (new_AGEMA_signal_35537), .Q (new_AGEMA_signal_35538) ) ;
    buf_clk new_AGEMA_reg_buffer_14586 ( .C (clk), .D (new_AGEMA_signal_35541), .Q (new_AGEMA_signal_35542) ) ;
    buf_clk new_AGEMA_reg_buffer_14590 ( .C (clk), .D (new_AGEMA_signal_35545), .Q (new_AGEMA_signal_35546) ) ;
    buf_clk new_AGEMA_reg_buffer_14594 ( .C (clk), .D (new_AGEMA_signal_35549), .Q (new_AGEMA_signal_35550) ) ;
    buf_clk new_AGEMA_reg_buffer_14598 ( .C (clk), .D (new_AGEMA_signal_35553), .Q (new_AGEMA_signal_35554) ) ;
    buf_clk new_AGEMA_reg_buffer_14602 ( .C (clk), .D (new_AGEMA_signal_35557), .Q (new_AGEMA_signal_35558) ) ;
    buf_clk new_AGEMA_reg_buffer_14606 ( .C (clk), .D (new_AGEMA_signal_35561), .Q (new_AGEMA_signal_35562) ) ;
    buf_clk new_AGEMA_reg_buffer_14610 ( .C (clk), .D (new_AGEMA_signal_35565), .Q (new_AGEMA_signal_35566) ) ;
    buf_clk new_AGEMA_reg_buffer_14614 ( .C (clk), .D (new_AGEMA_signal_35569), .Q (new_AGEMA_signal_35570) ) ;
    buf_clk new_AGEMA_reg_buffer_14618 ( .C (clk), .D (new_AGEMA_signal_35573), .Q (new_AGEMA_signal_35574) ) ;
    buf_clk new_AGEMA_reg_buffer_14622 ( .C (clk), .D (new_AGEMA_signal_35577), .Q (new_AGEMA_signal_35578) ) ;
    buf_clk new_AGEMA_reg_buffer_14626 ( .C (clk), .D (new_AGEMA_signal_35581), .Q (new_AGEMA_signal_35582) ) ;
    buf_clk new_AGEMA_reg_buffer_14630 ( .C (clk), .D (new_AGEMA_signal_35585), .Q (new_AGEMA_signal_35586) ) ;
    buf_clk new_AGEMA_reg_buffer_14634 ( .C (clk), .D (new_AGEMA_signal_35589), .Q (new_AGEMA_signal_35590) ) ;
    buf_clk new_AGEMA_reg_buffer_14638 ( .C (clk), .D (new_AGEMA_signal_35593), .Q (new_AGEMA_signal_35594) ) ;
    buf_clk new_AGEMA_reg_buffer_14642 ( .C (clk), .D (new_AGEMA_signal_35597), .Q (new_AGEMA_signal_35598) ) ;
    buf_clk new_AGEMA_reg_buffer_14646 ( .C (clk), .D (new_AGEMA_signal_35601), .Q (new_AGEMA_signal_35602) ) ;
    buf_clk new_AGEMA_reg_buffer_14650 ( .C (clk), .D (new_AGEMA_signal_35605), .Q (new_AGEMA_signal_35606) ) ;
    buf_clk new_AGEMA_reg_buffer_14654 ( .C (clk), .D (new_AGEMA_signal_35609), .Q (new_AGEMA_signal_35610) ) ;
    buf_clk new_AGEMA_reg_buffer_14658 ( .C (clk), .D (new_AGEMA_signal_35613), .Q (new_AGEMA_signal_35614) ) ;
    buf_clk new_AGEMA_reg_buffer_14662 ( .C (clk), .D (new_AGEMA_signal_35617), .Q (new_AGEMA_signal_35618) ) ;
    buf_clk new_AGEMA_reg_buffer_14666 ( .C (clk), .D (new_AGEMA_signal_35621), .Q (new_AGEMA_signal_35622) ) ;
    buf_clk new_AGEMA_reg_buffer_14670 ( .C (clk), .D (new_AGEMA_signal_35625), .Q (new_AGEMA_signal_35626) ) ;
    buf_clk new_AGEMA_reg_buffer_14674 ( .C (clk), .D (new_AGEMA_signal_35629), .Q (new_AGEMA_signal_35630) ) ;
    buf_clk new_AGEMA_reg_buffer_14678 ( .C (clk), .D (new_AGEMA_signal_35633), .Q (new_AGEMA_signal_35634) ) ;
    buf_clk new_AGEMA_reg_buffer_14682 ( .C (clk), .D (new_AGEMA_signal_35637), .Q (new_AGEMA_signal_35638) ) ;
    buf_clk new_AGEMA_reg_buffer_14686 ( .C (clk), .D (new_AGEMA_signal_35641), .Q (new_AGEMA_signal_35642) ) ;
    buf_clk new_AGEMA_reg_buffer_14690 ( .C (clk), .D (new_AGEMA_signal_35645), .Q (new_AGEMA_signal_35646) ) ;
    buf_clk new_AGEMA_reg_buffer_14694 ( .C (clk), .D (new_AGEMA_signal_35649), .Q (new_AGEMA_signal_35650) ) ;
    buf_clk new_AGEMA_reg_buffer_14698 ( .C (clk), .D (new_AGEMA_signal_35653), .Q (new_AGEMA_signal_35654) ) ;
    buf_clk new_AGEMA_reg_buffer_14702 ( .C (clk), .D (new_AGEMA_signal_35657), .Q (new_AGEMA_signal_35658) ) ;
    buf_clk new_AGEMA_reg_buffer_14706 ( .C (clk), .D (new_AGEMA_signal_35661), .Q (new_AGEMA_signal_35662) ) ;
    buf_clk new_AGEMA_reg_buffer_14710 ( .C (clk), .D (new_AGEMA_signal_35665), .Q (new_AGEMA_signal_35666) ) ;
    buf_clk new_AGEMA_reg_buffer_14714 ( .C (clk), .D (new_AGEMA_signal_35669), .Q (new_AGEMA_signal_35670) ) ;
    buf_clk new_AGEMA_reg_buffer_14718 ( .C (clk), .D (new_AGEMA_signal_35673), .Q (new_AGEMA_signal_35674) ) ;
    buf_clk new_AGEMA_reg_buffer_14722 ( .C (clk), .D (new_AGEMA_signal_35677), .Q (new_AGEMA_signal_35678) ) ;
    buf_clk new_AGEMA_reg_buffer_14726 ( .C (clk), .D (new_AGEMA_signal_35681), .Q (new_AGEMA_signal_35682) ) ;
    buf_clk new_AGEMA_reg_buffer_14730 ( .C (clk), .D (new_AGEMA_signal_35685), .Q (new_AGEMA_signal_35686) ) ;
    buf_clk new_AGEMA_reg_buffer_14734 ( .C (clk), .D (new_AGEMA_signal_35689), .Q (new_AGEMA_signal_35690) ) ;
    buf_clk new_AGEMA_reg_buffer_14738 ( .C (clk), .D (new_AGEMA_signal_35693), .Q (new_AGEMA_signal_35694) ) ;
    buf_clk new_AGEMA_reg_buffer_14742 ( .C (clk), .D (new_AGEMA_signal_35697), .Q (new_AGEMA_signal_35698) ) ;
    buf_clk new_AGEMA_reg_buffer_14746 ( .C (clk), .D (new_AGEMA_signal_35701), .Q (new_AGEMA_signal_35702) ) ;
    buf_clk new_AGEMA_reg_buffer_14750 ( .C (clk), .D (new_AGEMA_signal_35705), .Q (new_AGEMA_signal_35706) ) ;
    buf_clk new_AGEMA_reg_buffer_14754 ( .C (clk), .D (new_AGEMA_signal_35709), .Q (new_AGEMA_signal_35710) ) ;
    buf_clk new_AGEMA_reg_buffer_14758 ( .C (clk), .D (new_AGEMA_signal_35713), .Q (new_AGEMA_signal_35714) ) ;
    buf_clk new_AGEMA_reg_buffer_14762 ( .C (clk), .D (new_AGEMA_signal_35717), .Q (new_AGEMA_signal_35718) ) ;
    buf_clk new_AGEMA_reg_buffer_14766 ( .C (clk), .D (new_AGEMA_signal_35721), .Q (new_AGEMA_signal_35722) ) ;
    buf_clk new_AGEMA_reg_buffer_14770 ( .C (clk), .D (new_AGEMA_signal_35725), .Q (new_AGEMA_signal_35726) ) ;
    buf_clk new_AGEMA_reg_buffer_14774 ( .C (clk), .D (new_AGEMA_signal_35729), .Q (new_AGEMA_signal_35730) ) ;
    buf_clk new_AGEMA_reg_buffer_14778 ( .C (clk), .D (new_AGEMA_signal_35733), .Q (new_AGEMA_signal_35734) ) ;
    buf_clk new_AGEMA_reg_buffer_14782 ( .C (clk), .D (new_AGEMA_signal_35737), .Q (new_AGEMA_signal_35738) ) ;
    buf_clk new_AGEMA_reg_buffer_14786 ( .C (clk), .D (new_AGEMA_signal_35741), .Q (new_AGEMA_signal_35742) ) ;
    buf_clk new_AGEMA_reg_buffer_14790 ( .C (clk), .D (new_AGEMA_signal_35745), .Q (new_AGEMA_signal_35746) ) ;
    buf_clk new_AGEMA_reg_buffer_14794 ( .C (clk), .D (new_AGEMA_signal_35749), .Q (new_AGEMA_signal_35750) ) ;
    buf_clk new_AGEMA_reg_buffer_14798 ( .C (clk), .D (new_AGEMA_signal_35753), .Q (new_AGEMA_signal_35754) ) ;
    buf_clk new_AGEMA_reg_buffer_14802 ( .C (clk), .D (new_AGEMA_signal_35757), .Q (new_AGEMA_signal_35758) ) ;
    buf_clk new_AGEMA_reg_buffer_14806 ( .C (clk), .D (new_AGEMA_signal_35761), .Q (new_AGEMA_signal_35762) ) ;
    buf_clk new_AGEMA_reg_buffer_14810 ( .C (clk), .D (new_AGEMA_signal_35765), .Q (new_AGEMA_signal_35766) ) ;
    buf_clk new_AGEMA_reg_buffer_14814 ( .C (clk), .D (new_AGEMA_signal_35769), .Q (new_AGEMA_signal_35770) ) ;
    buf_clk new_AGEMA_reg_buffer_14818 ( .C (clk), .D (new_AGEMA_signal_35773), .Q (new_AGEMA_signal_35774) ) ;
    buf_clk new_AGEMA_reg_buffer_14822 ( .C (clk), .D (new_AGEMA_signal_35777), .Q (new_AGEMA_signal_35778) ) ;
    buf_clk new_AGEMA_reg_buffer_14826 ( .C (clk), .D (new_AGEMA_signal_35781), .Q (new_AGEMA_signal_35782) ) ;
    buf_clk new_AGEMA_reg_buffer_14830 ( .C (clk), .D (new_AGEMA_signal_35785), .Q (new_AGEMA_signal_35786) ) ;
    buf_clk new_AGEMA_reg_buffer_14834 ( .C (clk), .D (new_AGEMA_signal_35789), .Q (new_AGEMA_signal_35790) ) ;
    buf_clk new_AGEMA_reg_buffer_14837 ( .C (clk), .D (new_AGEMA_signal_35792), .Q (new_AGEMA_signal_35793) ) ;
    buf_clk new_AGEMA_reg_buffer_14840 ( .C (clk), .D (new_AGEMA_signal_35795), .Q (new_AGEMA_signal_35796) ) ;
    buf_clk new_AGEMA_reg_buffer_14843 ( .C (clk), .D (new_AGEMA_signal_35798), .Q (new_AGEMA_signal_35799) ) ;
    buf_clk new_AGEMA_reg_buffer_14846 ( .C (clk), .D (new_AGEMA_signal_35801), .Q (new_AGEMA_signal_35802) ) ;
    buf_clk new_AGEMA_reg_buffer_14849 ( .C (clk), .D (new_AGEMA_signal_35804), .Q (new_AGEMA_signal_35805) ) ;
    buf_clk new_AGEMA_reg_buffer_14852 ( .C (clk), .D (new_AGEMA_signal_35807), .Q (new_AGEMA_signal_35808) ) ;
    buf_clk new_AGEMA_reg_buffer_14855 ( .C (clk), .D (new_AGEMA_signal_35810), .Q (new_AGEMA_signal_35811) ) ;
    buf_clk new_AGEMA_reg_buffer_14858 ( .C (clk), .D (new_AGEMA_signal_35813), .Q (new_AGEMA_signal_35814) ) ;
    buf_clk new_AGEMA_reg_buffer_14861 ( .C (clk), .D (new_AGEMA_signal_35816), .Q (new_AGEMA_signal_35817) ) ;
    buf_clk new_AGEMA_reg_buffer_14864 ( .C (clk), .D (new_AGEMA_signal_35819), .Q (new_AGEMA_signal_35820) ) ;
    buf_clk new_AGEMA_reg_buffer_14867 ( .C (clk), .D (new_AGEMA_signal_35822), .Q (new_AGEMA_signal_35823) ) ;
    buf_clk new_AGEMA_reg_buffer_14870 ( .C (clk), .D (new_AGEMA_signal_35825), .Q (new_AGEMA_signal_35826) ) ;
    buf_clk new_AGEMA_reg_buffer_14873 ( .C (clk), .D (new_AGEMA_signal_35828), .Q (new_AGEMA_signal_35829) ) ;
    buf_clk new_AGEMA_reg_buffer_14876 ( .C (clk), .D (new_AGEMA_signal_35831), .Q (new_AGEMA_signal_35832) ) ;
    buf_clk new_AGEMA_reg_buffer_14879 ( .C (clk), .D (new_AGEMA_signal_35834), .Q (new_AGEMA_signal_35835) ) ;
    buf_clk new_AGEMA_reg_buffer_14882 ( .C (clk), .D (new_AGEMA_signal_35837), .Q (new_AGEMA_signal_35838) ) ;
    buf_clk new_AGEMA_reg_buffer_14885 ( .C (clk), .D (new_AGEMA_signal_35840), .Q (new_AGEMA_signal_35841) ) ;
    buf_clk new_AGEMA_reg_buffer_14888 ( .C (clk), .D (new_AGEMA_signal_35843), .Q (new_AGEMA_signal_35844) ) ;
    buf_clk new_AGEMA_reg_buffer_14891 ( .C (clk), .D (new_AGEMA_signal_35846), .Q (new_AGEMA_signal_35847) ) ;
    buf_clk new_AGEMA_reg_buffer_14894 ( .C (clk), .D (new_AGEMA_signal_35849), .Q (new_AGEMA_signal_35850) ) ;
    buf_clk new_AGEMA_reg_buffer_14897 ( .C (clk), .D (new_AGEMA_signal_35852), .Q (new_AGEMA_signal_35853) ) ;
    buf_clk new_AGEMA_reg_buffer_14900 ( .C (clk), .D (new_AGEMA_signal_35855), .Q (new_AGEMA_signal_35856) ) ;
    buf_clk new_AGEMA_reg_buffer_14903 ( .C (clk), .D (new_AGEMA_signal_35858), .Q (new_AGEMA_signal_35859) ) ;
    buf_clk new_AGEMA_reg_buffer_14906 ( .C (clk), .D (new_AGEMA_signal_35861), .Q (new_AGEMA_signal_35862) ) ;
    buf_clk new_AGEMA_reg_buffer_14909 ( .C (clk), .D (new_AGEMA_signal_35864), .Q (new_AGEMA_signal_35865) ) ;
    buf_clk new_AGEMA_reg_buffer_14912 ( .C (clk), .D (new_AGEMA_signal_35867), .Q (new_AGEMA_signal_35868) ) ;
    buf_clk new_AGEMA_reg_buffer_14915 ( .C (clk), .D (new_AGEMA_signal_35870), .Q (new_AGEMA_signal_35871) ) ;
    buf_clk new_AGEMA_reg_buffer_14918 ( .C (clk), .D (new_AGEMA_signal_35873), .Q (new_AGEMA_signal_35874) ) ;
    buf_clk new_AGEMA_reg_buffer_14921 ( .C (clk), .D (new_AGEMA_signal_35876), .Q (new_AGEMA_signal_35877) ) ;
    buf_clk new_AGEMA_reg_buffer_14924 ( .C (clk), .D (new_AGEMA_signal_35879), .Q (new_AGEMA_signal_35880) ) ;
    buf_clk new_AGEMA_reg_buffer_14927 ( .C (clk), .D (new_AGEMA_signal_35882), .Q (new_AGEMA_signal_35883) ) ;
    buf_clk new_AGEMA_reg_buffer_14930 ( .C (clk), .D (new_AGEMA_signal_35885), .Q (new_AGEMA_signal_35886) ) ;
    buf_clk new_AGEMA_reg_buffer_14933 ( .C (clk), .D (new_AGEMA_signal_35888), .Q (new_AGEMA_signal_35889) ) ;
    buf_clk new_AGEMA_reg_buffer_14936 ( .C (clk), .D (new_AGEMA_signal_35891), .Q (new_AGEMA_signal_35892) ) ;
    buf_clk new_AGEMA_reg_buffer_14939 ( .C (clk), .D (new_AGEMA_signal_35894), .Q (new_AGEMA_signal_35895) ) ;
    buf_clk new_AGEMA_reg_buffer_14942 ( .C (clk), .D (new_AGEMA_signal_35897), .Q (new_AGEMA_signal_35898) ) ;
    buf_clk new_AGEMA_reg_buffer_14945 ( .C (clk), .D (new_AGEMA_signal_35900), .Q (new_AGEMA_signal_35901) ) ;
    buf_clk new_AGEMA_reg_buffer_14948 ( .C (clk), .D (new_AGEMA_signal_35903), .Q (new_AGEMA_signal_35904) ) ;
    buf_clk new_AGEMA_reg_buffer_14951 ( .C (clk), .D (new_AGEMA_signal_35906), .Q (new_AGEMA_signal_35907) ) ;
    buf_clk new_AGEMA_reg_buffer_14954 ( .C (clk), .D (new_AGEMA_signal_35909), .Q (new_AGEMA_signal_35910) ) ;
    buf_clk new_AGEMA_reg_buffer_14957 ( .C (clk), .D (new_AGEMA_signal_35912), .Q (new_AGEMA_signal_35913) ) ;
    buf_clk new_AGEMA_reg_buffer_14960 ( .C (clk), .D (new_AGEMA_signal_35915), .Q (new_AGEMA_signal_35916) ) ;
    buf_clk new_AGEMA_reg_buffer_14963 ( .C (clk), .D (new_AGEMA_signal_35918), .Q (new_AGEMA_signal_35919) ) ;
    buf_clk new_AGEMA_reg_buffer_14966 ( .C (clk), .D (new_AGEMA_signal_35921), .Q (new_AGEMA_signal_35922) ) ;
    buf_clk new_AGEMA_reg_buffer_14969 ( .C (clk), .D (new_AGEMA_signal_35924), .Q (new_AGEMA_signal_35925) ) ;
    buf_clk new_AGEMA_reg_buffer_14972 ( .C (clk), .D (new_AGEMA_signal_35927), .Q (new_AGEMA_signal_35928) ) ;
    buf_clk new_AGEMA_reg_buffer_14975 ( .C (clk), .D (new_AGEMA_signal_35930), .Q (new_AGEMA_signal_35931) ) ;
    buf_clk new_AGEMA_reg_buffer_14978 ( .C (clk), .D (new_AGEMA_signal_35933), .Q (new_AGEMA_signal_35934) ) ;
    buf_clk new_AGEMA_reg_buffer_14981 ( .C (clk), .D (new_AGEMA_signal_35936), .Q (new_AGEMA_signal_35937) ) ;
    buf_clk new_AGEMA_reg_buffer_14984 ( .C (clk), .D (new_AGEMA_signal_35939), .Q (new_AGEMA_signal_35940) ) ;
    buf_clk new_AGEMA_reg_buffer_14987 ( .C (clk), .D (new_AGEMA_signal_35942), .Q (new_AGEMA_signal_35943) ) ;
    buf_clk new_AGEMA_reg_buffer_14990 ( .C (clk), .D (new_AGEMA_signal_35945), .Q (new_AGEMA_signal_35946) ) ;
    buf_clk new_AGEMA_reg_buffer_14993 ( .C (clk), .D (new_AGEMA_signal_35948), .Q (new_AGEMA_signal_35949) ) ;
    buf_clk new_AGEMA_reg_buffer_14996 ( .C (clk), .D (new_AGEMA_signal_35951), .Q (new_AGEMA_signal_35952) ) ;
    buf_clk new_AGEMA_reg_buffer_14999 ( .C (clk), .D (new_AGEMA_signal_35954), .Q (new_AGEMA_signal_35955) ) ;
    buf_clk new_AGEMA_reg_buffer_15002 ( .C (clk), .D (new_AGEMA_signal_35957), .Q (new_AGEMA_signal_35958) ) ;
    buf_clk new_AGEMA_reg_buffer_15005 ( .C (clk), .D (new_AGEMA_signal_35960), .Q (new_AGEMA_signal_35961) ) ;
    buf_clk new_AGEMA_reg_buffer_15008 ( .C (clk), .D (new_AGEMA_signal_35963), .Q (new_AGEMA_signal_35964) ) ;
    buf_clk new_AGEMA_reg_buffer_15011 ( .C (clk), .D (new_AGEMA_signal_35966), .Q (new_AGEMA_signal_35967) ) ;
    buf_clk new_AGEMA_reg_buffer_15014 ( .C (clk), .D (new_AGEMA_signal_35969), .Q (new_AGEMA_signal_35970) ) ;
    buf_clk new_AGEMA_reg_buffer_15017 ( .C (clk), .D (new_AGEMA_signal_35972), .Q (new_AGEMA_signal_35973) ) ;
    buf_clk new_AGEMA_reg_buffer_15020 ( .C (clk), .D (new_AGEMA_signal_35975), .Q (new_AGEMA_signal_35976) ) ;
    buf_clk new_AGEMA_reg_buffer_15023 ( .C (clk), .D (new_AGEMA_signal_35978), .Q (new_AGEMA_signal_35979) ) ;
    buf_clk new_AGEMA_reg_buffer_15026 ( .C (clk), .D (new_AGEMA_signal_35981), .Q (new_AGEMA_signal_35982) ) ;
    buf_clk new_AGEMA_reg_buffer_15029 ( .C (clk), .D (new_AGEMA_signal_35984), .Q (new_AGEMA_signal_35985) ) ;
    buf_clk new_AGEMA_reg_buffer_15032 ( .C (clk), .D (new_AGEMA_signal_35987), .Q (new_AGEMA_signal_35988) ) ;
    buf_clk new_AGEMA_reg_buffer_15035 ( .C (clk), .D (new_AGEMA_signal_35990), .Q (new_AGEMA_signal_35991) ) ;
    buf_clk new_AGEMA_reg_buffer_15038 ( .C (clk), .D (new_AGEMA_signal_35993), .Q (new_AGEMA_signal_35994) ) ;
    buf_clk new_AGEMA_reg_buffer_15041 ( .C (clk), .D (new_AGEMA_signal_35996), .Q (new_AGEMA_signal_35997) ) ;
    buf_clk new_AGEMA_reg_buffer_15044 ( .C (clk), .D (new_AGEMA_signal_35999), .Q (new_AGEMA_signal_36000) ) ;
    buf_clk new_AGEMA_reg_buffer_15047 ( .C (clk), .D (new_AGEMA_signal_36002), .Q (new_AGEMA_signal_36003) ) ;
    buf_clk new_AGEMA_reg_buffer_15050 ( .C (clk), .D (new_AGEMA_signal_36005), .Q (new_AGEMA_signal_36006) ) ;
    buf_clk new_AGEMA_reg_buffer_15053 ( .C (clk), .D (new_AGEMA_signal_36008), .Q (new_AGEMA_signal_36009) ) ;
    buf_clk new_AGEMA_reg_buffer_15056 ( .C (clk), .D (new_AGEMA_signal_36011), .Q (new_AGEMA_signal_36012) ) ;
    buf_clk new_AGEMA_reg_buffer_15059 ( .C (clk), .D (new_AGEMA_signal_36014), .Q (new_AGEMA_signal_36015) ) ;
    buf_clk new_AGEMA_reg_buffer_15062 ( .C (clk), .D (new_AGEMA_signal_36017), .Q (new_AGEMA_signal_36018) ) ;
    buf_clk new_AGEMA_reg_buffer_15065 ( .C (clk), .D (new_AGEMA_signal_36020), .Q (new_AGEMA_signal_36021) ) ;
    buf_clk new_AGEMA_reg_buffer_15068 ( .C (clk), .D (new_AGEMA_signal_36023), .Q (new_AGEMA_signal_36024) ) ;
    buf_clk new_AGEMA_reg_buffer_15071 ( .C (clk), .D (new_AGEMA_signal_36026), .Q (new_AGEMA_signal_36027) ) ;
    buf_clk new_AGEMA_reg_buffer_15074 ( .C (clk), .D (new_AGEMA_signal_36029), .Q (new_AGEMA_signal_36030) ) ;
    buf_clk new_AGEMA_reg_buffer_15077 ( .C (clk), .D (new_AGEMA_signal_36032), .Q (new_AGEMA_signal_36033) ) ;
    buf_clk new_AGEMA_reg_buffer_15080 ( .C (clk), .D (new_AGEMA_signal_36035), .Q (new_AGEMA_signal_36036) ) ;
    buf_clk new_AGEMA_reg_buffer_15083 ( .C (clk), .D (new_AGEMA_signal_36038), .Q (new_AGEMA_signal_36039) ) ;
    buf_clk new_AGEMA_reg_buffer_15086 ( .C (clk), .D (new_AGEMA_signal_36041), .Q (new_AGEMA_signal_36042) ) ;
    buf_clk new_AGEMA_reg_buffer_15089 ( .C (clk), .D (new_AGEMA_signal_36044), .Q (new_AGEMA_signal_36045) ) ;
    buf_clk new_AGEMA_reg_buffer_15092 ( .C (clk), .D (new_AGEMA_signal_36047), .Q (new_AGEMA_signal_36048) ) ;
    buf_clk new_AGEMA_reg_buffer_15095 ( .C (clk), .D (new_AGEMA_signal_36050), .Q (new_AGEMA_signal_36051) ) ;
    buf_clk new_AGEMA_reg_buffer_15098 ( .C (clk), .D (new_AGEMA_signal_36053), .Q (new_AGEMA_signal_36054) ) ;
    buf_clk new_AGEMA_reg_buffer_15101 ( .C (clk), .D (new_AGEMA_signal_36056), .Q (new_AGEMA_signal_36057) ) ;
    buf_clk new_AGEMA_reg_buffer_15104 ( .C (clk), .D (new_AGEMA_signal_36059), .Q (new_AGEMA_signal_36060) ) ;
    buf_clk new_AGEMA_reg_buffer_15107 ( .C (clk), .D (new_AGEMA_signal_36062), .Q (new_AGEMA_signal_36063) ) ;
    buf_clk new_AGEMA_reg_buffer_15110 ( .C (clk), .D (new_AGEMA_signal_36065), .Q (new_AGEMA_signal_36066) ) ;
    buf_clk new_AGEMA_reg_buffer_15113 ( .C (clk), .D (new_AGEMA_signal_36068), .Q (new_AGEMA_signal_36069) ) ;
    buf_clk new_AGEMA_reg_buffer_15116 ( .C (clk), .D (new_AGEMA_signal_36071), .Q (new_AGEMA_signal_36072) ) ;
    buf_clk new_AGEMA_reg_buffer_15119 ( .C (clk), .D (new_AGEMA_signal_36074), .Q (new_AGEMA_signal_36075) ) ;
    buf_clk new_AGEMA_reg_buffer_15122 ( .C (clk), .D (new_AGEMA_signal_36077), .Q (new_AGEMA_signal_36078) ) ;
    buf_clk new_AGEMA_reg_buffer_15125 ( .C (clk), .D (new_AGEMA_signal_36080), .Q (new_AGEMA_signal_36081) ) ;
    buf_clk new_AGEMA_reg_buffer_15128 ( .C (clk), .D (new_AGEMA_signal_36083), .Q (new_AGEMA_signal_36084) ) ;
    buf_clk new_AGEMA_reg_buffer_15131 ( .C (clk), .D (new_AGEMA_signal_36086), .Q (new_AGEMA_signal_36087) ) ;
    buf_clk new_AGEMA_reg_buffer_15134 ( .C (clk), .D (new_AGEMA_signal_36089), .Q (new_AGEMA_signal_36090) ) ;
    buf_clk new_AGEMA_reg_buffer_15137 ( .C (clk), .D (new_AGEMA_signal_36092), .Q (new_AGEMA_signal_36093) ) ;
    buf_clk new_AGEMA_reg_buffer_15140 ( .C (clk), .D (new_AGEMA_signal_36095), .Q (new_AGEMA_signal_36096) ) ;
    buf_clk new_AGEMA_reg_buffer_15143 ( .C (clk), .D (new_AGEMA_signal_36098), .Q (new_AGEMA_signal_36099) ) ;
    buf_clk new_AGEMA_reg_buffer_15146 ( .C (clk), .D (new_AGEMA_signal_36101), .Q (new_AGEMA_signal_36102) ) ;
    buf_clk new_AGEMA_reg_buffer_15149 ( .C (clk), .D (new_AGEMA_signal_36104), .Q (new_AGEMA_signal_36105) ) ;
    buf_clk new_AGEMA_reg_buffer_15152 ( .C (clk), .D (new_AGEMA_signal_36107), .Q (new_AGEMA_signal_36108) ) ;
    buf_clk new_AGEMA_reg_buffer_15155 ( .C (clk), .D (new_AGEMA_signal_36110), .Q (new_AGEMA_signal_36111) ) ;
    buf_clk new_AGEMA_reg_buffer_15158 ( .C (clk), .D (new_AGEMA_signal_36113), .Q (new_AGEMA_signal_36114) ) ;
    buf_clk new_AGEMA_reg_buffer_15161 ( .C (clk), .D (new_AGEMA_signal_36116), .Q (new_AGEMA_signal_36117) ) ;
    buf_clk new_AGEMA_reg_buffer_15164 ( .C (clk), .D (new_AGEMA_signal_36119), .Q (new_AGEMA_signal_36120) ) ;
    buf_clk new_AGEMA_reg_buffer_15167 ( .C (clk), .D (new_AGEMA_signal_36122), .Q (new_AGEMA_signal_36123) ) ;
    buf_clk new_AGEMA_reg_buffer_15170 ( .C (clk), .D (new_AGEMA_signal_36125), .Q (new_AGEMA_signal_36126) ) ;
    buf_clk new_AGEMA_reg_buffer_15173 ( .C (clk), .D (new_AGEMA_signal_36128), .Q (new_AGEMA_signal_36129) ) ;
    buf_clk new_AGEMA_reg_buffer_15176 ( .C (clk), .D (new_AGEMA_signal_36131), .Q (new_AGEMA_signal_36132) ) ;
    buf_clk new_AGEMA_reg_buffer_15179 ( .C (clk), .D (new_AGEMA_signal_36134), .Q (new_AGEMA_signal_36135) ) ;
    buf_clk new_AGEMA_reg_buffer_15182 ( .C (clk), .D (new_AGEMA_signal_36137), .Q (new_AGEMA_signal_36138) ) ;
    buf_clk new_AGEMA_reg_buffer_15185 ( .C (clk), .D (new_AGEMA_signal_36140), .Q (new_AGEMA_signal_36141) ) ;
    buf_clk new_AGEMA_reg_buffer_15188 ( .C (clk), .D (new_AGEMA_signal_36143), .Q (new_AGEMA_signal_36144) ) ;
    buf_clk new_AGEMA_reg_buffer_15191 ( .C (clk), .D (new_AGEMA_signal_36146), .Q (new_AGEMA_signal_36147) ) ;
    buf_clk new_AGEMA_reg_buffer_15194 ( .C (clk), .D (new_AGEMA_signal_36149), .Q (new_AGEMA_signal_36150) ) ;
    buf_clk new_AGEMA_reg_buffer_15197 ( .C (clk), .D (new_AGEMA_signal_36152), .Q (new_AGEMA_signal_36153) ) ;
    buf_clk new_AGEMA_reg_buffer_15200 ( .C (clk), .D (new_AGEMA_signal_36155), .Q (new_AGEMA_signal_36156) ) ;
    buf_clk new_AGEMA_reg_buffer_15203 ( .C (clk), .D (new_AGEMA_signal_36158), .Q (new_AGEMA_signal_36159) ) ;
    buf_clk new_AGEMA_reg_buffer_15206 ( .C (clk), .D (new_AGEMA_signal_36161), .Q (new_AGEMA_signal_36162) ) ;
    buf_clk new_AGEMA_reg_buffer_15209 ( .C (clk), .D (new_AGEMA_signal_36164), .Q (new_AGEMA_signal_36165) ) ;
    buf_clk new_AGEMA_reg_buffer_15212 ( .C (clk), .D (new_AGEMA_signal_36167), .Q (new_AGEMA_signal_36168) ) ;
    buf_clk new_AGEMA_reg_buffer_15215 ( .C (clk), .D (new_AGEMA_signal_36170), .Q (new_AGEMA_signal_36171) ) ;
    buf_clk new_AGEMA_reg_buffer_15218 ( .C (clk), .D (new_AGEMA_signal_36173), .Q (new_AGEMA_signal_36174) ) ;
    buf_clk new_AGEMA_reg_buffer_15221 ( .C (clk), .D (new_AGEMA_signal_36176), .Q (new_AGEMA_signal_36177) ) ;
    buf_clk new_AGEMA_reg_buffer_15224 ( .C (clk), .D (new_AGEMA_signal_36179), .Q (new_AGEMA_signal_36180) ) ;
    buf_clk new_AGEMA_reg_buffer_15227 ( .C (clk), .D (new_AGEMA_signal_36182), .Q (new_AGEMA_signal_36183) ) ;
    buf_clk new_AGEMA_reg_buffer_15230 ( .C (clk), .D (new_AGEMA_signal_36185), .Q (new_AGEMA_signal_36186) ) ;
    buf_clk new_AGEMA_reg_buffer_15233 ( .C (clk), .D (new_AGEMA_signal_36188), .Q (new_AGEMA_signal_36189) ) ;
    buf_clk new_AGEMA_reg_buffer_15236 ( .C (clk), .D (new_AGEMA_signal_36191), .Q (new_AGEMA_signal_36192) ) ;
    buf_clk new_AGEMA_reg_buffer_15239 ( .C (clk), .D (new_AGEMA_signal_36194), .Q (new_AGEMA_signal_36195) ) ;
    buf_clk new_AGEMA_reg_buffer_15242 ( .C (clk), .D (new_AGEMA_signal_36197), .Q (new_AGEMA_signal_36198) ) ;
    buf_clk new_AGEMA_reg_buffer_15245 ( .C (clk), .D (new_AGEMA_signal_36200), .Q (new_AGEMA_signal_36201) ) ;
    buf_clk new_AGEMA_reg_buffer_15248 ( .C (clk), .D (new_AGEMA_signal_36203), .Q (new_AGEMA_signal_36204) ) ;
    buf_clk new_AGEMA_reg_buffer_15251 ( .C (clk), .D (new_AGEMA_signal_36206), .Q (new_AGEMA_signal_36207) ) ;
    buf_clk new_AGEMA_reg_buffer_15254 ( .C (clk), .D (new_AGEMA_signal_36209), .Q (new_AGEMA_signal_36210) ) ;
    buf_clk new_AGEMA_reg_buffer_15257 ( .C (clk), .D (new_AGEMA_signal_36212), .Q (new_AGEMA_signal_36213) ) ;
    buf_clk new_AGEMA_reg_buffer_15260 ( .C (clk), .D (new_AGEMA_signal_36215), .Q (new_AGEMA_signal_36216) ) ;
    buf_clk new_AGEMA_reg_buffer_15263 ( .C (clk), .D (new_AGEMA_signal_36218), .Q (new_AGEMA_signal_36219) ) ;
    buf_clk new_AGEMA_reg_buffer_15266 ( .C (clk), .D (new_AGEMA_signal_36221), .Q (new_AGEMA_signal_36222) ) ;
    buf_clk new_AGEMA_reg_buffer_15269 ( .C (clk), .D (new_AGEMA_signal_36224), .Q (new_AGEMA_signal_36225) ) ;
    buf_clk new_AGEMA_reg_buffer_15272 ( .C (clk), .D (new_AGEMA_signal_36227), .Q (new_AGEMA_signal_36228) ) ;
    buf_clk new_AGEMA_reg_buffer_15275 ( .C (clk), .D (new_AGEMA_signal_36230), .Q (new_AGEMA_signal_36231) ) ;
    buf_clk new_AGEMA_reg_buffer_15278 ( .C (clk), .D (new_AGEMA_signal_36233), .Q (new_AGEMA_signal_36234) ) ;
    buf_clk new_AGEMA_reg_buffer_15281 ( .C (clk), .D (new_AGEMA_signal_36236), .Q (new_AGEMA_signal_36237) ) ;
    buf_clk new_AGEMA_reg_buffer_15284 ( .C (clk), .D (new_AGEMA_signal_36239), .Q (new_AGEMA_signal_36240) ) ;
    buf_clk new_AGEMA_reg_buffer_15287 ( .C (clk), .D (new_AGEMA_signal_36242), .Q (new_AGEMA_signal_36243) ) ;
    buf_clk new_AGEMA_reg_buffer_15290 ( .C (clk), .D (new_AGEMA_signal_36245), .Q (new_AGEMA_signal_36246) ) ;
    buf_clk new_AGEMA_reg_buffer_15293 ( .C (clk), .D (new_AGEMA_signal_36248), .Q (new_AGEMA_signal_36249) ) ;
    buf_clk new_AGEMA_reg_buffer_15296 ( .C (clk), .D (new_AGEMA_signal_36251), .Q (new_AGEMA_signal_36252) ) ;
    buf_clk new_AGEMA_reg_buffer_15299 ( .C (clk), .D (new_AGEMA_signal_36254), .Q (new_AGEMA_signal_36255) ) ;
    buf_clk new_AGEMA_reg_buffer_15302 ( .C (clk), .D (new_AGEMA_signal_36257), .Q (new_AGEMA_signal_36258) ) ;
    buf_clk new_AGEMA_reg_buffer_15305 ( .C (clk), .D (new_AGEMA_signal_36260), .Q (new_AGEMA_signal_36261) ) ;
    buf_clk new_AGEMA_reg_buffer_15308 ( .C (clk), .D (new_AGEMA_signal_36263), .Q (new_AGEMA_signal_36264) ) ;
    buf_clk new_AGEMA_reg_buffer_15311 ( .C (clk), .D (new_AGEMA_signal_36266), .Q (new_AGEMA_signal_36267) ) ;
    buf_clk new_AGEMA_reg_buffer_15314 ( .C (clk), .D (new_AGEMA_signal_36269), .Q (new_AGEMA_signal_36270) ) ;
    buf_clk new_AGEMA_reg_buffer_15317 ( .C (clk), .D (new_AGEMA_signal_36272), .Q (new_AGEMA_signal_36273) ) ;
    buf_clk new_AGEMA_reg_buffer_15320 ( .C (clk), .D (new_AGEMA_signal_36275), .Q (new_AGEMA_signal_36276) ) ;
    buf_clk new_AGEMA_reg_buffer_15323 ( .C (clk), .D (new_AGEMA_signal_36278), .Q (new_AGEMA_signal_36279) ) ;
    buf_clk new_AGEMA_reg_buffer_15326 ( .C (clk), .D (new_AGEMA_signal_36281), .Q (new_AGEMA_signal_36282) ) ;
    buf_clk new_AGEMA_reg_buffer_15329 ( .C (clk), .D (new_AGEMA_signal_36284), .Q (new_AGEMA_signal_36285) ) ;
    buf_clk new_AGEMA_reg_buffer_15332 ( .C (clk), .D (new_AGEMA_signal_36287), .Q (new_AGEMA_signal_36288) ) ;
    buf_clk new_AGEMA_reg_buffer_15335 ( .C (clk), .D (new_AGEMA_signal_36290), .Q (new_AGEMA_signal_36291) ) ;
    buf_clk new_AGEMA_reg_buffer_15338 ( .C (clk), .D (new_AGEMA_signal_36293), .Q (new_AGEMA_signal_36294) ) ;
    buf_clk new_AGEMA_reg_buffer_15341 ( .C (clk), .D (new_AGEMA_signal_36296), .Q (new_AGEMA_signal_36297) ) ;
    buf_clk new_AGEMA_reg_buffer_15344 ( .C (clk), .D (new_AGEMA_signal_36299), .Q (new_AGEMA_signal_36300) ) ;
    buf_clk new_AGEMA_reg_buffer_15347 ( .C (clk), .D (new_AGEMA_signal_36302), .Q (new_AGEMA_signal_36303) ) ;
    buf_clk new_AGEMA_reg_buffer_15350 ( .C (clk), .D (new_AGEMA_signal_36305), .Q (new_AGEMA_signal_36306) ) ;
    buf_clk new_AGEMA_reg_buffer_15353 ( .C (clk), .D (new_AGEMA_signal_36308), .Q (new_AGEMA_signal_36309) ) ;
    buf_clk new_AGEMA_reg_buffer_15356 ( .C (clk), .D (new_AGEMA_signal_36311), .Q (new_AGEMA_signal_36312) ) ;
    buf_clk new_AGEMA_reg_buffer_15359 ( .C (clk), .D (new_AGEMA_signal_36314), .Q (new_AGEMA_signal_36315) ) ;
    buf_clk new_AGEMA_reg_buffer_15362 ( .C (clk), .D (new_AGEMA_signal_36317), .Q (new_AGEMA_signal_36318) ) ;
    buf_clk new_AGEMA_reg_buffer_15365 ( .C (clk), .D (new_AGEMA_signal_36320), .Q (new_AGEMA_signal_36321) ) ;
    buf_clk new_AGEMA_reg_buffer_15368 ( .C (clk), .D (new_AGEMA_signal_36323), .Q (new_AGEMA_signal_36324) ) ;
    buf_clk new_AGEMA_reg_buffer_15371 ( .C (clk), .D (new_AGEMA_signal_36326), .Q (new_AGEMA_signal_36327) ) ;
    buf_clk new_AGEMA_reg_buffer_15374 ( .C (clk), .D (new_AGEMA_signal_36329), .Q (new_AGEMA_signal_36330) ) ;
    buf_clk new_AGEMA_reg_buffer_15377 ( .C (clk), .D (new_AGEMA_signal_36332), .Q (new_AGEMA_signal_36333) ) ;
    buf_clk new_AGEMA_reg_buffer_15380 ( .C (clk), .D (new_AGEMA_signal_36335), .Q (new_AGEMA_signal_36336) ) ;
    buf_clk new_AGEMA_reg_buffer_15383 ( .C (clk), .D (new_AGEMA_signal_36338), .Q (new_AGEMA_signal_36339) ) ;
    buf_clk new_AGEMA_reg_buffer_15386 ( .C (clk), .D (new_AGEMA_signal_36341), .Q (new_AGEMA_signal_36342) ) ;
    buf_clk new_AGEMA_reg_buffer_15389 ( .C (clk), .D (new_AGEMA_signal_36344), .Q (new_AGEMA_signal_36345) ) ;
    buf_clk new_AGEMA_reg_buffer_15392 ( .C (clk), .D (new_AGEMA_signal_36347), .Q (new_AGEMA_signal_36348) ) ;
    buf_clk new_AGEMA_reg_buffer_15395 ( .C (clk), .D (new_AGEMA_signal_36350), .Q (new_AGEMA_signal_36351) ) ;
    buf_clk new_AGEMA_reg_buffer_15398 ( .C (clk), .D (new_AGEMA_signal_36353), .Q (new_AGEMA_signal_36354) ) ;
    buf_clk new_AGEMA_reg_buffer_15401 ( .C (clk), .D (new_AGEMA_signal_36356), .Q (new_AGEMA_signal_36357) ) ;
    buf_clk new_AGEMA_reg_buffer_15404 ( .C (clk), .D (new_AGEMA_signal_36359), .Q (new_AGEMA_signal_36360) ) ;
    buf_clk new_AGEMA_reg_buffer_15407 ( .C (clk), .D (new_AGEMA_signal_36362), .Q (new_AGEMA_signal_36363) ) ;
    buf_clk new_AGEMA_reg_buffer_15410 ( .C (clk), .D (new_AGEMA_signal_36365), .Q (new_AGEMA_signal_36366) ) ;
    buf_clk new_AGEMA_reg_buffer_15413 ( .C (clk), .D (new_AGEMA_signal_36368), .Q (new_AGEMA_signal_36369) ) ;
    buf_clk new_AGEMA_reg_buffer_15416 ( .C (clk), .D (new_AGEMA_signal_36371), .Q (new_AGEMA_signal_36372) ) ;
    buf_clk new_AGEMA_reg_buffer_15419 ( .C (clk), .D (new_AGEMA_signal_36374), .Q (new_AGEMA_signal_36375) ) ;
    buf_clk new_AGEMA_reg_buffer_15422 ( .C (clk), .D (new_AGEMA_signal_36377), .Q (new_AGEMA_signal_36378) ) ;
    buf_clk new_AGEMA_reg_buffer_15425 ( .C (clk), .D (new_AGEMA_signal_36380), .Q (new_AGEMA_signal_36381) ) ;
    buf_clk new_AGEMA_reg_buffer_15428 ( .C (clk), .D (new_AGEMA_signal_36383), .Q (new_AGEMA_signal_36384) ) ;
    buf_clk new_AGEMA_reg_buffer_15431 ( .C (clk), .D (new_AGEMA_signal_36386), .Q (new_AGEMA_signal_36387) ) ;
    buf_clk new_AGEMA_reg_buffer_15434 ( .C (clk), .D (new_AGEMA_signal_36389), .Q (new_AGEMA_signal_36390) ) ;
    buf_clk new_AGEMA_reg_buffer_15437 ( .C (clk), .D (new_AGEMA_signal_36392), .Q (new_AGEMA_signal_36393) ) ;
    buf_clk new_AGEMA_reg_buffer_15440 ( .C (clk), .D (new_AGEMA_signal_36395), .Q (new_AGEMA_signal_36396) ) ;
    buf_clk new_AGEMA_reg_buffer_15443 ( .C (clk), .D (new_AGEMA_signal_36398), .Q (new_AGEMA_signal_36399) ) ;
    buf_clk new_AGEMA_reg_buffer_15446 ( .C (clk), .D (new_AGEMA_signal_36401), .Q (new_AGEMA_signal_36402) ) ;
    buf_clk new_AGEMA_reg_buffer_15449 ( .C (clk), .D (new_AGEMA_signal_36404), .Q (new_AGEMA_signal_36405) ) ;
    buf_clk new_AGEMA_reg_buffer_15452 ( .C (clk), .D (new_AGEMA_signal_36407), .Q (new_AGEMA_signal_36408) ) ;
    buf_clk new_AGEMA_reg_buffer_15455 ( .C (clk), .D (new_AGEMA_signal_36410), .Q (new_AGEMA_signal_36411) ) ;
    buf_clk new_AGEMA_reg_buffer_15458 ( .C (clk), .D (new_AGEMA_signal_36413), .Q (new_AGEMA_signal_36414) ) ;
    buf_clk new_AGEMA_reg_buffer_15461 ( .C (clk), .D (new_AGEMA_signal_36416), .Q (new_AGEMA_signal_36417) ) ;
    buf_clk new_AGEMA_reg_buffer_15464 ( .C (clk), .D (new_AGEMA_signal_36419), .Q (new_AGEMA_signal_36420) ) ;
    buf_clk new_AGEMA_reg_buffer_15467 ( .C (clk), .D (new_AGEMA_signal_36422), .Q (new_AGEMA_signal_36423) ) ;
    buf_clk new_AGEMA_reg_buffer_15470 ( .C (clk), .D (new_AGEMA_signal_36425), .Q (new_AGEMA_signal_36426) ) ;
    buf_clk new_AGEMA_reg_buffer_15473 ( .C (clk), .D (new_AGEMA_signal_36428), .Q (new_AGEMA_signal_36429) ) ;
    buf_clk new_AGEMA_reg_buffer_15476 ( .C (clk), .D (new_AGEMA_signal_36431), .Q (new_AGEMA_signal_36432) ) ;
    buf_clk new_AGEMA_reg_buffer_15479 ( .C (clk), .D (new_AGEMA_signal_36434), .Q (new_AGEMA_signal_36435) ) ;
    buf_clk new_AGEMA_reg_buffer_15482 ( .C (clk), .D (new_AGEMA_signal_36437), .Q (new_AGEMA_signal_36438) ) ;
    buf_clk new_AGEMA_reg_buffer_15485 ( .C (clk), .D (new_AGEMA_signal_36440), .Q (new_AGEMA_signal_36441) ) ;
    buf_clk new_AGEMA_reg_buffer_15488 ( .C (clk), .D (new_AGEMA_signal_36443), .Q (new_AGEMA_signal_36444) ) ;
    buf_clk new_AGEMA_reg_buffer_15491 ( .C (clk), .D (new_AGEMA_signal_36446), .Q (new_AGEMA_signal_36447) ) ;
    buf_clk new_AGEMA_reg_buffer_15494 ( .C (clk), .D (new_AGEMA_signal_36449), .Q (new_AGEMA_signal_36450) ) ;
    buf_clk new_AGEMA_reg_buffer_15497 ( .C (clk), .D (new_AGEMA_signal_36452), .Q (new_AGEMA_signal_36453) ) ;
    buf_clk new_AGEMA_reg_buffer_15500 ( .C (clk), .D (new_AGEMA_signal_36455), .Q (new_AGEMA_signal_36456) ) ;
    buf_clk new_AGEMA_reg_buffer_15503 ( .C (clk), .D (new_AGEMA_signal_36458), .Q (new_AGEMA_signal_36459) ) ;
    buf_clk new_AGEMA_reg_buffer_15506 ( .C (clk), .D (new_AGEMA_signal_36461), .Q (new_AGEMA_signal_36462) ) ;
    buf_clk new_AGEMA_reg_buffer_15509 ( .C (clk), .D (new_AGEMA_signal_36464), .Q (new_AGEMA_signal_36465) ) ;
    buf_clk new_AGEMA_reg_buffer_15512 ( .C (clk), .D (new_AGEMA_signal_36467), .Q (new_AGEMA_signal_36468) ) ;
    buf_clk new_AGEMA_reg_buffer_15515 ( .C (clk), .D (new_AGEMA_signal_36470), .Q (new_AGEMA_signal_36471) ) ;
    buf_clk new_AGEMA_reg_buffer_15518 ( .C (clk), .D (new_AGEMA_signal_36473), .Q (new_AGEMA_signal_36474) ) ;
    buf_clk new_AGEMA_reg_buffer_15521 ( .C (clk), .D (new_AGEMA_signal_36476), .Q (new_AGEMA_signal_36477) ) ;
    buf_clk new_AGEMA_reg_buffer_15524 ( .C (clk), .D (new_AGEMA_signal_36479), .Q (new_AGEMA_signal_36480) ) ;
    buf_clk new_AGEMA_reg_buffer_15527 ( .C (clk), .D (new_AGEMA_signal_36482), .Q (new_AGEMA_signal_36483) ) ;
    buf_clk new_AGEMA_reg_buffer_15530 ( .C (clk), .D (new_AGEMA_signal_36485), .Q (new_AGEMA_signal_36486) ) ;
    buf_clk new_AGEMA_reg_buffer_15533 ( .C (clk), .D (new_AGEMA_signal_36488), .Q (new_AGEMA_signal_36489) ) ;
    buf_clk new_AGEMA_reg_buffer_15536 ( .C (clk), .D (new_AGEMA_signal_36491), .Q (new_AGEMA_signal_36492) ) ;
    buf_clk new_AGEMA_reg_buffer_15539 ( .C (clk), .D (new_AGEMA_signal_36494), .Q (new_AGEMA_signal_36495) ) ;
    buf_clk new_AGEMA_reg_buffer_15542 ( .C (clk), .D (new_AGEMA_signal_36497), .Q (new_AGEMA_signal_36498) ) ;
    buf_clk new_AGEMA_reg_buffer_15545 ( .C (clk), .D (new_AGEMA_signal_36500), .Q (new_AGEMA_signal_36501) ) ;
    buf_clk new_AGEMA_reg_buffer_15548 ( .C (clk), .D (new_AGEMA_signal_36503), .Q (new_AGEMA_signal_36504) ) ;
    buf_clk new_AGEMA_reg_buffer_15551 ( .C (clk), .D (new_AGEMA_signal_36506), .Q (new_AGEMA_signal_36507) ) ;
    buf_clk new_AGEMA_reg_buffer_15554 ( .C (clk), .D (new_AGEMA_signal_36509), .Q (new_AGEMA_signal_36510) ) ;
    buf_clk new_AGEMA_reg_buffer_15557 ( .C (clk), .D (new_AGEMA_signal_36512), .Q (new_AGEMA_signal_36513) ) ;
    buf_clk new_AGEMA_reg_buffer_15560 ( .C (clk), .D (new_AGEMA_signal_36515), .Q (new_AGEMA_signal_36516) ) ;
    buf_clk new_AGEMA_reg_buffer_15563 ( .C (clk), .D (new_AGEMA_signal_36518), .Q (new_AGEMA_signal_36519) ) ;
    buf_clk new_AGEMA_reg_buffer_15566 ( .C (clk), .D (new_AGEMA_signal_36521), .Q (new_AGEMA_signal_36522) ) ;
    buf_clk new_AGEMA_reg_buffer_15569 ( .C (clk), .D (new_AGEMA_signal_36524), .Q (new_AGEMA_signal_36525) ) ;
    buf_clk new_AGEMA_reg_buffer_15572 ( .C (clk), .D (new_AGEMA_signal_36527), .Q (new_AGEMA_signal_36528) ) ;
    buf_clk new_AGEMA_reg_buffer_15575 ( .C (clk), .D (new_AGEMA_signal_36530), .Q (new_AGEMA_signal_36531) ) ;
    buf_clk new_AGEMA_reg_buffer_15578 ( .C (clk), .D (new_AGEMA_signal_36533), .Q (new_AGEMA_signal_36534) ) ;
    buf_clk new_AGEMA_reg_buffer_15581 ( .C (clk), .D (new_AGEMA_signal_36536), .Q (new_AGEMA_signal_36537) ) ;
    buf_clk new_AGEMA_reg_buffer_15584 ( .C (clk), .D (new_AGEMA_signal_36539), .Q (new_AGEMA_signal_36540) ) ;
    buf_clk new_AGEMA_reg_buffer_15587 ( .C (clk), .D (new_AGEMA_signal_36542), .Q (new_AGEMA_signal_36543) ) ;
    buf_clk new_AGEMA_reg_buffer_15590 ( .C (clk), .D (new_AGEMA_signal_36545), .Q (new_AGEMA_signal_36546) ) ;
    buf_clk new_AGEMA_reg_buffer_15593 ( .C (clk), .D (new_AGEMA_signal_36548), .Q (new_AGEMA_signal_36549) ) ;
    buf_clk new_AGEMA_reg_buffer_15596 ( .C (clk), .D (new_AGEMA_signal_36551), .Q (new_AGEMA_signal_36552) ) ;
    buf_clk new_AGEMA_reg_buffer_15599 ( .C (clk), .D (new_AGEMA_signal_36554), .Q (new_AGEMA_signal_36555) ) ;
    buf_clk new_AGEMA_reg_buffer_15602 ( .C (clk), .D (new_AGEMA_signal_36557), .Q (new_AGEMA_signal_36558) ) ;
    buf_clk new_AGEMA_reg_buffer_15605 ( .C (clk), .D (new_AGEMA_signal_36560), .Q (new_AGEMA_signal_36561) ) ;
    buf_clk new_AGEMA_reg_buffer_15608 ( .C (clk), .D (new_AGEMA_signal_36563), .Q (new_AGEMA_signal_36564) ) ;
    buf_clk new_AGEMA_reg_buffer_15611 ( .C (clk), .D (new_AGEMA_signal_36566), .Q (new_AGEMA_signal_36567) ) ;
    buf_clk new_AGEMA_reg_buffer_15614 ( .C (clk), .D (new_AGEMA_signal_36569), .Q (new_AGEMA_signal_36570) ) ;
    buf_clk new_AGEMA_reg_buffer_15617 ( .C (clk), .D (new_AGEMA_signal_36572), .Q (new_AGEMA_signal_36573) ) ;
    buf_clk new_AGEMA_reg_buffer_15620 ( .C (clk), .D (new_AGEMA_signal_36575), .Q (new_AGEMA_signal_36576) ) ;
    buf_clk new_AGEMA_reg_buffer_15623 ( .C (clk), .D (new_AGEMA_signal_36578), .Q (new_AGEMA_signal_36579) ) ;
    buf_clk new_AGEMA_reg_buffer_15626 ( .C (clk), .D (new_AGEMA_signal_36581), .Q (new_AGEMA_signal_36582) ) ;
    buf_clk new_AGEMA_reg_buffer_15629 ( .C (clk), .D (new_AGEMA_signal_36584), .Q (new_AGEMA_signal_36585) ) ;
    buf_clk new_AGEMA_reg_buffer_15632 ( .C (clk), .D (new_AGEMA_signal_36587), .Q (new_AGEMA_signal_36588) ) ;
    buf_clk new_AGEMA_reg_buffer_15635 ( .C (clk), .D (new_AGEMA_signal_36590), .Q (new_AGEMA_signal_36591) ) ;
    buf_clk new_AGEMA_reg_buffer_15638 ( .C (clk), .D (new_AGEMA_signal_36593), .Q (new_AGEMA_signal_36594) ) ;
    buf_clk new_AGEMA_reg_buffer_15641 ( .C (clk), .D (new_AGEMA_signal_36596), .Q (new_AGEMA_signal_36597) ) ;
    buf_clk new_AGEMA_reg_buffer_15644 ( .C (clk), .D (new_AGEMA_signal_36599), .Q (new_AGEMA_signal_36600) ) ;
    buf_clk new_AGEMA_reg_buffer_15647 ( .C (clk), .D (new_AGEMA_signal_36602), .Q (new_AGEMA_signal_36603) ) ;
    buf_clk new_AGEMA_reg_buffer_15650 ( .C (clk), .D (new_AGEMA_signal_36605), .Q (new_AGEMA_signal_36606) ) ;
    buf_clk new_AGEMA_reg_buffer_15654 ( .C (clk), .D (new_AGEMA_signal_36609), .Q (new_AGEMA_signal_36610) ) ;
    buf_clk new_AGEMA_reg_buffer_15658 ( .C (clk), .D (new_AGEMA_signal_36613), .Q (new_AGEMA_signal_36614) ) ;
    buf_clk new_AGEMA_reg_buffer_15662 ( .C (clk), .D (new_AGEMA_signal_36617), .Q (new_AGEMA_signal_36618) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_25496, new_AGEMA_signal_25495, new_AGEMA_signal_25494, new_AGEMA_signal_25493}), .clk (clk), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, new_AGEMA_signal_8944, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_25500, new_AGEMA_signal_25499, new_AGEMA_signal_25498, new_AGEMA_signal_25497}), .clk (clk), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, new_AGEMA_signal_9244, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_25496, new_AGEMA_signal_25495, new_AGEMA_signal_25494, new_AGEMA_signal_25493}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, new_AGEMA_signal_8950, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910], Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_25500, new_AGEMA_signal_25499, new_AGEMA_signal_25498, new_AGEMA_signal_25497}), .b ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, new_AGEMA_signal_8698, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, new_AGEMA_signal_9250, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_25808, new_AGEMA_signal_25807, new_AGEMA_signal_25806, new_AGEMA_signal_25805}), .b ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_25812, new_AGEMA_signal_25811, new_AGEMA_signal_25810, new_AGEMA_signal_25809}), .c ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_25816, new_AGEMA_signal_25815, new_AGEMA_signal_25814, new_AGEMA_signal_25813}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, new_AGEMA_signal_9244, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, new_AGEMA_signal_9250, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_25820, new_AGEMA_signal_25819, new_AGEMA_signal_25818, new_AGEMA_signal_25817}), .c ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, new_AGEMA_signal_8962, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_25512, new_AGEMA_signal_25511, new_AGEMA_signal_25510, new_AGEMA_signal_25509}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, new_AGEMA_signal_9256, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, new_AGEMA_signal_8959, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_25516, new_AGEMA_signal_25515, new_AGEMA_signal_25514, new_AGEMA_signal_25513}), .clk (clk), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_25512, new_AGEMA_signal_25511, new_AGEMA_signal_25510, new_AGEMA_signal_25509}), .b ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, new_AGEMA_signal_8965, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, new_AGEMA_signal_9262, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_25516, new_AGEMA_signal_25515, new_AGEMA_signal_25514, new_AGEMA_signal_25513}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, new_AGEMA_signal_8710, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970], Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_25824, new_AGEMA_signal_25823, new_AGEMA_signal_25822, new_AGEMA_signal_25821}), .b ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, new_AGEMA_signal_9256, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, new_AGEMA_signal_9262, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_25828, new_AGEMA_signal_25827, new_AGEMA_signal_25826, new_AGEMA_signal_25825}), .c ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_25832, new_AGEMA_signal_25831, new_AGEMA_signal_25830, new_AGEMA_signal_25829}), .b ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_25836, new_AGEMA_signal_25835, new_AGEMA_signal_25834, new_AGEMA_signal_25833}), .c ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, new_AGEMA_signal_8977, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_25528, new_AGEMA_signal_25527, new_AGEMA_signal_25526, new_AGEMA_signal_25525}), .clk (clk), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, new_AGEMA_signal_8974, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_25532, new_AGEMA_signal_25531, new_AGEMA_signal_25530, new_AGEMA_signal_25529}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, new_AGEMA_signal_9274, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_25528, new_AGEMA_signal_25527, new_AGEMA_signal_25526, new_AGEMA_signal_25525}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, new_AGEMA_signal_8980, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_25532, new_AGEMA_signal_25531, new_AGEMA_signal_25530, new_AGEMA_signal_25529}), .b ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, new_AGEMA_signal_8722, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, new_AGEMA_signal_9280, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_25840, new_AGEMA_signal_25839, new_AGEMA_signal_25838, new_AGEMA_signal_25837}), .b ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_25844, new_AGEMA_signal_25843, new_AGEMA_signal_25842, new_AGEMA_signal_25841}), .c ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_25848, new_AGEMA_signal_25847, new_AGEMA_signal_25846, new_AGEMA_signal_25845}), .b ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, new_AGEMA_signal_9274, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, new_AGEMA_signal_9280, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_25852, new_AGEMA_signal_25851, new_AGEMA_signal_25850, new_AGEMA_signal_25849}), .c ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, new_AGEMA_signal_8992, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_25544, new_AGEMA_signal_25543, new_AGEMA_signal_25542, new_AGEMA_signal_25541}), .clk (clk), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030], Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, new_AGEMA_signal_9286, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, new_AGEMA_signal_8989, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_25548, new_AGEMA_signal_25547, new_AGEMA_signal_25546, new_AGEMA_signal_25545}), .clk (clk), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_25544, new_AGEMA_signal_25543, new_AGEMA_signal_25542, new_AGEMA_signal_25541}), .b ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, new_AGEMA_signal_8995, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, new_AGEMA_signal_9292, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_25548, new_AGEMA_signal_25547, new_AGEMA_signal_25546, new_AGEMA_signal_25545}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, new_AGEMA_signal_8734, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_25856, new_AGEMA_signal_25855, new_AGEMA_signal_25854, new_AGEMA_signal_25853}), .b ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, new_AGEMA_signal_9286, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, new_AGEMA_signal_9292, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_25860, new_AGEMA_signal_25859, new_AGEMA_signal_25858, new_AGEMA_signal_25857}), .c ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_25864, new_AGEMA_signal_25863, new_AGEMA_signal_25862, new_AGEMA_signal_25861}), .b ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_25868, new_AGEMA_signal_25867, new_AGEMA_signal_25866, new_AGEMA_signal_25865}), .c ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, new_AGEMA_signal_9007, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_25560, new_AGEMA_signal_25559, new_AGEMA_signal_25558, new_AGEMA_signal_25557}), .clk (clk), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, new_AGEMA_signal_9004, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_25564, new_AGEMA_signal_25563, new_AGEMA_signal_25562, new_AGEMA_signal_25561}), .clk (clk), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090], Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, new_AGEMA_signal_9304, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_25560, new_AGEMA_signal_25559, new_AGEMA_signal_25558, new_AGEMA_signal_25557}), .b ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, new_AGEMA_signal_9010, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_25564, new_AGEMA_signal_25563, new_AGEMA_signal_25562, new_AGEMA_signal_25561}), .b ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, new_AGEMA_signal_8746, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, new_AGEMA_signal_9310, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_25872, new_AGEMA_signal_25871, new_AGEMA_signal_25870, new_AGEMA_signal_25869}), .b ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_25876, new_AGEMA_signal_25875, new_AGEMA_signal_25874, new_AGEMA_signal_25873}), .c ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_25880, new_AGEMA_signal_25879, new_AGEMA_signal_25878, new_AGEMA_signal_25877}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, new_AGEMA_signal_9304, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, new_AGEMA_signal_9310, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_25884, new_AGEMA_signal_25883, new_AGEMA_signal_25882, new_AGEMA_signal_25881}), .c ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, new_AGEMA_signal_9022, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_25576, new_AGEMA_signal_25575, new_AGEMA_signal_25574, new_AGEMA_signal_25573}), .clk (clk), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, new_AGEMA_signal_9316, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, new_AGEMA_signal_9019, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_25580, new_AGEMA_signal_25579, new_AGEMA_signal_25578, new_AGEMA_signal_25577}), .clk (clk), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_25576, new_AGEMA_signal_25575, new_AGEMA_signal_25574, new_AGEMA_signal_25573}), .b ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, new_AGEMA_signal_9025, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150], Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, new_AGEMA_signal_9322, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_25580, new_AGEMA_signal_25579, new_AGEMA_signal_25578, new_AGEMA_signal_25577}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, new_AGEMA_signal_8758, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_25888, new_AGEMA_signal_25887, new_AGEMA_signal_25886, new_AGEMA_signal_25885}), .b ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, new_AGEMA_signal_9316, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, new_AGEMA_signal_9322, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_25892, new_AGEMA_signal_25891, new_AGEMA_signal_25890, new_AGEMA_signal_25889}), .c ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_25896, new_AGEMA_signal_25895, new_AGEMA_signal_25894, new_AGEMA_signal_25893}), .b ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_25900, new_AGEMA_signal_25899, new_AGEMA_signal_25898, new_AGEMA_signal_25897}), .c ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_25592, new_AGEMA_signal_25591, new_AGEMA_signal_25590, new_AGEMA_signal_25589}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, new_AGEMA_signal_9034, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_25596, new_AGEMA_signal_25595, new_AGEMA_signal_25594, new_AGEMA_signal_25593}), .clk (clk), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, new_AGEMA_signal_9334, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_25592, new_AGEMA_signal_25591, new_AGEMA_signal_25590, new_AGEMA_signal_25589}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, new_AGEMA_signal_9040, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_25596, new_AGEMA_signal_25595, new_AGEMA_signal_25594, new_AGEMA_signal_25593}), .b ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, new_AGEMA_signal_8770, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210], Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, new_AGEMA_signal_9340, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_25904, new_AGEMA_signal_25903, new_AGEMA_signal_25902, new_AGEMA_signal_25901}), .b ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_25908, new_AGEMA_signal_25907, new_AGEMA_signal_25906, new_AGEMA_signal_25905}), .c ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_25912, new_AGEMA_signal_25911, new_AGEMA_signal_25910, new_AGEMA_signal_25909}), .b ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, new_AGEMA_signal_9334, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, new_AGEMA_signal_9340, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_25916, new_AGEMA_signal_25915, new_AGEMA_signal_25914, new_AGEMA_signal_25913}), .c ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, new_AGEMA_signal_9052, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_25608, new_AGEMA_signal_25607, new_AGEMA_signal_25606, new_AGEMA_signal_25605}), .clk (clk), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, new_AGEMA_signal_9346, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_25612, new_AGEMA_signal_25611, new_AGEMA_signal_25610, new_AGEMA_signal_25609}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_25608, new_AGEMA_signal_25607, new_AGEMA_signal_25606, new_AGEMA_signal_25605}), .b ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, new_AGEMA_signal_9352, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_25612, new_AGEMA_signal_25611, new_AGEMA_signal_25610, new_AGEMA_signal_25609}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, new_AGEMA_signal_8782, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_25920, new_AGEMA_signal_25919, new_AGEMA_signal_25918, new_AGEMA_signal_25917}), .b ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, new_AGEMA_signal_9346, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, new_AGEMA_signal_9352, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_25924, new_AGEMA_signal_25923, new_AGEMA_signal_25922, new_AGEMA_signal_25921}), .c ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_25928, new_AGEMA_signal_25927, new_AGEMA_signal_25926, new_AGEMA_signal_25925}), .b ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_25932, new_AGEMA_signal_25931, new_AGEMA_signal_25930, new_AGEMA_signal_25929}), .c ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_25624, new_AGEMA_signal_25623, new_AGEMA_signal_25622, new_AGEMA_signal_25621}), .clk (clk), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270], Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, new_AGEMA_signal_9361, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, new_AGEMA_signal_9064, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_25628, new_AGEMA_signal_25627, new_AGEMA_signal_25626, new_AGEMA_signal_25625}), .clk (clk), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, new_AGEMA_signal_9364, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_25624, new_AGEMA_signal_25623, new_AGEMA_signal_25622, new_AGEMA_signal_25621}), .b ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, new_AGEMA_signal_9070, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, new_AGEMA_signal_9367, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_25628, new_AGEMA_signal_25627, new_AGEMA_signal_25626, new_AGEMA_signal_25625}), .b ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, new_AGEMA_signal_8794, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, new_AGEMA_signal_9370, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_25936, new_AGEMA_signal_25935, new_AGEMA_signal_25934, new_AGEMA_signal_25933}), .b ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, new_AGEMA_signal_9361, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, new_AGEMA_signal_9367, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_25940, new_AGEMA_signal_25939, new_AGEMA_signal_25938, new_AGEMA_signal_25937}), .c ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_25944, new_AGEMA_signal_25943, new_AGEMA_signal_25942, new_AGEMA_signal_25941}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, new_AGEMA_signal_9364, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, new_AGEMA_signal_9370, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_25948, new_AGEMA_signal_25947, new_AGEMA_signal_25946, new_AGEMA_signal_25945}), .c ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, new_AGEMA_signal_9082, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_25640, new_AGEMA_signal_25639, new_AGEMA_signal_25638, new_AGEMA_signal_25637}), .clk (clk), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, new_AGEMA_signal_9376, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_25644, new_AGEMA_signal_25643, new_AGEMA_signal_25642, new_AGEMA_signal_25641}), .clk (clk), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330], Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, new_AGEMA_signal_9379, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_25640, new_AGEMA_signal_25639, new_AGEMA_signal_25638, new_AGEMA_signal_25637}), .b ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, new_AGEMA_signal_9382, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_25644, new_AGEMA_signal_25643, new_AGEMA_signal_25642, new_AGEMA_signal_25641}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, new_AGEMA_signal_8806, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, new_AGEMA_signal_9385, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_25952, new_AGEMA_signal_25951, new_AGEMA_signal_25950, new_AGEMA_signal_25949}), .b ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, new_AGEMA_signal_9376, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, new_AGEMA_signal_9382, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_25956, new_AGEMA_signal_25955, new_AGEMA_signal_25954, new_AGEMA_signal_25953}), .c ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_25960, new_AGEMA_signal_25959, new_AGEMA_signal_25958, new_AGEMA_signal_25957}), .b ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, new_AGEMA_signal_9379, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, new_AGEMA_signal_9385, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_25964, new_AGEMA_signal_25963, new_AGEMA_signal_25962, new_AGEMA_signal_25961}), .c ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_25656, new_AGEMA_signal_25655, new_AGEMA_signal_25654, new_AGEMA_signal_25653}), .clk (clk), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, new_AGEMA_signal_9391, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, new_AGEMA_signal_9094, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_25660, new_AGEMA_signal_25659, new_AGEMA_signal_25658, new_AGEMA_signal_25657}), .clk (clk), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, new_AGEMA_signal_9394, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_25656, new_AGEMA_signal_25655, new_AGEMA_signal_25654, new_AGEMA_signal_25653}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, new_AGEMA_signal_9100, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390], Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, new_AGEMA_signal_9397, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_25660, new_AGEMA_signal_25659, new_AGEMA_signal_25658, new_AGEMA_signal_25657}), .b ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, new_AGEMA_signal_8818, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, new_AGEMA_signal_9400, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_25968, new_AGEMA_signal_25967, new_AGEMA_signal_25966, new_AGEMA_signal_25965}), .b ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, new_AGEMA_signal_9391, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, new_AGEMA_signal_9397, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_25972, new_AGEMA_signal_25971, new_AGEMA_signal_25970, new_AGEMA_signal_25969}), .c ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_25976, new_AGEMA_signal_25975, new_AGEMA_signal_25974, new_AGEMA_signal_25973}), .b ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, new_AGEMA_signal_9394, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, new_AGEMA_signal_9400, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_25980, new_AGEMA_signal_25979, new_AGEMA_signal_25978, new_AGEMA_signal_25977}), .c ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, new_AGEMA_signal_9112, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_25672, new_AGEMA_signal_25671, new_AGEMA_signal_25670, new_AGEMA_signal_25669}), .clk (clk), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, new_AGEMA_signal_9406, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_25676, new_AGEMA_signal_25675, new_AGEMA_signal_25674, new_AGEMA_signal_25673}), .clk (clk), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, new_AGEMA_signal_9409, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_25672, new_AGEMA_signal_25671, new_AGEMA_signal_25670, new_AGEMA_signal_25669}), .b ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, new_AGEMA_signal_9412, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_25676, new_AGEMA_signal_25675, new_AGEMA_signal_25674, new_AGEMA_signal_25673}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, new_AGEMA_signal_8830, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450], Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, new_AGEMA_signal_9415, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_25984, new_AGEMA_signal_25983, new_AGEMA_signal_25982, new_AGEMA_signal_25981}), .b ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, new_AGEMA_signal_9406, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, new_AGEMA_signal_9412, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_25988, new_AGEMA_signal_25987, new_AGEMA_signal_25986, new_AGEMA_signal_25985}), .c ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_25992, new_AGEMA_signal_25991, new_AGEMA_signal_25990, new_AGEMA_signal_25989}), .b ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, new_AGEMA_signal_9409, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, new_AGEMA_signal_9415, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_25996, new_AGEMA_signal_25995, new_AGEMA_signal_25994, new_AGEMA_signal_25993}), .c ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_25688, new_AGEMA_signal_25687, new_AGEMA_signal_25686, new_AGEMA_signal_25685}), .clk (clk), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, new_AGEMA_signal_9421, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, new_AGEMA_signal_9124, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_25692, new_AGEMA_signal_25691, new_AGEMA_signal_25690, new_AGEMA_signal_25689}), .clk (clk), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, new_AGEMA_signal_9424, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_25688, new_AGEMA_signal_25687, new_AGEMA_signal_25686, new_AGEMA_signal_25685}), .b ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, new_AGEMA_signal_9130, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, new_AGEMA_signal_9427, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_25692, new_AGEMA_signal_25691, new_AGEMA_signal_25690, new_AGEMA_signal_25689}), .b ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, new_AGEMA_signal_8842, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, new_AGEMA_signal_9430, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_26000, new_AGEMA_signal_25999, new_AGEMA_signal_25998, new_AGEMA_signal_25997}), .b ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, new_AGEMA_signal_9421, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, new_AGEMA_signal_9427, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_26004, new_AGEMA_signal_26003, new_AGEMA_signal_26002, new_AGEMA_signal_26001}), .c ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_26008, new_AGEMA_signal_26007, new_AGEMA_signal_26006, new_AGEMA_signal_26005}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, new_AGEMA_signal_9424, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, new_AGEMA_signal_9430, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_26012, new_AGEMA_signal_26011, new_AGEMA_signal_26010, new_AGEMA_signal_26009}), .c ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, new_AGEMA_signal_9142, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_25704, new_AGEMA_signal_25703, new_AGEMA_signal_25702, new_AGEMA_signal_25701}), .clk (clk), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510], Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, new_AGEMA_signal_9436, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_25708, new_AGEMA_signal_25707, new_AGEMA_signal_25706, new_AGEMA_signal_25705}), .clk (clk), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_25704, new_AGEMA_signal_25703, new_AGEMA_signal_25702, new_AGEMA_signal_25701}), .b ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, new_AGEMA_signal_9442, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_25708, new_AGEMA_signal_25707, new_AGEMA_signal_25706, new_AGEMA_signal_25705}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, new_AGEMA_signal_8854, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_26016, new_AGEMA_signal_26015, new_AGEMA_signal_26014, new_AGEMA_signal_26013}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, new_AGEMA_signal_9436, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, new_AGEMA_signal_9442, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_26020, new_AGEMA_signal_26019, new_AGEMA_signal_26018, new_AGEMA_signal_26017}), .c ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_26024, new_AGEMA_signal_26023, new_AGEMA_signal_26022, new_AGEMA_signal_26021}), .b ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_26028, new_AGEMA_signal_26027, new_AGEMA_signal_26026, new_AGEMA_signal_26025}), .c ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_25720, new_AGEMA_signal_25719, new_AGEMA_signal_25718, new_AGEMA_signal_25717}), .clk (clk), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, new_AGEMA_signal_9154, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_25724, new_AGEMA_signal_25723, new_AGEMA_signal_25722, new_AGEMA_signal_25721}), .clk (clk), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570], Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, new_AGEMA_signal_9454, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_25720, new_AGEMA_signal_25719, new_AGEMA_signal_25718, new_AGEMA_signal_25717}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, new_AGEMA_signal_9160, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_25724, new_AGEMA_signal_25723, new_AGEMA_signal_25722, new_AGEMA_signal_25721}), .b ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, new_AGEMA_signal_8866, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, new_AGEMA_signal_9460, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_26032, new_AGEMA_signal_26031, new_AGEMA_signal_26030, new_AGEMA_signal_26029}), .b ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_26036, new_AGEMA_signal_26035, new_AGEMA_signal_26034, new_AGEMA_signal_26033}), .c ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_26040, new_AGEMA_signal_26039, new_AGEMA_signal_26038, new_AGEMA_signal_26037}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, new_AGEMA_signal_9454, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, new_AGEMA_signal_9460, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_26044, new_AGEMA_signal_26043, new_AGEMA_signal_26042, new_AGEMA_signal_26041}), .c ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, new_AGEMA_signal_9172, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_25736, new_AGEMA_signal_25735, new_AGEMA_signal_25734, new_AGEMA_signal_25733}), .clk (clk), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, new_AGEMA_signal_9466, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_25740, new_AGEMA_signal_25739, new_AGEMA_signal_25738, new_AGEMA_signal_25737}), .clk (clk), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_25736, new_AGEMA_signal_25735, new_AGEMA_signal_25734, new_AGEMA_signal_25733}), .b ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630], Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, new_AGEMA_signal_9472, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_25740, new_AGEMA_signal_25739, new_AGEMA_signal_25738, new_AGEMA_signal_25737}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, new_AGEMA_signal_8878, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_26048, new_AGEMA_signal_26047, new_AGEMA_signal_26046, new_AGEMA_signal_26045}), .b ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, new_AGEMA_signal_9466, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, new_AGEMA_signal_9472, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_26052, new_AGEMA_signal_26051, new_AGEMA_signal_26050, new_AGEMA_signal_26049}), .c ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_26056, new_AGEMA_signal_26055, new_AGEMA_signal_26054, new_AGEMA_signal_26053}), .b ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_26060, new_AGEMA_signal_26059, new_AGEMA_signal_26058, new_AGEMA_signal_26057}), .c ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, new_AGEMA_signal_8887, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_25752, new_AGEMA_signal_25751, new_AGEMA_signal_25750, new_AGEMA_signal_25749}), .clk (clk), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, new_AGEMA_signal_9181, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, new_AGEMA_signal_8884, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_25756, new_AGEMA_signal_25755, new_AGEMA_signal_25754, new_AGEMA_signal_25753}), .clk (clk), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, new_AGEMA_signal_9184, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_25752, new_AGEMA_signal_25751, new_AGEMA_signal_25750, new_AGEMA_signal_25749}), .b ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, new_AGEMA_signal_8890, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, new_AGEMA_signal_9187, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_25756, new_AGEMA_signal_25755, new_AGEMA_signal_25754, new_AGEMA_signal_25753}), .b ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, new_AGEMA_signal_8650, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690], Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, new_AGEMA_signal_9190, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_26064, new_AGEMA_signal_26063, new_AGEMA_signal_26062, new_AGEMA_signal_26061}), .b ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, new_AGEMA_signal_9181, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, new_AGEMA_signal_9187, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_26068, new_AGEMA_signal_26067, new_AGEMA_signal_26066, new_AGEMA_signal_26065}), .c ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_26072, new_AGEMA_signal_26071, new_AGEMA_signal_26070, new_AGEMA_signal_26069}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, new_AGEMA_signal_9184, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, new_AGEMA_signal_9190, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_26076, new_AGEMA_signal_26075, new_AGEMA_signal_26074, new_AGEMA_signal_26073}), .c ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, new_AGEMA_signal_8902, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_25768, new_AGEMA_signal_25767, new_AGEMA_signal_25766, new_AGEMA_signal_25765}), .clk (clk), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, new_AGEMA_signal_9196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, new_AGEMA_signal_8899, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_25772, new_AGEMA_signal_25771, new_AGEMA_signal_25770, new_AGEMA_signal_25769}), .clk (clk), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, new_AGEMA_signal_9199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_25768, new_AGEMA_signal_25767, new_AGEMA_signal_25766, new_AGEMA_signal_25765}), .b ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, new_AGEMA_signal_8905, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, new_AGEMA_signal_9202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_25772, new_AGEMA_signal_25771, new_AGEMA_signal_25770, new_AGEMA_signal_25769}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, new_AGEMA_signal_8662, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, new_AGEMA_signal_9205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_26080, new_AGEMA_signal_26079, new_AGEMA_signal_26078, new_AGEMA_signal_26077}), .b ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, new_AGEMA_signal_9196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, new_AGEMA_signal_9202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_26084, new_AGEMA_signal_26083, new_AGEMA_signal_26082, new_AGEMA_signal_26081}), .c ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_26088, new_AGEMA_signal_26087, new_AGEMA_signal_26086, new_AGEMA_signal_26085}), .b ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, new_AGEMA_signal_9199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, new_AGEMA_signal_9205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_26092, new_AGEMA_signal_26091, new_AGEMA_signal_26090, new_AGEMA_signal_26089}), .c ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, new_AGEMA_signal_8917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_25784, new_AGEMA_signal_25783, new_AGEMA_signal_25782, new_AGEMA_signal_25781}), .clk (clk), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750], Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, new_AGEMA_signal_9211, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, new_AGEMA_signal_8914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_25788, new_AGEMA_signal_25787, new_AGEMA_signal_25786, new_AGEMA_signal_25785}), .clk (clk), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, new_AGEMA_signal_9214, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_25784, new_AGEMA_signal_25783, new_AGEMA_signal_25782, new_AGEMA_signal_25781}), .b ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, new_AGEMA_signal_8920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, new_AGEMA_signal_9217, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_25788, new_AGEMA_signal_25787, new_AGEMA_signal_25786, new_AGEMA_signal_25785}), .b ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, new_AGEMA_signal_8674, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, new_AGEMA_signal_9220, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_26096, new_AGEMA_signal_26095, new_AGEMA_signal_26094, new_AGEMA_signal_26093}), .b ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, new_AGEMA_signal_9211, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, new_AGEMA_signal_9217, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_26100, new_AGEMA_signal_26099, new_AGEMA_signal_26098, new_AGEMA_signal_26097}), .c ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_26104, new_AGEMA_signal_26103, new_AGEMA_signal_26102, new_AGEMA_signal_26101}), .b ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, new_AGEMA_signal_9214, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, new_AGEMA_signal_9220, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_26108, new_AGEMA_signal_26107, new_AGEMA_signal_26106, new_AGEMA_signal_26105}), .c ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, new_AGEMA_signal_8932, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_25800, new_AGEMA_signal_25799, new_AGEMA_signal_25798, new_AGEMA_signal_25797}), .clk (clk), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, new_AGEMA_signal_9226, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, new_AGEMA_signal_8929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_25804, new_AGEMA_signal_25803, new_AGEMA_signal_25802, new_AGEMA_signal_25801}), .clk (clk), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810], Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, new_AGEMA_signal_9229, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_25800, new_AGEMA_signal_25799, new_AGEMA_signal_25798, new_AGEMA_signal_25797}), .b ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, new_AGEMA_signal_8935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, new_AGEMA_signal_9232, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_25804, new_AGEMA_signal_25803, new_AGEMA_signal_25802, new_AGEMA_signal_25801}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, new_AGEMA_signal_8686, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, new_AGEMA_signal_9235, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_26112, new_AGEMA_signal_26111, new_AGEMA_signal_26110, new_AGEMA_signal_26109}), .b ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, new_AGEMA_signal_9226, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, new_AGEMA_signal_9232, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_26116, new_AGEMA_signal_26115, new_AGEMA_signal_26114, new_AGEMA_signal_26113}), .c ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_26120, new_AGEMA_signal_26119, new_AGEMA_signal_26118, new_AGEMA_signal_26117}), .b ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, new_AGEMA_signal_9229, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, new_AGEMA_signal_9235, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_26124, new_AGEMA_signal_26123, new_AGEMA_signal_26122, new_AGEMA_signal_26121}), .c ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C (clk), .D (new_AGEMA_signal_25485), .Q (new_AGEMA_signal_25805) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_25486), .Q (new_AGEMA_signal_25806) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_25487), .Q (new_AGEMA_signal_25807) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_25488), .Q (new_AGEMA_signal_25808) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_25809) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_8953), .Q (new_AGEMA_signal_25810) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_8954), .Q (new_AGEMA_signal_25811) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_8955), .Q (new_AGEMA_signal_25812) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C (clk), .D (new_AGEMA_signal_25489), .Q (new_AGEMA_signal_25813) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_25490), .Q (new_AGEMA_signal_25814) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_25491), .Q (new_AGEMA_signal_25815) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_25492), .Q (new_AGEMA_signal_25816) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_25817) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_9253), .Q (new_AGEMA_signal_25818) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_9254), .Q (new_AGEMA_signal_25819) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_9255), .Q (new_AGEMA_signal_25820) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C (clk), .D (new_AGEMA_signal_25501), .Q (new_AGEMA_signal_25821) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_25502), .Q (new_AGEMA_signal_25822) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_25503), .Q (new_AGEMA_signal_25823) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_25504), .Q (new_AGEMA_signal_25824) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_25825) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_8968), .Q (new_AGEMA_signal_25826) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_8969), .Q (new_AGEMA_signal_25827) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_8970), .Q (new_AGEMA_signal_25828) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C (clk), .D (new_AGEMA_signal_25505), .Q (new_AGEMA_signal_25829) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_25506), .Q (new_AGEMA_signal_25830) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_25507), .Q (new_AGEMA_signal_25831) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_25508), .Q (new_AGEMA_signal_25832) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_25833) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_9268), .Q (new_AGEMA_signal_25834) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_9269), .Q (new_AGEMA_signal_25835) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_9270), .Q (new_AGEMA_signal_25836) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C (clk), .D (new_AGEMA_signal_25517), .Q (new_AGEMA_signal_25837) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_25518), .Q (new_AGEMA_signal_25838) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_25519), .Q (new_AGEMA_signal_25839) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_25520), .Q (new_AGEMA_signal_25840) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_25841) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_8983), .Q (new_AGEMA_signal_25842) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_8984), .Q (new_AGEMA_signal_25843) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_8985), .Q (new_AGEMA_signal_25844) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C (clk), .D (new_AGEMA_signal_25521), .Q (new_AGEMA_signal_25845) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_25522), .Q (new_AGEMA_signal_25846) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_25523), .Q (new_AGEMA_signal_25847) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_25524), .Q (new_AGEMA_signal_25848) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_25849) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_9283), .Q (new_AGEMA_signal_25850) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_9284), .Q (new_AGEMA_signal_25851) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_9285), .Q (new_AGEMA_signal_25852) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C (clk), .D (new_AGEMA_signal_25533), .Q (new_AGEMA_signal_25853) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_25534), .Q (new_AGEMA_signal_25854) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_25535), .Q (new_AGEMA_signal_25855) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_25536), .Q (new_AGEMA_signal_25856) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_25857) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_8998), .Q (new_AGEMA_signal_25858) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_8999), .Q (new_AGEMA_signal_25859) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_9000), .Q (new_AGEMA_signal_25860) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C (clk), .D (new_AGEMA_signal_25537), .Q (new_AGEMA_signal_25861) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_25538), .Q (new_AGEMA_signal_25862) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_25539), .Q (new_AGEMA_signal_25863) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_25540), .Q (new_AGEMA_signal_25864) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_25865) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_9298), .Q (new_AGEMA_signal_25866) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_9299), .Q (new_AGEMA_signal_25867) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_9300), .Q (new_AGEMA_signal_25868) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C (clk), .D (new_AGEMA_signal_25549), .Q (new_AGEMA_signal_25869) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_25550), .Q (new_AGEMA_signal_25870) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_25551), .Q (new_AGEMA_signal_25871) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_25552), .Q (new_AGEMA_signal_25872) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M33), .Q (new_AGEMA_signal_25873) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_9013), .Q (new_AGEMA_signal_25874) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_9014), .Q (new_AGEMA_signal_25875) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_9015), .Q (new_AGEMA_signal_25876) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C (clk), .D (new_AGEMA_signal_25553), .Q (new_AGEMA_signal_25877) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_25554), .Q (new_AGEMA_signal_25878) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_25555), .Q (new_AGEMA_signal_25879) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_25556), .Q (new_AGEMA_signal_25880) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M36), .Q (new_AGEMA_signal_25881) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_9313), .Q (new_AGEMA_signal_25882) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_9314), .Q (new_AGEMA_signal_25883) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_9315), .Q (new_AGEMA_signal_25884) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C (clk), .D (new_AGEMA_signal_25565), .Q (new_AGEMA_signal_25885) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_25566), .Q (new_AGEMA_signal_25886) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_25567), .Q (new_AGEMA_signal_25887) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_25568), .Q (new_AGEMA_signal_25888) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M33), .Q (new_AGEMA_signal_25889) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_9028), .Q (new_AGEMA_signal_25890) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_9029), .Q (new_AGEMA_signal_25891) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_9030), .Q (new_AGEMA_signal_25892) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C (clk), .D (new_AGEMA_signal_25569), .Q (new_AGEMA_signal_25893) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_25570), .Q (new_AGEMA_signal_25894) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_25571), .Q (new_AGEMA_signal_25895) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_25572), .Q (new_AGEMA_signal_25896) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M36), .Q (new_AGEMA_signal_25897) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_9328), .Q (new_AGEMA_signal_25898) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_9329), .Q (new_AGEMA_signal_25899) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_9330), .Q (new_AGEMA_signal_25900) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C (clk), .D (new_AGEMA_signal_25581), .Q (new_AGEMA_signal_25901) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_25582), .Q (new_AGEMA_signal_25902) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_25583), .Q (new_AGEMA_signal_25903) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_25584), .Q (new_AGEMA_signal_25904) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M33), .Q (new_AGEMA_signal_25905) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_9043), .Q (new_AGEMA_signal_25906) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_9044), .Q (new_AGEMA_signal_25907) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_9045), .Q (new_AGEMA_signal_25908) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C (clk), .D (new_AGEMA_signal_25585), .Q (new_AGEMA_signal_25909) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_25586), .Q (new_AGEMA_signal_25910) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_25587), .Q (new_AGEMA_signal_25911) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_25588), .Q (new_AGEMA_signal_25912) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M36), .Q (new_AGEMA_signal_25913) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_9343), .Q (new_AGEMA_signal_25914) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_9344), .Q (new_AGEMA_signal_25915) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_9345), .Q (new_AGEMA_signal_25916) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C (clk), .D (new_AGEMA_signal_25597), .Q (new_AGEMA_signal_25917) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_25598), .Q (new_AGEMA_signal_25918) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_25599), .Q (new_AGEMA_signal_25919) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_25600), .Q (new_AGEMA_signal_25920) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M33), .Q (new_AGEMA_signal_25921) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_9058), .Q (new_AGEMA_signal_25922) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_9059), .Q (new_AGEMA_signal_25923) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_9060), .Q (new_AGEMA_signal_25924) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C (clk), .D (new_AGEMA_signal_25601), .Q (new_AGEMA_signal_25925) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_25602), .Q (new_AGEMA_signal_25926) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_25603), .Q (new_AGEMA_signal_25927) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_25604), .Q (new_AGEMA_signal_25928) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M36), .Q (new_AGEMA_signal_25929) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_9358), .Q (new_AGEMA_signal_25930) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_9359), .Q (new_AGEMA_signal_25931) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_9360), .Q (new_AGEMA_signal_25932) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C (clk), .D (new_AGEMA_signal_25613), .Q (new_AGEMA_signal_25933) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_25614), .Q (new_AGEMA_signal_25934) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_25615), .Q (new_AGEMA_signal_25935) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_25616), .Q (new_AGEMA_signal_25936) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M33), .Q (new_AGEMA_signal_25937) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_9073), .Q (new_AGEMA_signal_25938) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_9074), .Q (new_AGEMA_signal_25939) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_9075), .Q (new_AGEMA_signal_25940) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C (clk), .D (new_AGEMA_signal_25617), .Q (new_AGEMA_signal_25941) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_25618), .Q (new_AGEMA_signal_25942) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_25619), .Q (new_AGEMA_signal_25943) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_25620), .Q (new_AGEMA_signal_25944) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M36), .Q (new_AGEMA_signal_25945) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_9373), .Q (new_AGEMA_signal_25946) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_9374), .Q (new_AGEMA_signal_25947) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_9375), .Q (new_AGEMA_signal_25948) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C (clk), .D (new_AGEMA_signal_25629), .Q (new_AGEMA_signal_25949) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_25630), .Q (new_AGEMA_signal_25950) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_25631), .Q (new_AGEMA_signal_25951) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_25632), .Q (new_AGEMA_signal_25952) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M33), .Q (new_AGEMA_signal_25953) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_9088), .Q (new_AGEMA_signal_25954) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_9089), .Q (new_AGEMA_signal_25955) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_9090), .Q (new_AGEMA_signal_25956) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C (clk), .D (new_AGEMA_signal_25633), .Q (new_AGEMA_signal_25957) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_25634), .Q (new_AGEMA_signal_25958) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_25635), .Q (new_AGEMA_signal_25959) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_25636), .Q (new_AGEMA_signal_25960) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M36), .Q (new_AGEMA_signal_25961) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_9388), .Q (new_AGEMA_signal_25962) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_9389), .Q (new_AGEMA_signal_25963) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_9390), .Q (new_AGEMA_signal_25964) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C (clk), .D (new_AGEMA_signal_25645), .Q (new_AGEMA_signal_25965) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_25646), .Q (new_AGEMA_signal_25966) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_25647), .Q (new_AGEMA_signal_25967) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_25648), .Q (new_AGEMA_signal_25968) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M33), .Q (new_AGEMA_signal_25969) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_9103), .Q (new_AGEMA_signal_25970) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_9104), .Q (new_AGEMA_signal_25971) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_9105), .Q (new_AGEMA_signal_25972) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C (clk), .D (new_AGEMA_signal_25649), .Q (new_AGEMA_signal_25973) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_25650), .Q (new_AGEMA_signal_25974) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_25651), .Q (new_AGEMA_signal_25975) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_25652), .Q (new_AGEMA_signal_25976) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M36), .Q (new_AGEMA_signal_25977) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_9403), .Q (new_AGEMA_signal_25978) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_9404), .Q (new_AGEMA_signal_25979) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_9405), .Q (new_AGEMA_signal_25980) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C (clk), .D (new_AGEMA_signal_25661), .Q (new_AGEMA_signal_25981) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_25662), .Q (new_AGEMA_signal_25982) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_25663), .Q (new_AGEMA_signal_25983) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_25664), .Q (new_AGEMA_signal_25984) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M33), .Q (new_AGEMA_signal_25985) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_9118), .Q (new_AGEMA_signal_25986) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_9119), .Q (new_AGEMA_signal_25987) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_9120), .Q (new_AGEMA_signal_25988) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C (clk), .D (new_AGEMA_signal_25665), .Q (new_AGEMA_signal_25989) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_25666), .Q (new_AGEMA_signal_25990) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_25667), .Q (new_AGEMA_signal_25991) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_25668), .Q (new_AGEMA_signal_25992) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M36), .Q (new_AGEMA_signal_25993) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_9418), .Q (new_AGEMA_signal_25994) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_9419), .Q (new_AGEMA_signal_25995) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_9420), .Q (new_AGEMA_signal_25996) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C (clk), .D (new_AGEMA_signal_25677), .Q (new_AGEMA_signal_25997) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_25678), .Q (new_AGEMA_signal_25998) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_25679), .Q (new_AGEMA_signal_25999) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_25680), .Q (new_AGEMA_signal_26000) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M33), .Q (new_AGEMA_signal_26001) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_9133), .Q (new_AGEMA_signal_26002) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_9134), .Q (new_AGEMA_signal_26003) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_9135), .Q (new_AGEMA_signal_26004) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C (clk), .D (new_AGEMA_signal_25681), .Q (new_AGEMA_signal_26005) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_25682), .Q (new_AGEMA_signal_26006) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_25683), .Q (new_AGEMA_signal_26007) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_25684), .Q (new_AGEMA_signal_26008) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M36), .Q (new_AGEMA_signal_26009) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_9433), .Q (new_AGEMA_signal_26010) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_9434), .Q (new_AGEMA_signal_26011) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_9435), .Q (new_AGEMA_signal_26012) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C (clk), .D (new_AGEMA_signal_25693), .Q (new_AGEMA_signal_26013) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_25694), .Q (new_AGEMA_signal_26014) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_25695), .Q (new_AGEMA_signal_26015) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_25696), .Q (new_AGEMA_signal_26016) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M33), .Q (new_AGEMA_signal_26017) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_9148), .Q (new_AGEMA_signal_26018) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_9149), .Q (new_AGEMA_signal_26019) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_9150), .Q (new_AGEMA_signal_26020) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C (clk), .D (new_AGEMA_signal_25697), .Q (new_AGEMA_signal_26021) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_25698), .Q (new_AGEMA_signal_26022) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_25699), .Q (new_AGEMA_signal_26023) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_25700), .Q (new_AGEMA_signal_26024) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M36), .Q (new_AGEMA_signal_26025) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_9448), .Q (new_AGEMA_signal_26026) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_9449), .Q (new_AGEMA_signal_26027) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_9450), .Q (new_AGEMA_signal_26028) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C (clk), .D (new_AGEMA_signal_25709), .Q (new_AGEMA_signal_26029) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_25710), .Q (new_AGEMA_signal_26030) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_25711), .Q (new_AGEMA_signal_26031) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_25712), .Q (new_AGEMA_signal_26032) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M33), .Q (new_AGEMA_signal_26033) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_9163), .Q (new_AGEMA_signal_26034) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_9164), .Q (new_AGEMA_signal_26035) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_9165), .Q (new_AGEMA_signal_26036) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C (clk), .D (new_AGEMA_signal_25713), .Q (new_AGEMA_signal_26037) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_25714), .Q (new_AGEMA_signal_26038) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_25715), .Q (new_AGEMA_signal_26039) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_25716), .Q (new_AGEMA_signal_26040) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M36), .Q (new_AGEMA_signal_26041) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_9463), .Q (new_AGEMA_signal_26042) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_9464), .Q (new_AGEMA_signal_26043) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_9465), .Q (new_AGEMA_signal_26044) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C (clk), .D (new_AGEMA_signal_25725), .Q (new_AGEMA_signal_26045) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_25726), .Q (new_AGEMA_signal_26046) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_25727), .Q (new_AGEMA_signal_26047) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_25728), .Q (new_AGEMA_signal_26048) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M33), .Q (new_AGEMA_signal_26049) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_9178), .Q (new_AGEMA_signal_26050) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_9179), .Q (new_AGEMA_signal_26051) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_9180), .Q (new_AGEMA_signal_26052) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C (clk), .D (new_AGEMA_signal_25729), .Q (new_AGEMA_signal_26053) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_25730), .Q (new_AGEMA_signal_26054) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_25731), .Q (new_AGEMA_signal_26055) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_25732), .Q (new_AGEMA_signal_26056) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M36), .Q (new_AGEMA_signal_26057) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_9478), .Q (new_AGEMA_signal_26058) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_9479), .Q (new_AGEMA_signal_26059) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_9480), .Q (new_AGEMA_signal_26060) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C (clk), .D (new_AGEMA_signal_25741), .Q (new_AGEMA_signal_26061) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_25742), .Q (new_AGEMA_signal_26062) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_25743), .Q (new_AGEMA_signal_26063) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_25744), .Q (new_AGEMA_signal_26064) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_26065) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_8893), .Q (new_AGEMA_signal_26066) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_8894), .Q (new_AGEMA_signal_26067) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_8895), .Q (new_AGEMA_signal_26068) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C (clk), .D (new_AGEMA_signal_25745), .Q (new_AGEMA_signal_26069) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_25746), .Q (new_AGEMA_signal_26070) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_25747), .Q (new_AGEMA_signal_26071) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_25748), .Q (new_AGEMA_signal_26072) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_26073) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_9193), .Q (new_AGEMA_signal_26074) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_9194), .Q (new_AGEMA_signal_26075) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_9195), .Q (new_AGEMA_signal_26076) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C (clk), .D (new_AGEMA_signal_25757), .Q (new_AGEMA_signal_26077) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_25758), .Q (new_AGEMA_signal_26078) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_25759), .Q (new_AGEMA_signal_26079) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_25760), .Q (new_AGEMA_signal_26080) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_26081) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_8908), .Q (new_AGEMA_signal_26082) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_8909), .Q (new_AGEMA_signal_26083) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_8910), .Q (new_AGEMA_signal_26084) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C (clk), .D (new_AGEMA_signal_25761), .Q (new_AGEMA_signal_26085) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_25762), .Q (new_AGEMA_signal_26086) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_25763), .Q (new_AGEMA_signal_26087) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_25764), .Q (new_AGEMA_signal_26088) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_26089) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_9208), .Q (new_AGEMA_signal_26090) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_9209), .Q (new_AGEMA_signal_26091) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_9210), .Q (new_AGEMA_signal_26092) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C (clk), .D (new_AGEMA_signal_25773), .Q (new_AGEMA_signal_26093) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_25774), .Q (new_AGEMA_signal_26094) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_25775), .Q (new_AGEMA_signal_26095) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_25776), .Q (new_AGEMA_signal_26096) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_26097) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_8923), .Q (new_AGEMA_signal_26098) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_8924), .Q (new_AGEMA_signal_26099) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_8925), .Q (new_AGEMA_signal_26100) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C (clk), .D (new_AGEMA_signal_25777), .Q (new_AGEMA_signal_26101) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_25778), .Q (new_AGEMA_signal_26102) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_25779), .Q (new_AGEMA_signal_26103) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_25780), .Q (new_AGEMA_signal_26104) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_26105) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_9223), .Q (new_AGEMA_signal_26106) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_9224), .Q (new_AGEMA_signal_26107) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_9225), .Q (new_AGEMA_signal_26108) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C (clk), .D (new_AGEMA_signal_25789), .Q (new_AGEMA_signal_26109) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_25790), .Q (new_AGEMA_signal_26110) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_25791), .Q (new_AGEMA_signal_26111) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_25792), .Q (new_AGEMA_signal_26112) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_26113) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_8938), .Q (new_AGEMA_signal_26114) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_8939), .Q (new_AGEMA_signal_26115) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_8940), .Q (new_AGEMA_signal_26116) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C (clk), .D (new_AGEMA_signal_25793), .Q (new_AGEMA_signal_26117) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_25794), .Q (new_AGEMA_signal_26118) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_25795), .Q (new_AGEMA_signal_26119) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_25796), .Q (new_AGEMA_signal_26120) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_26121) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_9238), .Q (new_AGEMA_signal_26122) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_9239), .Q (new_AGEMA_signal_26123) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_9240), .Q (new_AGEMA_signal_26124) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_26126), .Q (new_AGEMA_signal_26127) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_26130), .Q (new_AGEMA_signal_26131) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_26134), .Q (new_AGEMA_signal_26135) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_26138), .Q (new_AGEMA_signal_26139) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_26142), .Q (new_AGEMA_signal_26143) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_26146), .Q (new_AGEMA_signal_26147) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_26150), .Q (new_AGEMA_signal_26151) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_26154), .Q (new_AGEMA_signal_26155) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_26158), .Q (new_AGEMA_signal_26159) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_26162), .Q (new_AGEMA_signal_26163) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_26166), .Q (new_AGEMA_signal_26167) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_26170), .Q (new_AGEMA_signal_26171) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_26174), .Q (new_AGEMA_signal_26175) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_26178), .Q (new_AGEMA_signal_26179) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_26182), .Q (new_AGEMA_signal_26183) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_26186), .Q (new_AGEMA_signal_26187) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_26190), .Q (new_AGEMA_signal_26191) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_26194), .Q (new_AGEMA_signal_26195) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_26198), .Q (new_AGEMA_signal_26199) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_26202), .Q (new_AGEMA_signal_26203) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_26206), .Q (new_AGEMA_signal_26207) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_26210), .Q (new_AGEMA_signal_26211) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_26214), .Q (new_AGEMA_signal_26215) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_26218), .Q (new_AGEMA_signal_26219) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_26222), .Q (new_AGEMA_signal_26223) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_26226), .Q (new_AGEMA_signal_26227) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_26230), .Q (new_AGEMA_signal_26231) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_26234), .Q (new_AGEMA_signal_26235) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_26238), .Q (new_AGEMA_signal_26239) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_26242), .Q (new_AGEMA_signal_26243) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_26246), .Q (new_AGEMA_signal_26247) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_26250), .Q (new_AGEMA_signal_26251) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_26254), .Q (new_AGEMA_signal_26255) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_26258), .Q (new_AGEMA_signal_26259) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_26262), .Q (new_AGEMA_signal_26263) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_26266), .Q (new_AGEMA_signal_26267) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_26270), .Q (new_AGEMA_signal_26271) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_26274), .Q (new_AGEMA_signal_26275) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_26278), .Q (new_AGEMA_signal_26279) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_26282), .Q (new_AGEMA_signal_26283) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_26286), .Q (new_AGEMA_signal_26287) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_26290), .Q (new_AGEMA_signal_26291) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_26294), .Q (new_AGEMA_signal_26295) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_26298), .Q (new_AGEMA_signal_26299) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_26302), .Q (new_AGEMA_signal_26303) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_26306), .Q (new_AGEMA_signal_26307) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_26310), .Q (new_AGEMA_signal_26311) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_26314), .Q (new_AGEMA_signal_26315) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_26318), .Q (new_AGEMA_signal_26319) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_26322), .Q (new_AGEMA_signal_26323) ) ;
    buf_clk new_AGEMA_reg_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_26326), .Q (new_AGEMA_signal_26327) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_26330), .Q (new_AGEMA_signal_26331) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_26334), .Q (new_AGEMA_signal_26335) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_26338), .Q (new_AGEMA_signal_26339) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_26342), .Q (new_AGEMA_signal_26343) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_26346), .Q (new_AGEMA_signal_26347) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_26350), .Q (new_AGEMA_signal_26351) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_26354), .Q (new_AGEMA_signal_26355) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_26358), .Q (new_AGEMA_signal_26359) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_26362), .Q (new_AGEMA_signal_26363) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_26366), .Q (new_AGEMA_signal_26367) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_26370), .Q (new_AGEMA_signal_26371) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_26374), .Q (new_AGEMA_signal_26375) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_26378), .Q (new_AGEMA_signal_26379) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_26382), .Q (new_AGEMA_signal_26383) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_26386), .Q (new_AGEMA_signal_26387) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_26390), .Q (new_AGEMA_signal_26391) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_26394), .Q (new_AGEMA_signal_26395) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_26398), .Q (new_AGEMA_signal_26399) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_26402), .Q (new_AGEMA_signal_26403) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_26406), .Q (new_AGEMA_signal_26407) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_26410), .Q (new_AGEMA_signal_26411) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_26414), .Q (new_AGEMA_signal_26415) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_26418), .Q (new_AGEMA_signal_26419) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_26422), .Q (new_AGEMA_signal_26423) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_26426), .Q (new_AGEMA_signal_26427) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_26430), .Q (new_AGEMA_signal_26431) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_26434), .Q (new_AGEMA_signal_26435) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_26438), .Q (new_AGEMA_signal_26439) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_26442), .Q (new_AGEMA_signal_26443) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_26446), .Q (new_AGEMA_signal_26447) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_26450), .Q (new_AGEMA_signal_26451) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_26454), .Q (new_AGEMA_signal_26455) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_26458), .Q (new_AGEMA_signal_26459) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_26462), .Q (new_AGEMA_signal_26463) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_26466), .Q (new_AGEMA_signal_26467) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_26470), .Q (new_AGEMA_signal_26471) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_26474), .Q (new_AGEMA_signal_26475) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_26478), .Q (new_AGEMA_signal_26479) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_26482), .Q (new_AGEMA_signal_26483) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_26486), .Q (new_AGEMA_signal_26487) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_26490), .Q (new_AGEMA_signal_26491) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_26494), .Q (new_AGEMA_signal_26495) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_26498), .Q (new_AGEMA_signal_26499) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_26502), .Q (new_AGEMA_signal_26503) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_26506), .Q (new_AGEMA_signal_26507) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_26510), .Q (new_AGEMA_signal_26511) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_26514), .Q (new_AGEMA_signal_26515) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_26518), .Q (new_AGEMA_signal_26519) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_26522), .Q (new_AGEMA_signal_26523) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_26526), .Q (new_AGEMA_signal_26527) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_26530), .Q (new_AGEMA_signal_26531) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_26534), .Q (new_AGEMA_signal_26535) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_26538), .Q (new_AGEMA_signal_26539) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_26542), .Q (new_AGEMA_signal_26543) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_26546), .Q (new_AGEMA_signal_26547) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_26550), .Q (new_AGEMA_signal_26551) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_26554), .Q (new_AGEMA_signal_26555) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_26558), .Q (new_AGEMA_signal_26559) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_26562), .Q (new_AGEMA_signal_26563) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_26566), .Q (new_AGEMA_signal_26567) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_26570), .Q (new_AGEMA_signal_26571) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_26574), .Q (new_AGEMA_signal_26575) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_26578), .Q (new_AGEMA_signal_26579) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_26582), .Q (new_AGEMA_signal_26583) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_26586), .Q (new_AGEMA_signal_26587) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_26590), .Q (new_AGEMA_signal_26591) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_26594), .Q (new_AGEMA_signal_26595) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_26598), .Q (new_AGEMA_signal_26599) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_26602), .Q (new_AGEMA_signal_26603) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_26606), .Q (new_AGEMA_signal_26607) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_26610), .Q (new_AGEMA_signal_26611) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_26614), .Q (new_AGEMA_signal_26615) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_26618), .Q (new_AGEMA_signal_26619) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_26622), .Q (new_AGEMA_signal_26623) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_26626), .Q (new_AGEMA_signal_26627) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_26630), .Q (new_AGEMA_signal_26631) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_26634), .Q (new_AGEMA_signal_26635) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_26638), .Q (new_AGEMA_signal_26639) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_26642), .Q (new_AGEMA_signal_26643) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_26646), .Q (new_AGEMA_signal_26647) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_26650), .Q (new_AGEMA_signal_26651) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_26654), .Q (new_AGEMA_signal_26655) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_26658), .Q (new_AGEMA_signal_26659) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_26662), .Q (new_AGEMA_signal_26663) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_26666), .Q (new_AGEMA_signal_26667) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_26670), .Q (new_AGEMA_signal_26671) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_26674), .Q (new_AGEMA_signal_26675) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_26678), .Q (new_AGEMA_signal_26679) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_26682), .Q (new_AGEMA_signal_26683) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_26686), .Q (new_AGEMA_signal_26687) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_26690), .Q (new_AGEMA_signal_26691) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_26694), .Q (new_AGEMA_signal_26695) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_26698), .Q (new_AGEMA_signal_26699) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_26702), .Q (new_AGEMA_signal_26703) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_26706), .Q (new_AGEMA_signal_26707) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_26710), .Q (new_AGEMA_signal_26711) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_26714), .Q (new_AGEMA_signal_26715) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_26718), .Q (new_AGEMA_signal_26719) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_26722), .Q (new_AGEMA_signal_26723) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_26726), .Q (new_AGEMA_signal_26727) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_26730), .Q (new_AGEMA_signal_26731) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_26734), .Q (new_AGEMA_signal_26735) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_26738), .Q (new_AGEMA_signal_26739) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_26742), .Q (new_AGEMA_signal_26743) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_26746), .Q (new_AGEMA_signal_26747) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_26750), .Q (new_AGEMA_signal_26751) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_26754), .Q (new_AGEMA_signal_26755) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_26758), .Q (new_AGEMA_signal_26759) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_26762), .Q (new_AGEMA_signal_26763) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_26766), .Q (new_AGEMA_signal_26767) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_26770), .Q (new_AGEMA_signal_26771) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_26774), .Q (new_AGEMA_signal_26775) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_26778), .Q (new_AGEMA_signal_26779) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_26782), .Q (new_AGEMA_signal_26783) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_26786), .Q (new_AGEMA_signal_26787) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_26790), .Q (new_AGEMA_signal_26791) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_26794), .Q (new_AGEMA_signal_26795) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_26798), .Q (new_AGEMA_signal_26799) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_26802), .Q (new_AGEMA_signal_26803) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_26806), .Q (new_AGEMA_signal_26807) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_26810), .Q (new_AGEMA_signal_26811) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_26814), .Q (new_AGEMA_signal_26815) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_26818), .Q (new_AGEMA_signal_26819) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_26822), .Q (new_AGEMA_signal_26823) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_26826), .Q (new_AGEMA_signal_26827) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_26830), .Q (new_AGEMA_signal_26831) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_26834), .Q (new_AGEMA_signal_26835) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_26838), .Q (new_AGEMA_signal_26839) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_26842), .Q (new_AGEMA_signal_26843) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_26846), .Q (new_AGEMA_signal_26847) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_26850), .Q (new_AGEMA_signal_26851) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_26854), .Q (new_AGEMA_signal_26855) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_26858), .Q (new_AGEMA_signal_26859) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_26862), .Q (new_AGEMA_signal_26863) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_26866), .Q (new_AGEMA_signal_26867) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_26870), .Q (new_AGEMA_signal_26871) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_26874), .Q (new_AGEMA_signal_26875) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_26878), .Q (new_AGEMA_signal_26879) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_26882), .Q (new_AGEMA_signal_26883) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_26886), .Q (new_AGEMA_signal_26887) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_26890), .Q (new_AGEMA_signal_26891) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_26894), .Q (new_AGEMA_signal_26895) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_26898), .Q (new_AGEMA_signal_26899) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_26902), .Q (new_AGEMA_signal_26903) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_26906), .Q (new_AGEMA_signal_26907) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_26910), .Q (new_AGEMA_signal_26911) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_26914), .Q (new_AGEMA_signal_26915) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_26918), .Q (new_AGEMA_signal_26919) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_26922), .Q (new_AGEMA_signal_26923) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_26926), .Q (new_AGEMA_signal_26927) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_26930), .Q (new_AGEMA_signal_26931) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_26934), .Q (new_AGEMA_signal_26935) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_26938), .Q (new_AGEMA_signal_26939) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_26942), .Q (new_AGEMA_signal_26943) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_26946), .Q (new_AGEMA_signal_26947) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_26950), .Q (new_AGEMA_signal_26951) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_26954), .Q (new_AGEMA_signal_26955) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_26958), .Q (new_AGEMA_signal_26959) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_26962), .Q (new_AGEMA_signal_26963) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_26966), .Q (new_AGEMA_signal_26967) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_26970), .Q (new_AGEMA_signal_26971) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_26974), .Q (new_AGEMA_signal_26975) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_26978), .Q (new_AGEMA_signal_26979) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_26982), .Q (new_AGEMA_signal_26983) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_26986), .Q (new_AGEMA_signal_26987) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_26990), .Q (new_AGEMA_signal_26991) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_26994), .Q (new_AGEMA_signal_26995) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_26998), .Q (new_AGEMA_signal_26999) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_27002), .Q (new_AGEMA_signal_27003) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C (clk), .D (new_AGEMA_signal_27006), .Q (new_AGEMA_signal_27007) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_27010), .Q (new_AGEMA_signal_27011) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_27014), .Q (new_AGEMA_signal_27015) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C (clk), .D (new_AGEMA_signal_27018), .Q (new_AGEMA_signal_27019) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_27022), .Q (new_AGEMA_signal_27023) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_27026), .Q (new_AGEMA_signal_27027) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C (clk), .D (new_AGEMA_signal_27030), .Q (new_AGEMA_signal_27031) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_27034), .Q (new_AGEMA_signal_27035) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_27038), .Q (new_AGEMA_signal_27039) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C (clk), .D (new_AGEMA_signal_27042), .Q (new_AGEMA_signal_27043) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_27046), .Q (new_AGEMA_signal_27047) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_27050), .Q (new_AGEMA_signal_27051) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C (clk), .D (new_AGEMA_signal_27054), .Q (new_AGEMA_signal_27055) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_27058), .Q (new_AGEMA_signal_27059) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_27062), .Q (new_AGEMA_signal_27063) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C (clk), .D (new_AGEMA_signal_27066), .Q (new_AGEMA_signal_27067) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_27070), .Q (new_AGEMA_signal_27071) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_27074), .Q (new_AGEMA_signal_27075) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C (clk), .D (new_AGEMA_signal_27078), .Q (new_AGEMA_signal_27079) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_27082), .Q (new_AGEMA_signal_27083) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_27086), .Q (new_AGEMA_signal_27087) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C (clk), .D (new_AGEMA_signal_27090), .Q (new_AGEMA_signal_27091) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_27094), .Q (new_AGEMA_signal_27095) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_27098), .Q (new_AGEMA_signal_27099) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C (clk), .D (new_AGEMA_signal_27102), .Q (new_AGEMA_signal_27103) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_27106), .Q (new_AGEMA_signal_27107) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_27110), .Q (new_AGEMA_signal_27111) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C (clk), .D (new_AGEMA_signal_27114), .Q (new_AGEMA_signal_27115) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_27118), .Q (new_AGEMA_signal_27119) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_27122), .Q (new_AGEMA_signal_27123) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C (clk), .D (new_AGEMA_signal_27126), .Q (new_AGEMA_signal_27127) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_27130), .Q (new_AGEMA_signal_27131) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C (clk), .D (new_AGEMA_signal_27134), .Q (new_AGEMA_signal_27135) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C (clk), .D (new_AGEMA_signal_27138), .Q (new_AGEMA_signal_27139) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_27142), .Q (new_AGEMA_signal_27143) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_27146), .Q (new_AGEMA_signal_27147) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C (clk), .D (new_AGEMA_signal_27150), .Q (new_AGEMA_signal_27151) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_27154), .Q (new_AGEMA_signal_27155) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_27158), .Q (new_AGEMA_signal_27159) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C (clk), .D (new_AGEMA_signal_27162), .Q (new_AGEMA_signal_27163) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_27166), .Q (new_AGEMA_signal_27167) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C (clk), .D (new_AGEMA_signal_27170), .Q (new_AGEMA_signal_27171) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C (clk), .D (new_AGEMA_signal_27174), .Q (new_AGEMA_signal_27175) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_27178), .Q (new_AGEMA_signal_27179) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_27182), .Q (new_AGEMA_signal_27183) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C (clk), .D (new_AGEMA_signal_27186), .Q (new_AGEMA_signal_27187) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_27190), .Q (new_AGEMA_signal_27191) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_27194), .Q (new_AGEMA_signal_27195) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C (clk), .D (new_AGEMA_signal_27198), .Q (new_AGEMA_signal_27199) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_27202), .Q (new_AGEMA_signal_27203) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C (clk), .D (new_AGEMA_signal_27206), .Q (new_AGEMA_signal_27207) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C (clk), .D (new_AGEMA_signal_27210), .Q (new_AGEMA_signal_27211) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_27214), .Q (new_AGEMA_signal_27215) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_27218), .Q (new_AGEMA_signal_27219) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C (clk), .D (new_AGEMA_signal_27222), .Q (new_AGEMA_signal_27223) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_27226), .Q (new_AGEMA_signal_27227) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_27230), .Q (new_AGEMA_signal_27231) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C (clk), .D (new_AGEMA_signal_27234), .Q (new_AGEMA_signal_27235) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_27238), .Q (new_AGEMA_signal_27239) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C (clk), .D (new_AGEMA_signal_27242), .Q (new_AGEMA_signal_27243) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C (clk), .D (new_AGEMA_signal_27246), .Q (new_AGEMA_signal_27247) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_27250), .Q (new_AGEMA_signal_27251) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_27254), .Q (new_AGEMA_signal_27255) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C (clk), .D (new_AGEMA_signal_27258), .Q (new_AGEMA_signal_27259) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_27262), .Q (new_AGEMA_signal_27263) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_27266), .Q (new_AGEMA_signal_27267) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C (clk), .D (new_AGEMA_signal_27270), .Q (new_AGEMA_signal_27271) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_27274), .Q (new_AGEMA_signal_27275) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C (clk), .D (new_AGEMA_signal_27278), .Q (new_AGEMA_signal_27279) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C (clk), .D (new_AGEMA_signal_27282), .Q (new_AGEMA_signal_27283) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_27286), .Q (new_AGEMA_signal_27287) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_27290), .Q (new_AGEMA_signal_27291) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C (clk), .D (new_AGEMA_signal_27294), .Q (new_AGEMA_signal_27295) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_27298), .Q (new_AGEMA_signal_27299) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_27302), .Q (new_AGEMA_signal_27303) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C (clk), .D (new_AGEMA_signal_27306), .Q (new_AGEMA_signal_27307) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_27310), .Q (new_AGEMA_signal_27311) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C (clk), .D (new_AGEMA_signal_27314), .Q (new_AGEMA_signal_27315) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C (clk), .D (new_AGEMA_signal_27318), .Q (new_AGEMA_signal_27319) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_27322), .Q (new_AGEMA_signal_27323) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_27326), .Q (new_AGEMA_signal_27327) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C (clk), .D (new_AGEMA_signal_27330), .Q (new_AGEMA_signal_27331) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_27334), .Q (new_AGEMA_signal_27335) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_27338), .Q (new_AGEMA_signal_27339) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C (clk), .D (new_AGEMA_signal_27342), .Q (new_AGEMA_signal_27343) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_27346), .Q (new_AGEMA_signal_27347) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C (clk), .D (new_AGEMA_signal_27350), .Q (new_AGEMA_signal_27351) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C (clk), .D (new_AGEMA_signal_27354), .Q (new_AGEMA_signal_27355) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_27358), .Q (new_AGEMA_signal_27359) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_27362), .Q (new_AGEMA_signal_27363) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C (clk), .D (new_AGEMA_signal_27366), .Q (new_AGEMA_signal_27367) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_27370), .Q (new_AGEMA_signal_27371) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_27374), .Q (new_AGEMA_signal_27375) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C (clk), .D (new_AGEMA_signal_27378), .Q (new_AGEMA_signal_27379) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_27382), .Q (new_AGEMA_signal_27383) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C (clk), .D (new_AGEMA_signal_27386), .Q (new_AGEMA_signal_27387) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C (clk), .D (new_AGEMA_signal_27390), .Q (new_AGEMA_signal_27391) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_27394), .Q (new_AGEMA_signal_27395) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_27398), .Q (new_AGEMA_signal_27399) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C (clk), .D (new_AGEMA_signal_27402), .Q (new_AGEMA_signal_27403) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_27406), .Q (new_AGEMA_signal_27407) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_27410), .Q (new_AGEMA_signal_27411) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C (clk), .D (new_AGEMA_signal_27414), .Q (new_AGEMA_signal_27415) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C (clk), .D (new_AGEMA_signal_27418), .Q (new_AGEMA_signal_27419) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_27422), .Q (new_AGEMA_signal_27423) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C (clk), .D (new_AGEMA_signal_27426), .Q (new_AGEMA_signal_27427) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_27430), .Q (new_AGEMA_signal_27431) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C (clk), .D (new_AGEMA_signal_27434), .Q (new_AGEMA_signal_27435) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C (clk), .D (new_AGEMA_signal_27438), .Q (new_AGEMA_signal_27439) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C (clk), .D (new_AGEMA_signal_27442), .Q (new_AGEMA_signal_27443) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_27446), .Q (new_AGEMA_signal_27447) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C (clk), .D (new_AGEMA_signal_27450), .Q (new_AGEMA_signal_27451) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_27454), .Q (new_AGEMA_signal_27455) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_27458), .Q (new_AGEMA_signal_27459) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C (clk), .D (new_AGEMA_signal_27462), .Q (new_AGEMA_signal_27463) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_27466), .Q (new_AGEMA_signal_27467) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C (clk), .D (new_AGEMA_signal_27470), .Q (new_AGEMA_signal_27471) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C (clk), .D (new_AGEMA_signal_27474), .Q (new_AGEMA_signal_27475) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_27478), .Q (new_AGEMA_signal_27479) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_27482), .Q (new_AGEMA_signal_27483) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C (clk), .D (new_AGEMA_signal_27486), .Q (new_AGEMA_signal_27487) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_27490), .Q (new_AGEMA_signal_27491) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_27494), .Q (new_AGEMA_signal_27495) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C (clk), .D (new_AGEMA_signal_27498), .Q (new_AGEMA_signal_27499) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_27502), .Q (new_AGEMA_signal_27503) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C (clk), .D (new_AGEMA_signal_27506), .Q (new_AGEMA_signal_27507) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C (clk), .D (new_AGEMA_signal_27510), .Q (new_AGEMA_signal_27511) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_27514), .Q (new_AGEMA_signal_27515) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_27518), .Q (new_AGEMA_signal_27519) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C (clk), .D (new_AGEMA_signal_27522), .Q (new_AGEMA_signal_27523) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_27526), .Q (new_AGEMA_signal_27527) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_27530), .Q (new_AGEMA_signal_27531) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C (clk), .D (new_AGEMA_signal_27534), .Q (new_AGEMA_signal_27535) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_27538), .Q (new_AGEMA_signal_27539) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C (clk), .D (new_AGEMA_signal_27542), .Q (new_AGEMA_signal_27543) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C (clk), .D (new_AGEMA_signal_27546), .Q (new_AGEMA_signal_27547) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_27550), .Q (new_AGEMA_signal_27551) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_27554), .Q (new_AGEMA_signal_27555) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C (clk), .D (new_AGEMA_signal_27558), .Q (new_AGEMA_signal_27559) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_27562), .Q (new_AGEMA_signal_27563) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_27566), .Q (new_AGEMA_signal_27567) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C (clk), .D (new_AGEMA_signal_27570), .Q (new_AGEMA_signal_27571) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_27574), .Q (new_AGEMA_signal_27575) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C (clk), .D (new_AGEMA_signal_27578), .Q (new_AGEMA_signal_27579) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C (clk), .D (new_AGEMA_signal_27582), .Q (new_AGEMA_signal_27583) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_27586), .Q (new_AGEMA_signal_27587) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_27590), .Q (new_AGEMA_signal_27591) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C (clk), .D (new_AGEMA_signal_27594), .Q (new_AGEMA_signal_27595) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_27598), .Q (new_AGEMA_signal_27599) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_27602), .Q (new_AGEMA_signal_27603) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C (clk), .D (new_AGEMA_signal_27606), .Q (new_AGEMA_signal_27607) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_27610), .Q (new_AGEMA_signal_27611) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C (clk), .D (new_AGEMA_signal_27614), .Q (new_AGEMA_signal_27615) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C (clk), .D (new_AGEMA_signal_27618), .Q (new_AGEMA_signal_27619) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_27622), .Q (new_AGEMA_signal_27623) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_27626), .Q (new_AGEMA_signal_27627) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C (clk), .D (new_AGEMA_signal_27630), .Q (new_AGEMA_signal_27631) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_27634), .Q (new_AGEMA_signal_27635) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C (clk), .D (new_AGEMA_signal_27638), .Q (new_AGEMA_signal_27639) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C (clk), .D (new_AGEMA_signal_27642), .Q (new_AGEMA_signal_27643) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C (clk), .D (new_AGEMA_signal_27646), .Q (new_AGEMA_signal_27647) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C (clk), .D (new_AGEMA_signal_27650), .Q (new_AGEMA_signal_27651) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C (clk), .D (new_AGEMA_signal_27654), .Q (new_AGEMA_signal_27655) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C (clk), .D (new_AGEMA_signal_27658), .Q (new_AGEMA_signal_27659) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C (clk), .D (new_AGEMA_signal_27662), .Q (new_AGEMA_signal_27663) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C (clk), .D (new_AGEMA_signal_27666), .Q (new_AGEMA_signal_27667) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C (clk), .D (new_AGEMA_signal_27670), .Q (new_AGEMA_signal_27671) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C (clk), .D (new_AGEMA_signal_27674), .Q (new_AGEMA_signal_27675) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C (clk), .D (new_AGEMA_signal_27678), .Q (new_AGEMA_signal_27679) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C (clk), .D (new_AGEMA_signal_27682), .Q (new_AGEMA_signal_27683) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C (clk), .D (new_AGEMA_signal_27686), .Q (new_AGEMA_signal_27687) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C (clk), .D (new_AGEMA_signal_27690), .Q (new_AGEMA_signal_27691) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C (clk), .D (new_AGEMA_signal_27694), .Q (new_AGEMA_signal_27695) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C (clk), .D (new_AGEMA_signal_27698), .Q (new_AGEMA_signal_27699) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C (clk), .D (new_AGEMA_signal_27702), .Q (new_AGEMA_signal_27703) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C (clk), .D (new_AGEMA_signal_27706), .Q (new_AGEMA_signal_27707) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C (clk), .D (new_AGEMA_signal_27710), .Q (new_AGEMA_signal_27711) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C (clk), .D (new_AGEMA_signal_27714), .Q (new_AGEMA_signal_27715) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C (clk), .D (new_AGEMA_signal_27718), .Q (new_AGEMA_signal_27719) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C (clk), .D (new_AGEMA_signal_27722), .Q (new_AGEMA_signal_27723) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C (clk), .D (new_AGEMA_signal_27726), .Q (new_AGEMA_signal_27727) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C (clk), .D (new_AGEMA_signal_27730), .Q (new_AGEMA_signal_27731) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C (clk), .D (new_AGEMA_signal_27734), .Q (new_AGEMA_signal_27735) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C (clk), .D (new_AGEMA_signal_27738), .Q (new_AGEMA_signal_27739) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C (clk), .D (new_AGEMA_signal_27742), .Q (new_AGEMA_signal_27743) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C (clk), .D (new_AGEMA_signal_27746), .Q (new_AGEMA_signal_27747) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C (clk), .D (new_AGEMA_signal_27750), .Q (new_AGEMA_signal_27751) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C (clk), .D (new_AGEMA_signal_27754), .Q (new_AGEMA_signal_27755) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C (clk), .D (new_AGEMA_signal_27758), .Q (new_AGEMA_signal_27759) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C (clk), .D (new_AGEMA_signal_27762), .Q (new_AGEMA_signal_27763) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C (clk), .D (new_AGEMA_signal_27766), .Q (new_AGEMA_signal_27767) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C (clk), .D (new_AGEMA_signal_27770), .Q (new_AGEMA_signal_27771) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C (clk), .D (new_AGEMA_signal_27774), .Q (new_AGEMA_signal_27775) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C (clk), .D (new_AGEMA_signal_27778), .Q (new_AGEMA_signal_27779) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C (clk), .D (new_AGEMA_signal_27782), .Q (new_AGEMA_signal_27783) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C (clk), .D (new_AGEMA_signal_27786), .Q (new_AGEMA_signal_27787) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C (clk), .D (new_AGEMA_signal_27790), .Q (new_AGEMA_signal_27791) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C (clk), .D (new_AGEMA_signal_27794), .Q (new_AGEMA_signal_27795) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C (clk), .D (new_AGEMA_signal_27798), .Q (new_AGEMA_signal_27799) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C (clk), .D (new_AGEMA_signal_27802), .Q (new_AGEMA_signal_27803) ) ;
    buf_clk new_AGEMA_reg_buffer_6851 ( .C (clk), .D (new_AGEMA_signal_27806), .Q (new_AGEMA_signal_27807) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C (clk), .D (new_AGEMA_signal_27810), .Q (new_AGEMA_signal_27811) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C (clk), .D (new_AGEMA_signal_27814), .Q (new_AGEMA_signal_27815) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C (clk), .D (new_AGEMA_signal_27818), .Q (new_AGEMA_signal_27819) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C (clk), .D (new_AGEMA_signal_27822), .Q (new_AGEMA_signal_27823) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C (clk), .D (new_AGEMA_signal_27826), .Q (new_AGEMA_signal_27827) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C (clk), .D (new_AGEMA_signal_27830), .Q (new_AGEMA_signal_27831) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C (clk), .D (new_AGEMA_signal_27834), .Q (new_AGEMA_signal_27835) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C (clk), .D (new_AGEMA_signal_27838), .Q (new_AGEMA_signal_27839) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C (clk), .D (new_AGEMA_signal_27842), .Q (new_AGEMA_signal_27843) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C (clk), .D (new_AGEMA_signal_27846), .Q (new_AGEMA_signal_27847) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C (clk), .D (new_AGEMA_signal_27850), .Q (new_AGEMA_signal_27851) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C (clk), .D (new_AGEMA_signal_27854), .Q (new_AGEMA_signal_27855) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C (clk), .D (new_AGEMA_signal_27858), .Q (new_AGEMA_signal_27859) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C (clk), .D (new_AGEMA_signal_27862), .Q (new_AGEMA_signal_27863) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C (clk), .D (new_AGEMA_signal_27866), .Q (new_AGEMA_signal_27867) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C (clk), .D (new_AGEMA_signal_27870), .Q (new_AGEMA_signal_27871) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C (clk), .D (new_AGEMA_signal_27874), .Q (new_AGEMA_signal_27875) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C (clk), .D (new_AGEMA_signal_27878), .Q (new_AGEMA_signal_27879) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C (clk), .D (new_AGEMA_signal_27882), .Q (new_AGEMA_signal_27883) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C (clk), .D (new_AGEMA_signal_27886), .Q (new_AGEMA_signal_27887) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C (clk), .D (new_AGEMA_signal_27890), .Q (new_AGEMA_signal_27891) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C (clk), .D (new_AGEMA_signal_27894), .Q (new_AGEMA_signal_27895) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C (clk), .D (new_AGEMA_signal_27898), .Q (new_AGEMA_signal_27899) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C (clk), .D (new_AGEMA_signal_27902), .Q (new_AGEMA_signal_27903) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C (clk), .D (new_AGEMA_signal_27906), .Q (new_AGEMA_signal_27907) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C (clk), .D (new_AGEMA_signal_27910), .Q (new_AGEMA_signal_27911) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C (clk), .D (new_AGEMA_signal_27914), .Q (new_AGEMA_signal_27915) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C (clk), .D (new_AGEMA_signal_27918), .Q (new_AGEMA_signal_27919) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C (clk), .D (new_AGEMA_signal_27922), .Q (new_AGEMA_signal_27923) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C (clk), .D (new_AGEMA_signal_27926), .Q (new_AGEMA_signal_27927) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C (clk), .D (new_AGEMA_signal_27930), .Q (new_AGEMA_signal_27931) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C (clk), .D (new_AGEMA_signal_27934), .Q (new_AGEMA_signal_27935) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C (clk), .D (new_AGEMA_signal_27938), .Q (new_AGEMA_signal_27939) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C (clk), .D (new_AGEMA_signal_27942), .Q (new_AGEMA_signal_27943) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C (clk), .D (new_AGEMA_signal_27946), .Q (new_AGEMA_signal_27947) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C (clk), .D (new_AGEMA_signal_27950), .Q (new_AGEMA_signal_27951) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C (clk), .D (new_AGEMA_signal_27954), .Q (new_AGEMA_signal_27955) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C (clk), .D (new_AGEMA_signal_27958), .Q (new_AGEMA_signal_27959) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C (clk), .D (new_AGEMA_signal_27962), .Q (new_AGEMA_signal_27963) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C (clk), .D (new_AGEMA_signal_27966), .Q (new_AGEMA_signal_27967) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C (clk), .D (new_AGEMA_signal_27970), .Q (new_AGEMA_signal_27971) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C (clk), .D (new_AGEMA_signal_27974), .Q (new_AGEMA_signal_27975) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C (clk), .D (new_AGEMA_signal_27978), .Q (new_AGEMA_signal_27979) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C (clk), .D (new_AGEMA_signal_27982), .Q (new_AGEMA_signal_27983) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C (clk), .D (new_AGEMA_signal_27986), .Q (new_AGEMA_signal_27987) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C (clk), .D (new_AGEMA_signal_27990), .Q (new_AGEMA_signal_27991) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C (clk), .D (new_AGEMA_signal_27994), .Q (new_AGEMA_signal_27995) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C (clk), .D (new_AGEMA_signal_27998), .Q (new_AGEMA_signal_27999) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C (clk), .D (new_AGEMA_signal_28002), .Q (new_AGEMA_signal_28003) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C (clk), .D (new_AGEMA_signal_28006), .Q (new_AGEMA_signal_28007) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C (clk), .D (new_AGEMA_signal_28010), .Q (new_AGEMA_signal_28011) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C (clk), .D (new_AGEMA_signal_28014), .Q (new_AGEMA_signal_28015) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C (clk), .D (new_AGEMA_signal_28018), .Q (new_AGEMA_signal_28019) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C (clk), .D (new_AGEMA_signal_28022), .Q (new_AGEMA_signal_28023) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C (clk), .D (new_AGEMA_signal_28026), .Q (new_AGEMA_signal_28027) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C (clk), .D (new_AGEMA_signal_28030), .Q (new_AGEMA_signal_28031) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C (clk), .D (new_AGEMA_signal_28034), .Q (new_AGEMA_signal_28035) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C (clk), .D (new_AGEMA_signal_28038), .Q (new_AGEMA_signal_28039) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C (clk), .D (new_AGEMA_signal_28042), .Q (new_AGEMA_signal_28043) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C (clk), .D (new_AGEMA_signal_28046), .Q (new_AGEMA_signal_28047) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C (clk), .D (new_AGEMA_signal_28050), .Q (new_AGEMA_signal_28051) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C (clk), .D (new_AGEMA_signal_28054), .Q (new_AGEMA_signal_28055) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C (clk), .D (new_AGEMA_signal_28058), .Q (new_AGEMA_signal_28059) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C (clk), .D (new_AGEMA_signal_28062), .Q (new_AGEMA_signal_28063) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C (clk), .D (new_AGEMA_signal_28066), .Q (new_AGEMA_signal_28067) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C (clk), .D (new_AGEMA_signal_28070), .Q (new_AGEMA_signal_28071) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C (clk), .D (new_AGEMA_signal_28074), .Q (new_AGEMA_signal_28075) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C (clk), .D (new_AGEMA_signal_28078), .Q (new_AGEMA_signal_28079) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C (clk), .D (new_AGEMA_signal_28082), .Q (new_AGEMA_signal_28083) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C (clk), .D (new_AGEMA_signal_28086), .Q (new_AGEMA_signal_28087) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C (clk), .D (new_AGEMA_signal_28090), .Q (new_AGEMA_signal_28091) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C (clk), .D (new_AGEMA_signal_28094), .Q (new_AGEMA_signal_28095) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C (clk), .D (new_AGEMA_signal_28098), .Q (new_AGEMA_signal_28099) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C (clk), .D (new_AGEMA_signal_28102), .Q (new_AGEMA_signal_28103) ) ;
    buf_clk new_AGEMA_reg_buffer_7151 ( .C (clk), .D (new_AGEMA_signal_28106), .Q (new_AGEMA_signal_28107) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C (clk), .D (new_AGEMA_signal_28110), .Q (new_AGEMA_signal_28111) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C (clk), .D (new_AGEMA_signal_28114), .Q (new_AGEMA_signal_28115) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C (clk), .D (new_AGEMA_signal_28118), .Q (new_AGEMA_signal_28119) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C (clk), .D (new_AGEMA_signal_28122), .Q (new_AGEMA_signal_28123) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C (clk), .D (new_AGEMA_signal_28126), .Q (new_AGEMA_signal_28127) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C (clk), .D (new_AGEMA_signal_28130), .Q (new_AGEMA_signal_28131) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C (clk), .D (new_AGEMA_signal_28134), .Q (new_AGEMA_signal_28135) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C (clk), .D (new_AGEMA_signal_28138), .Q (new_AGEMA_signal_28139) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C (clk), .D (new_AGEMA_signal_28142), .Q (new_AGEMA_signal_28143) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C (clk), .D (new_AGEMA_signal_28146), .Q (new_AGEMA_signal_28147) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C (clk), .D (new_AGEMA_signal_28150), .Q (new_AGEMA_signal_28151) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C (clk), .D (new_AGEMA_signal_28154), .Q (new_AGEMA_signal_28155) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C (clk), .D (new_AGEMA_signal_28158), .Q (new_AGEMA_signal_28159) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C (clk), .D (new_AGEMA_signal_28162), .Q (new_AGEMA_signal_28163) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C (clk), .D (new_AGEMA_signal_28166), .Q (new_AGEMA_signal_28167) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C (clk), .D (new_AGEMA_signal_28170), .Q (new_AGEMA_signal_28171) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C (clk), .D (new_AGEMA_signal_28174), .Q (new_AGEMA_signal_28175) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C (clk), .D (new_AGEMA_signal_28178), .Q (new_AGEMA_signal_28179) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C (clk), .D (new_AGEMA_signal_28182), .Q (new_AGEMA_signal_28183) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C (clk), .D (new_AGEMA_signal_28186), .Q (new_AGEMA_signal_28187) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C (clk), .D (new_AGEMA_signal_28190), .Q (new_AGEMA_signal_28191) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C (clk), .D (new_AGEMA_signal_28194), .Q (new_AGEMA_signal_28195) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C (clk), .D (new_AGEMA_signal_28198), .Q (new_AGEMA_signal_28199) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C (clk), .D (new_AGEMA_signal_28202), .Q (new_AGEMA_signal_28203) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C (clk), .D (new_AGEMA_signal_28206), .Q (new_AGEMA_signal_28207) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C (clk), .D (new_AGEMA_signal_28209), .Q (new_AGEMA_signal_28210) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C (clk), .D (new_AGEMA_signal_28212), .Q (new_AGEMA_signal_28213) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C (clk), .D (new_AGEMA_signal_28215), .Q (new_AGEMA_signal_28216) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C (clk), .D (new_AGEMA_signal_28218), .Q (new_AGEMA_signal_28219) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C (clk), .D (new_AGEMA_signal_28221), .Q (new_AGEMA_signal_28222) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C (clk), .D (new_AGEMA_signal_28224), .Q (new_AGEMA_signal_28225) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C (clk), .D (new_AGEMA_signal_28227), .Q (new_AGEMA_signal_28228) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C (clk), .D (new_AGEMA_signal_28230), .Q (new_AGEMA_signal_28231) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C (clk), .D (new_AGEMA_signal_28233), .Q (new_AGEMA_signal_28234) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C (clk), .D (new_AGEMA_signal_28236), .Q (new_AGEMA_signal_28237) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C (clk), .D (new_AGEMA_signal_28239), .Q (new_AGEMA_signal_28240) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C (clk), .D (new_AGEMA_signal_28242), .Q (new_AGEMA_signal_28243) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C (clk), .D (new_AGEMA_signal_28245), .Q (new_AGEMA_signal_28246) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C (clk), .D (new_AGEMA_signal_28248), .Q (new_AGEMA_signal_28249) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C (clk), .D (new_AGEMA_signal_28251), .Q (new_AGEMA_signal_28252) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C (clk), .D (new_AGEMA_signal_28254), .Q (new_AGEMA_signal_28255) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C (clk), .D (new_AGEMA_signal_28257), .Q (new_AGEMA_signal_28258) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C (clk), .D (new_AGEMA_signal_28260), .Q (new_AGEMA_signal_28261) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C (clk), .D (new_AGEMA_signal_28263), .Q (new_AGEMA_signal_28264) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C (clk), .D (new_AGEMA_signal_28266), .Q (new_AGEMA_signal_28267) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C (clk), .D (new_AGEMA_signal_28269), .Q (new_AGEMA_signal_28270) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C (clk), .D (new_AGEMA_signal_28272), .Q (new_AGEMA_signal_28273) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C (clk), .D (new_AGEMA_signal_28275), .Q (new_AGEMA_signal_28276) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C (clk), .D (new_AGEMA_signal_28278), .Q (new_AGEMA_signal_28279) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C (clk), .D (new_AGEMA_signal_28281), .Q (new_AGEMA_signal_28282) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C (clk), .D (new_AGEMA_signal_28284), .Q (new_AGEMA_signal_28285) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C (clk), .D (new_AGEMA_signal_28287), .Q (new_AGEMA_signal_28288) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C (clk), .D (new_AGEMA_signal_28290), .Q (new_AGEMA_signal_28291) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C (clk), .D (new_AGEMA_signal_28293), .Q (new_AGEMA_signal_28294) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C (clk), .D (new_AGEMA_signal_28296), .Q (new_AGEMA_signal_28297) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C (clk), .D (new_AGEMA_signal_28299), .Q (new_AGEMA_signal_28300) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C (clk), .D (new_AGEMA_signal_28302), .Q (new_AGEMA_signal_28303) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C (clk), .D (new_AGEMA_signal_28305), .Q (new_AGEMA_signal_28306) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C (clk), .D (new_AGEMA_signal_28308), .Q (new_AGEMA_signal_28309) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C (clk), .D (new_AGEMA_signal_28311), .Q (new_AGEMA_signal_28312) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C (clk), .D (new_AGEMA_signal_28314), .Q (new_AGEMA_signal_28315) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C (clk), .D (new_AGEMA_signal_28317), .Q (new_AGEMA_signal_28318) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C (clk), .D (new_AGEMA_signal_28320), .Q (new_AGEMA_signal_28321) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C (clk), .D (new_AGEMA_signal_28323), .Q (new_AGEMA_signal_28324) ) ;
    buf_clk new_AGEMA_reg_buffer_7371 ( .C (clk), .D (new_AGEMA_signal_28326), .Q (new_AGEMA_signal_28327) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C (clk), .D (new_AGEMA_signal_28329), .Q (new_AGEMA_signal_28330) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C (clk), .D (new_AGEMA_signal_28332), .Q (new_AGEMA_signal_28333) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C (clk), .D (new_AGEMA_signal_28335), .Q (new_AGEMA_signal_28336) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C (clk), .D (new_AGEMA_signal_28338), .Q (new_AGEMA_signal_28339) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C (clk), .D (new_AGEMA_signal_28341), .Q (new_AGEMA_signal_28342) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C (clk), .D (new_AGEMA_signal_28344), .Q (new_AGEMA_signal_28345) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C (clk), .D (new_AGEMA_signal_28347), .Q (new_AGEMA_signal_28348) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C (clk), .D (new_AGEMA_signal_28350), .Q (new_AGEMA_signal_28351) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C (clk), .D (new_AGEMA_signal_28353), .Q (new_AGEMA_signal_28354) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C (clk), .D (new_AGEMA_signal_28356), .Q (new_AGEMA_signal_28357) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C (clk), .D (new_AGEMA_signal_28359), .Q (new_AGEMA_signal_28360) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C (clk), .D (new_AGEMA_signal_28362), .Q (new_AGEMA_signal_28363) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C (clk), .D (new_AGEMA_signal_28365), .Q (new_AGEMA_signal_28366) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C (clk), .D (new_AGEMA_signal_28368), .Q (new_AGEMA_signal_28369) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C (clk), .D (new_AGEMA_signal_28371), .Q (new_AGEMA_signal_28372) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C (clk), .D (new_AGEMA_signal_28374), .Q (new_AGEMA_signal_28375) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C (clk), .D (new_AGEMA_signal_28377), .Q (new_AGEMA_signal_28378) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C (clk), .D (new_AGEMA_signal_28380), .Q (new_AGEMA_signal_28381) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C (clk), .D (new_AGEMA_signal_28383), .Q (new_AGEMA_signal_28384) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C (clk), .D (new_AGEMA_signal_28386), .Q (new_AGEMA_signal_28387) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C (clk), .D (new_AGEMA_signal_28389), .Q (new_AGEMA_signal_28390) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C (clk), .D (new_AGEMA_signal_28392), .Q (new_AGEMA_signal_28393) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C (clk), .D (new_AGEMA_signal_28395), .Q (new_AGEMA_signal_28396) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C (clk), .D (new_AGEMA_signal_28398), .Q (new_AGEMA_signal_28399) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C (clk), .D (new_AGEMA_signal_28401), .Q (new_AGEMA_signal_28402) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C (clk), .D (new_AGEMA_signal_28404), .Q (new_AGEMA_signal_28405) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C (clk), .D (new_AGEMA_signal_28407), .Q (new_AGEMA_signal_28408) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C (clk), .D (new_AGEMA_signal_28410), .Q (new_AGEMA_signal_28411) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C (clk), .D (new_AGEMA_signal_28413), .Q (new_AGEMA_signal_28414) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C (clk), .D (new_AGEMA_signal_28416), .Q (new_AGEMA_signal_28417) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C (clk), .D (new_AGEMA_signal_28419), .Q (new_AGEMA_signal_28420) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C (clk), .D (new_AGEMA_signal_28422), .Q (new_AGEMA_signal_28423) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C (clk), .D (new_AGEMA_signal_28425), .Q (new_AGEMA_signal_28426) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C (clk), .D (new_AGEMA_signal_28428), .Q (new_AGEMA_signal_28429) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C (clk), .D (new_AGEMA_signal_28431), .Q (new_AGEMA_signal_28432) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C (clk), .D (new_AGEMA_signal_28434), .Q (new_AGEMA_signal_28435) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C (clk), .D (new_AGEMA_signal_28437), .Q (new_AGEMA_signal_28438) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C (clk), .D (new_AGEMA_signal_28440), .Q (new_AGEMA_signal_28441) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C (clk), .D (new_AGEMA_signal_28443), .Q (new_AGEMA_signal_28444) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C (clk), .D (new_AGEMA_signal_28446), .Q (new_AGEMA_signal_28447) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C (clk), .D (new_AGEMA_signal_28449), .Q (new_AGEMA_signal_28450) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C (clk), .D (new_AGEMA_signal_28452), .Q (new_AGEMA_signal_28453) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C (clk), .D (new_AGEMA_signal_28455), .Q (new_AGEMA_signal_28456) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C (clk), .D (new_AGEMA_signal_28458), .Q (new_AGEMA_signal_28459) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C (clk), .D (new_AGEMA_signal_28461), .Q (new_AGEMA_signal_28462) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C (clk), .D (new_AGEMA_signal_28464), .Q (new_AGEMA_signal_28465) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C (clk), .D (new_AGEMA_signal_28467), .Q (new_AGEMA_signal_28468) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C (clk), .D (new_AGEMA_signal_28470), .Q (new_AGEMA_signal_28471) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C (clk), .D (new_AGEMA_signal_28473), .Q (new_AGEMA_signal_28474) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C (clk), .D (new_AGEMA_signal_28476), .Q (new_AGEMA_signal_28477) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C (clk), .D (new_AGEMA_signal_28479), .Q (new_AGEMA_signal_28480) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C (clk), .D (new_AGEMA_signal_28482), .Q (new_AGEMA_signal_28483) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C (clk), .D (new_AGEMA_signal_28485), .Q (new_AGEMA_signal_28486) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C (clk), .D (new_AGEMA_signal_28488), .Q (new_AGEMA_signal_28489) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C (clk), .D (new_AGEMA_signal_28491), .Q (new_AGEMA_signal_28492) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C (clk), .D (new_AGEMA_signal_28494), .Q (new_AGEMA_signal_28495) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C (clk), .D (new_AGEMA_signal_28497), .Q (new_AGEMA_signal_28498) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C (clk), .D (new_AGEMA_signal_28500), .Q (new_AGEMA_signal_28501) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C (clk), .D (new_AGEMA_signal_28503), .Q (new_AGEMA_signal_28504) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C (clk), .D (new_AGEMA_signal_28506), .Q (new_AGEMA_signal_28507) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C (clk), .D (new_AGEMA_signal_28509), .Q (new_AGEMA_signal_28510) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C (clk), .D (new_AGEMA_signal_28512), .Q (new_AGEMA_signal_28513) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C (clk), .D (new_AGEMA_signal_28515), .Q (new_AGEMA_signal_28516) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C (clk), .D (new_AGEMA_signal_28518), .Q (new_AGEMA_signal_28519) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C (clk), .D (new_AGEMA_signal_28521), .Q (new_AGEMA_signal_28522) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C (clk), .D (new_AGEMA_signal_28524), .Q (new_AGEMA_signal_28525) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C (clk), .D (new_AGEMA_signal_28527), .Q (new_AGEMA_signal_28528) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C (clk), .D (new_AGEMA_signal_28530), .Q (new_AGEMA_signal_28531) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C (clk), .D (new_AGEMA_signal_28533), .Q (new_AGEMA_signal_28534) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C (clk), .D (new_AGEMA_signal_28536), .Q (new_AGEMA_signal_28537) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C (clk), .D (new_AGEMA_signal_28539), .Q (new_AGEMA_signal_28540) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C (clk), .D (new_AGEMA_signal_28542), .Q (new_AGEMA_signal_28543) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C (clk), .D (new_AGEMA_signal_28545), .Q (new_AGEMA_signal_28546) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C (clk), .D (new_AGEMA_signal_28548), .Q (new_AGEMA_signal_28549) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C (clk), .D (new_AGEMA_signal_28551), .Q (new_AGEMA_signal_28552) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C (clk), .D (new_AGEMA_signal_28554), .Q (new_AGEMA_signal_28555) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C (clk), .D (new_AGEMA_signal_28557), .Q (new_AGEMA_signal_28558) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C (clk), .D (new_AGEMA_signal_28560), .Q (new_AGEMA_signal_28561) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C (clk), .D (new_AGEMA_signal_28563), .Q (new_AGEMA_signal_28564) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C (clk), .D (new_AGEMA_signal_28566), .Q (new_AGEMA_signal_28567) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C (clk), .D (new_AGEMA_signal_28569), .Q (new_AGEMA_signal_28570) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C (clk), .D (new_AGEMA_signal_28572), .Q (new_AGEMA_signal_28573) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C (clk), .D (new_AGEMA_signal_28575), .Q (new_AGEMA_signal_28576) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C (clk), .D (new_AGEMA_signal_28578), .Q (new_AGEMA_signal_28579) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C (clk), .D (new_AGEMA_signal_28581), .Q (new_AGEMA_signal_28582) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C (clk), .D (new_AGEMA_signal_28584), .Q (new_AGEMA_signal_28585) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C (clk), .D (new_AGEMA_signal_28587), .Q (new_AGEMA_signal_28588) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C (clk), .D (new_AGEMA_signal_28590), .Q (new_AGEMA_signal_28591) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C (clk), .D (new_AGEMA_signal_28593), .Q (new_AGEMA_signal_28594) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C (clk), .D (new_AGEMA_signal_28596), .Q (new_AGEMA_signal_28597) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C (clk), .D (new_AGEMA_signal_28599), .Q (new_AGEMA_signal_28600) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C (clk), .D (new_AGEMA_signal_28602), .Q (new_AGEMA_signal_28603) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C (clk), .D (new_AGEMA_signal_28605), .Q (new_AGEMA_signal_28606) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C (clk), .D (new_AGEMA_signal_28608), .Q (new_AGEMA_signal_28609) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C (clk), .D (new_AGEMA_signal_28611), .Q (new_AGEMA_signal_28612) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C (clk), .D (new_AGEMA_signal_28614), .Q (new_AGEMA_signal_28615) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C (clk), .D (new_AGEMA_signal_28617), .Q (new_AGEMA_signal_28618) ) ;
    buf_clk new_AGEMA_reg_buffer_7665 ( .C (clk), .D (new_AGEMA_signal_28620), .Q (new_AGEMA_signal_28621) ) ;
    buf_clk new_AGEMA_reg_buffer_7668 ( .C (clk), .D (new_AGEMA_signal_28623), .Q (new_AGEMA_signal_28624) ) ;
    buf_clk new_AGEMA_reg_buffer_7671 ( .C (clk), .D (new_AGEMA_signal_28626), .Q (new_AGEMA_signal_28627) ) ;
    buf_clk new_AGEMA_reg_buffer_7674 ( .C (clk), .D (new_AGEMA_signal_28629), .Q (new_AGEMA_signal_28630) ) ;
    buf_clk new_AGEMA_reg_buffer_7677 ( .C (clk), .D (new_AGEMA_signal_28632), .Q (new_AGEMA_signal_28633) ) ;
    buf_clk new_AGEMA_reg_buffer_7680 ( .C (clk), .D (new_AGEMA_signal_28635), .Q (new_AGEMA_signal_28636) ) ;
    buf_clk new_AGEMA_reg_buffer_7683 ( .C (clk), .D (new_AGEMA_signal_28638), .Q (new_AGEMA_signal_28639) ) ;
    buf_clk new_AGEMA_reg_buffer_7686 ( .C (clk), .D (new_AGEMA_signal_28641), .Q (new_AGEMA_signal_28642) ) ;
    buf_clk new_AGEMA_reg_buffer_7689 ( .C (clk), .D (new_AGEMA_signal_28644), .Q (new_AGEMA_signal_28645) ) ;
    buf_clk new_AGEMA_reg_buffer_7692 ( .C (clk), .D (new_AGEMA_signal_28647), .Q (new_AGEMA_signal_28648) ) ;
    buf_clk new_AGEMA_reg_buffer_7695 ( .C (clk), .D (new_AGEMA_signal_28650), .Q (new_AGEMA_signal_28651) ) ;
    buf_clk new_AGEMA_reg_buffer_7698 ( .C (clk), .D (new_AGEMA_signal_28653), .Q (new_AGEMA_signal_28654) ) ;
    buf_clk new_AGEMA_reg_buffer_7701 ( .C (clk), .D (new_AGEMA_signal_28656), .Q (new_AGEMA_signal_28657) ) ;
    buf_clk new_AGEMA_reg_buffer_7704 ( .C (clk), .D (new_AGEMA_signal_28659), .Q (new_AGEMA_signal_28660) ) ;
    buf_clk new_AGEMA_reg_buffer_7707 ( .C (clk), .D (new_AGEMA_signal_28662), .Q (new_AGEMA_signal_28663) ) ;
    buf_clk new_AGEMA_reg_buffer_7710 ( .C (clk), .D (new_AGEMA_signal_28665), .Q (new_AGEMA_signal_28666) ) ;
    buf_clk new_AGEMA_reg_buffer_7713 ( .C (clk), .D (new_AGEMA_signal_28668), .Q (new_AGEMA_signal_28669) ) ;
    buf_clk new_AGEMA_reg_buffer_7716 ( .C (clk), .D (new_AGEMA_signal_28671), .Q (new_AGEMA_signal_28672) ) ;
    buf_clk new_AGEMA_reg_buffer_7719 ( .C (clk), .D (new_AGEMA_signal_28674), .Q (new_AGEMA_signal_28675) ) ;
    buf_clk new_AGEMA_reg_buffer_7722 ( .C (clk), .D (new_AGEMA_signal_28677), .Q (new_AGEMA_signal_28678) ) ;
    buf_clk new_AGEMA_reg_buffer_7725 ( .C (clk), .D (new_AGEMA_signal_28680), .Q (new_AGEMA_signal_28681) ) ;
    buf_clk new_AGEMA_reg_buffer_7728 ( .C (clk), .D (new_AGEMA_signal_28683), .Q (new_AGEMA_signal_28684) ) ;
    buf_clk new_AGEMA_reg_buffer_7731 ( .C (clk), .D (new_AGEMA_signal_28686), .Q (new_AGEMA_signal_28687) ) ;
    buf_clk new_AGEMA_reg_buffer_7734 ( .C (clk), .D (new_AGEMA_signal_28689), .Q (new_AGEMA_signal_28690) ) ;
    buf_clk new_AGEMA_reg_buffer_7737 ( .C (clk), .D (new_AGEMA_signal_28692), .Q (new_AGEMA_signal_28693) ) ;
    buf_clk new_AGEMA_reg_buffer_7740 ( .C (clk), .D (new_AGEMA_signal_28695), .Q (new_AGEMA_signal_28696) ) ;
    buf_clk new_AGEMA_reg_buffer_7743 ( .C (clk), .D (new_AGEMA_signal_28698), .Q (new_AGEMA_signal_28699) ) ;
    buf_clk new_AGEMA_reg_buffer_7746 ( .C (clk), .D (new_AGEMA_signal_28701), .Q (new_AGEMA_signal_28702) ) ;
    buf_clk new_AGEMA_reg_buffer_7749 ( .C (clk), .D (new_AGEMA_signal_28704), .Q (new_AGEMA_signal_28705) ) ;
    buf_clk new_AGEMA_reg_buffer_7752 ( .C (clk), .D (new_AGEMA_signal_28707), .Q (new_AGEMA_signal_28708) ) ;
    buf_clk new_AGEMA_reg_buffer_7755 ( .C (clk), .D (new_AGEMA_signal_28710), .Q (new_AGEMA_signal_28711) ) ;
    buf_clk new_AGEMA_reg_buffer_7758 ( .C (clk), .D (new_AGEMA_signal_28713), .Q (new_AGEMA_signal_28714) ) ;
    buf_clk new_AGEMA_reg_buffer_7761 ( .C (clk), .D (new_AGEMA_signal_28716), .Q (new_AGEMA_signal_28717) ) ;
    buf_clk new_AGEMA_reg_buffer_7764 ( .C (clk), .D (new_AGEMA_signal_28719), .Q (new_AGEMA_signal_28720) ) ;
    buf_clk new_AGEMA_reg_buffer_7767 ( .C (clk), .D (new_AGEMA_signal_28722), .Q (new_AGEMA_signal_28723) ) ;
    buf_clk new_AGEMA_reg_buffer_7770 ( .C (clk), .D (new_AGEMA_signal_28725), .Q (new_AGEMA_signal_28726) ) ;
    buf_clk new_AGEMA_reg_buffer_7773 ( .C (clk), .D (new_AGEMA_signal_28728), .Q (new_AGEMA_signal_28729) ) ;
    buf_clk new_AGEMA_reg_buffer_7776 ( .C (clk), .D (new_AGEMA_signal_28731), .Q (new_AGEMA_signal_28732) ) ;
    buf_clk new_AGEMA_reg_buffer_7779 ( .C (clk), .D (new_AGEMA_signal_28734), .Q (new_AGEMA_signal_28735) ) ;
    buf_clk new_AGEMA_reg_buffer_7782 ( .C (clk), .D (new_AGEMA_signal_28737), .Q (new_AGEMA_signal_28738) ) ;
    buf_clk new_AGEMA_reg_buffer_7785 ( .C (clk), .D (new_AGEMA_signal_28740), .Q (new_AGEMA_signal_28741) ) ;
    buf_clk new_AGEMA_reg_buffer_7788 ( .C (clk), .D (new_AGEMA_signal_28743), .Q (new_AGEMA_signal_28744) ) ;
    buf_clk new_AGEMA_reg_buffer_7791 ( .C (clk), .D (new_AGEMA_signal_28746), .Q (new_AGEMA_signal_28747) ) ;
    buf_clk new_AGEMA_reg_buffer_7794 ( .C (clk), .D (new_AGEMA_signal_28749), .Q (new_AGEMA_signal_28750) ) ;
    buf_clk new_AGEMA_reg_buffer_7797 ( .C (clk), .D (new_AGEMA_signal_28752), .Q (new_AGEMA_signal_28753) ) ;
    buf_clk new_AGEMA_reg_buffer_7800 ( .C (clk), .D (new_AGEMA_signal_28755), .Q (new_AGEMA_signal_28756) ) ;
    buf_clk new_AGEMA_reg_buffer_7803 ( .C (clk), .D (new_AGEMA_signal_28758), .Q (new_AGEMA_signal_28759) ) ;
    buf_clk new_AGEMA_reg_buffer_7806 ( .C (clk), .D (new_AGEMA_signal_28761), .Q (new_AGEMA_signal_28762) ) ;
    buf_clk new_AGEMA_reg_buffer_7809 ( .C (clk), .D (new_AGEMA_signal_28764), .Q (new_AGEMA_signal_28765) ) ;
    buf_clk new_AGEMA_reg_buffer_7812 ( .C (clk), .D (new_AGEMA_signal_28767), .Q (new_AGEMA_signal_28768) ) ;
    buf_clk new_AGEMA_reg_buffer_7815 ( .C (clk), .D (new_AGEMA_signal_28770), .Q (new_AGEMA_signal_28771) ) ;
    buf_clk new_AGEMA_reg_buffer_7818 ( .C (clk), .D (new_AGEMA_signal_28773), .Q (new_AGEMA_signal_28774) ) ;
    buf_clk new_AGEMA_reg_buffer_7821 ( .C (clk), .D (new_AGEMA_signal_28776), .Q (new_AGEMA_signal_28777) ) ;
    buf_clk new_AGEMA_reg_buffer_7824 ( .C (clk), .D (new_AGEMA_signal_28779), .Q (new_AGEMA_signal_28780) ) ;
    buf_clk new_AGEMA_reg_buffer_7827 ( .C (clk), .D (new_AGEMA_signal_28782), .Q (new_AGEMA_signal_28783) ) ;
    buf_clk new_AGEMA_reg_buffer_7830 ( .C (clk), .D (new_AGEMA_signal_28785), .Q (new_AGEMA_signal_28786) ) ;
    buf_clk new_AGEMA_reg_buffer_7833 ( .C (clk), .D (new_AGEMA_signal_28788), .Q (new_AGEMA_signal_28789) ) ;
    buf_clk new_AGEMA_reg_buffer_7836 ( .C (clk), .D (new_AGEMA_signal_28791), .Q (new_AGEMA_signal_28792) ) ;
    buf_clk new_AGEMA_reg_buffer_7839 ( .C (clk), .D (new_AGEMA_signal_28794), .Q (new_AGEMA_signal_28795) ) ;
    buf_clk new_AGEMA_reg_buffer_7842 ( .C (clk), .D (new_AGEMA_signal_28797), .Q (new_AGEMA_signal_28798) ) ;
    buf_clk new_AGEMA_reg_buffer_7845 ( .C (clk), .D (new_AGEMA_signal_28800), .Q (new_AGEMA_signal_28801) ) ;
    buf_clk new_AGEMA_reg_buffer_7848 ( .C (clk), .D (new_AGEMA_signal_28803), .Q (new_AGEMA_signal_28804) ) ;
    buf_clk new_AGEMA_reg_buffer_7851 ( .C (clk), .D (new_AGEMA_signal_28806), .Q (new_AGEMA_signal_28807) ) ;
    buf_clk new_AGEMA_reg_buffer_7854 ( .C (clk), .D (new_AGEMA_signal_28809), .Q (new_AGEMA_signal_28810) ) ;
    buf_clk new_AGEMA_reg_buffer_7857 ( .C (clk), .D (new_AGEMA_signal_28812), .Q (new_AGEMA_signal_28813) ) ;
    buf_clk new_AGEMA_reg_buffer_7860 ( .C (clk), .D (new_AGEMA_signal_28815), .Q (new_AGEMA_signal_28816) ) ;
    buf_clk new_AGEMA_reg_buffer_7863 ( .C (clk), .D (new_AGEMA_signal_28818), .Q (new_AGEMA_signal_28819) ) ;
    buf_clk new_AGEMA_reg_buffer_7866 ( .C (clk), .D (new_AGEMA_signal_28821), .Q (new_AGEMA_signal_28822) ) ;
    buf_clk new_AGEMA_reg_buffer_7869 ( .C (clk), .D (new_AGEMA_signal_28824), .Q (new_AGEMA_signal_28825) ) ;
    buf_clk new_AGEMA_reg_buffer_7872 ( .C (clk), .D (new_AGEMA_signal_28827), .Q (new_AGEMA_signal_28828) ) ;
    buf_clk new_AGEMA_reg_buffer_7875 ( .C (clk), .D (new_AGEMA_signal_28830), .Q (new_AGEMA_signal_28831) ) ;
    buf_clk new_AGEMA_reg_buffer_7878 ( .C (clk), .D (new_AGEMA_signal_28833), .Q (new_AGEMA_signal_28834) ) ;
    buf_clk new_AGEMA_reg_buffer_7881 ( .C (clk), .D (new_AGEMA_signal_28836), .Q (new_AGEMA_signal_28837) ) ;
    buf_clk new_AGEMA_reg_buffer_7884 ( .C (clk), .D (new_AGEMA_signal_28839), .Q (new_AGEMA_signal_28840) ) ;
    buf_clk new_AGEMA_reg_buffer_7887 ( .C (clk), .D (new_AGEMA_signal_28842), .Q (new_AGEMA_signal_28843) ) ;
    buf_clk new_AGEMA_reg_buffer_7890 ( .C (clk), .D (new_AGEMA_signal_28845), .Q (new_AGEMA_signal_28846) ) ;
    buf_clk new_AGEMA_reg_buffer_7893 ( .C (clk), .D (new_AGEMA_signal_28848), .Q (new_AGEMA_signal_28849) ) ;
    buf_clk new_AGEMA_reg_buffer_7896 ( .C (clk), .D (new_AGEMA_signal_28851), .Q (new_AGEMA_signal_28852) ) ;
    buf_clk new_AGEMA_reg_buffer_7899 ( .C (clk), .D (new_AGEMA_signal_28854), .Q (new_AGEMA_signal_28855) ) ;
    buf_clk new_AGEMA_reg_buffer_7902 ( .C (clk), .D (new_AGEMA_signal_28857), .Q (new_AGEMA_signal_28858) ) ;
    buf_clk new_AGEMA_reg_buffer_7905 ( .C (clk), .D (new_AGEMA_signal_28860), .Q (new_AGEMA_signal_28861) ) ;
    buf_clk new_AGEMA_reg_buffer_7908 ( .C (clk), .D (new_AGEMA_signal_28863), .Q (new_AGEMA_signal_28864) ) ;
    buf_clk new_AGEMA_reg_buffer_7911 ( .C (clk), .D (new_AGEMA_signal_28866), .Q (new_AGEMA_signal_28867) ) ;
    buf_clk new_AGEMA_reg_buffer_7914 ( .C (clk), .D (new_AGEMA_signal_28869), .Q (new_AGEMA_signal_28870) ) ;
    buf_clk new_AGEMA_reg_buffer_7917 ( .C (clk), .D (new_AGEMA_signal_28872), .Q (new_AGEMA_signal_28873) ) ;
    buf_clk new_AGEMA_reg_buffer_7920 ( .C (clk), .D (new_AGEMA_signal_28875), .Q (new_AGEMA_signal_28876) ) ;
    buf_clk new_AGEMA_reg_buffer_7923 ( .C (clk), .D (new_AGEMA_signal_28878), .Q (new_AGEMA_signal_28879) ) ;
    buf_clk new_AGEMA_reg_buffer_7926 ( .C (clk), .D (new_AGEMA_signal_28881), .Q (new_AGEMA_signal_28882) ) ;
    buf_clk new_AGEMA_reg_buffer_7929 ( .C (clk), .D (new_AGEMA_signal_28884), .Q (new_AGEMA_signal_28885) ) ;
    buf_clk new_AGEMA_reg_buffer_7932 ( .C (clk), .D (new_AGEMA_signal_28887), .Q (new_AGEMA_signal_28888) ) ;
    buf_clk new_AGEMA_reg_buffer_7935 ( .C (clk), .D (new_AGEMA_signal_28890), .Q (new_AGEMA_signal_28891) ) ;
    buf_clk new_AGEMA_reg_buffer_7938 ( .C (clk), .D (new_AGEMA_signal_28893), .Q (new_AGEMA_signal_28894) ) ;
    buf_clk new_AGEMA_reg_buffer_7941 ( .C (clk), .D (new_AGEMA_signal_28896), .Q (new_AGEMA_signal_28897) ) ;
    buf_clk new_AGEMA_reg_buffer_7944 ( .C (clk), .D (new_AGEMA_signal_28899), .Q (new_AGEMA_signal_28900) ) ;
    buf_clk new_AGEMA_reg_buffer_7947 ( .C (clk), .D (new_AGEMA_signal_28902), .Q (new_AGEMA_signal_28903) ) ;
    buf_clk new_AGEMA_reg_buffer_7950 ( .C (clk), .D (new_AGEMA_signal_28905), .Q (new_AGEMA_signal_28906) ) ;
    buf_clk new_AGEMA_reg_buffer_7953 ( .C (clk), .D (new_AGEMA_signal_28908), .Q (new_AGEMA_signal_28909) ) ;
    buf_clk new_AGEMA_reg_buffer_7956 ( .C (clk), .D (new_AGEMA_signal_28911), .Q (new_AGEMA_signal_28912) ) ;
    buf_clk new_AGEMA_reg_buffer_7959 ( .C (clk), .D (new_AGEMA_signal_28914), .Q (new_AGEMA_signal_28915) ) ;
    buf_clk new_AGEMA_reg_buffer_7962 ( .C (clk), .D (new_AGEMA_signal_28917), .Q (new_AGEMA_signal_28918) ) ;
    buf_clk new_AGEMA_reg_buffer_7965 ( .C (clk), .D (new_AGEMA_signal_28920), .Q (new_AGEMA_signal_28921) ) ;
    buf_clk new_AGEMA_reg_buffer_7968 ( .C (clk), .D (new_AGEMA_signal_28923), .Q (new_AGEMA_signal_28924) ) ;
    buf_clk new_AGEMA_reg_buffer_7971 ( .C (clk), .D (new_AGEMA_signal_28926), .Q (new_AGEMA_signal_28927) ) ;
    buf_clk new_AGEMA_reg_buffer_7974 ( .C (clk), .D (new_AGEMA_signal_28929), .Q (new_AGEMA_signal_28930) ) ;
    buf_clk new_AGEMA_reg_buffer_7977 ( .C (clk), .D (new_AGEMA_signal_28932), .Q (new_AGEMA_signal_28933) ) ;
    buf_clk new_AGEMA_reg_buffer_7980 ( .C (clk), .D (new_AGEMA_signal_28935), .Q (new_AGEMA_signal_28936) ) ;
    buf_clk new_AGEMA_reg_buffer_7983 ( .C (clk), .D (new_AGEMA_signal_28938), .Q (new_AGEMA_signal_28939) ) ;
    buf_clk new_AGEMA_reg_buffer_7986 ( .C (clk), .D (new_AGEMA_signal_28941), .Q (new_AGEMA_signal_28942) ) ;
    buf_clk new_AGEMA_reg_buffer_7989 ( .C (clk), .D (new_AGEMA_signal_28944), .Q (new_AGEMA_signal_28945) ) ;
    buf_clk new_AGEMA_reg_buffer_7992 ( .C (clk), .D (new_AGEMA_signal_28947), .Q (new_AGEMA_signal_28948) ) ;
    buf_clk new_AGEMA_reg_buffer_7995 ( .C (clk), .D (new_AGEMA_signal_28950), .Q (new_AGEMA_signal_28951) ) ;
    buf_clk new_AGEMA_reg_buffer_7998 ( .C (clk), .D (new_AGEMA_signal_28953), .Q (new_AGEMA_signal_28954) ) ;
    buf_clk new_AGEMA_reg_buffer_8001 ( .C (clk), .D (new_AGEMA_signal_28956), .Q (new_AGEMA_signal_28957) ) ;
    buf_clk new_AGEMA_reg_buffer_8004 ( .C (clk), .D (new_AGEMA_signal_28959), .Q (new_AGEMA_signal_28960) ) ;
    buf_clk new_AGEMA_reg_buffer_8007 ( .C (clk), .D (new_AGEMA_signal_28962), .Q (new_AGEMA_signal_28963) ) ;
    buf_clk new_AGEMA_reg_buffer_8010 ( .C (clk), .D (new_AGEMA_signal_28965), .Q (new_AGEMA_signal_28966) ) ;
    buf_clk new_AGEMA_reg_buffer_8013 ( .C (clk), .D (new_AGEMA_signal_28968), .Q (new_AGEMA_signal_28969) ) ;
    buf_clk new_AGEMA_reg_buffer_8016 ( .C (clk), .D (new_AGEMA_signal_28971), .Q (new_AGEMA_signal_28972) ) ;
    buf_clk new_AGEMA_reg_buffer_8019 ( .C (clk), .D (new_AGEMA_signal_28974), .Q (new_AGEMA_signal_28975) ) ;
    buf_clk new_AGEMA_reg_buffer_8022 ( .C (clk), .D (new_AGEMA_signal_28977), .Q (new_AGEMA_signal_28978) ) ;
    buf_clk new_AGEMA_reg_buffer_8025 ( .C (clk), .D (new_AGEMA_signal_28980), .Q (new_AGEMA_signal_28981) ) ;
    buf_clk new_AGEMA_reg_buffer_8028 ( .C (clk), .D (new_AGEMA_signal_28983), .Q (new_AGEMA_signal_28984) ) ;
    buf_clk new_AGEMA_reg_buffer_8031 ( .C (clk), .D (new_AGEMA_signal_28986), .Q (new_AGEMA_signal_28987) ) ;
    buf_clk new_AGEMA_reg_buffer_8034 ( .C (clk), .D (new_AGEMA_signal_28989), .Q (new_AGEMA_signal_28990) ) ;
    buf_clk new_AGEMA_reg_buffer_8037 ( .C (clk), .D (new_AGEMA_signal_28992), .Q (new_AGEMA_signal_28993) ) ;
    buf_clk new_AGEMA_reg_buffer_8040 ( .C (clk), .D (new_AGEMA_signal_28995), .Q (new_AGEMA_signal_28996) ) ;
    buf_clk new_AGEMA_reg_buffer_8043 ( .C (clk), .D (new_AGEMA_signal_28998), .Q (new_AGEMA_signal_28999) ) ;
    buf_clk new_AGEMA_reg_buffer_8046 ( .C (clk), .D (new_AGEMA_signal_29001), .Q (new_AGEMA_signal_29002) ) ;
    buf_clk new_AGEMA_reg_buffer_8049 ( .C (clk), .D (new_AGEMA_signal_29004), .Q (new_AGEMA_signal_29005) ) ;
    buf_clk new_AGEMA_reg_buffer_8052 ( .C (clk), .D (new_AGEMA_signal_29007), .Q (new_AGEMA_signal_29008) ) ;
    buf_clk new_AGEMA_reg_buffer_8055 ( .C (clk), .D (new_AGEMA_signal_29010), .Q (new_AGEMA_signal_29011) ) ;
    buf_clk new_AGEMA_reg_buffer_8058 ( .C (clk), .D (new_AGEMA_signal_29013), .Q (new_AGEMA_signal_29014) ) ;
    buf_clk new_AGEMA_reg_buffer_8061 ( .C (clk), .D (new_AGEMA_signal_29016), .Q (new_AGEMA_signal_29017) ) ;
    buf_clk new_AGEMA_reg_buffer_8064 ( .C (clk), .D (new_AGEMA_signal_29019), .Q (new_AGEMA_signal_29020) ) ;
    buf_clk new_AGEMA_reg_buffer_8067 ( .C (clk), .D (new_AGEMA_signal_29022), .Q (new_AGEMA_signal_29023) ) ;
    buf_clk new_AGEMA_reg_buffer_8070 ( .C (clk), .D (new_AGEMA_signal_29025), .Q (new_AGEMA_signal_29026) ) ;
    buf_clk new_AGEMA_reg_buffer_8073 ( .C (clk), .D (new_AGEMA_signal_29028), .Q (new_AGEMA_signal_29029) ) ;
    buf_clk new_AGEMA_reg_buffer_8076 ( .C (clk), .D (new_AGEMA_signal_29031), .Q (new_AGEMA_signal_29032) ) ;
    buf_clk new_AGEMA_reg_buffer_8079 ( .C (clk), .D (new_AGEMA_signal_29034), .Q (new_AGEMA_signal_29035) ) ;
    buf_clk new_AGEMA_reg_buffer_8082 ( .C (clk), .D (new_AGEMA_signal_29037), .Q (new_AGEMA_signal_29038) ) ;
    buf_clk new_AGEMA_reg_buffer_8085 ( .C (clk), .D (new_AGEMA_signal_29040), .Q (new_AGEMA_signal_29041) ) ;
    buf_clk new_AGEMA_reg_buffer_8088 ( .C (clk), .D (new_AGEMA_signal_29043), .Q (new_AGEMA_signal_29044) ) ;
    buf_clk new_AGEMA_reg_buffer_8091 ( .C (clk), .D (new_AGEMA_signal_29046), .Q (new_AGEMA_signal_29047) ) ;
    buf_clk new_AGEMA_reg_buffer_8094 ( .C (clk), .D (new_AGEMA_signal_29049), .Q (new_AGEMA_signal_29050) ) ;
    buf_clk new_AGEMA_reg_buffer_8097 ( .C (clk), .D (new_AGEMA_signal_29052), .Q (new_AGEMA_signal_29053) ) ;
    buf_clk new_AGEMA_reg_buffer_8100 ( .C (clk), .D (new_AGEMA_signal_29055), .Q (new_AGEMA_signal_29056) ) ;
    buf_clk new_AGEMA_reg_buffer_8103 ( .C (clk), .D (new_AGEMA_signal_29058), .Q (new_AGEMA_signal_29059) ) ;
    buf_clk new_AGEMA_reg_buffer_8106 ( .C (clk), .D (new_AGEMA_signal_29061), .Q (new_AGEMA_signal_29062) ) ;
    buf_clk new_AGEMA_reg_buffer_8109 ( .C (clk), .D (new_AGEMA_signal_29064), .Q (new_AGEMA_signal_29065) ) ;
    buf_clk new_AGEMA_reg_buffer_8112 ( .C (clk), .D (new_AGEMA_signal_29067), .Q (new_AGEMA_signal_29068) ) ;
    buf_clk new_AGEMA_reg_buffer_8115 ( .C (clk), .D (new_AGEMA_signal_29070), .Q (new_AGEMA_signal_29071) ) ;
    buf_clk new_AGEMA_reg_buffer_8118 ( .C (clk), .D (new_AGEMA_signal_29073), .Q (new_AGEMA_signal_29074) ) ;
    buf_clk new_AGEMA_reg_buffer_8121 ( .C (clk), .D (new_AGEMA_signal_29076), .Q (new_AGEMA_signal_29077) ) ;
    buf_clk new_AGEMA_reg_buffer_8124 ( .C (clk), .D (new_AGEMA_signal_29079), .Q (new_AGEMA_signal_29080) ) ;
    buf_clk new_AGEMA_reg_buffer_8127 ( .C (clk), .D (new_AGEMA_signal_29082), .Q (new_AGEMA_signal_29083) ) ;
    buf_clk new_AGEMA_reg_buffer_8130 ( .C (clk), .D (new_AGEMA_signal_29085), .Q (new_AGEMA_signal_29086) ) ;
    buf_clk new_AGEMA_reg_buffer_8133 ( .C (clk), .D (new_AGEMA_signal_29088), .Q (new_AGEMA_signal_29089) ) ;
    buf_clk new_AGEMA_reg_buffer_8136 ( .C (clk), .D (new_AGEMA_signal_29091), .Q (new_AGEMA_signal_29092) ) ;
    buf_clk new_AGEMA_reg_buffer_8139 ( .C (clk), .D (new_AGEMA_signal_29094), .Q (new_AGEMA_signal_29095) ) ;
    buf_clk new_AGEMA_reg_buffer_8142 ( .C (clk), .D (new_AGEMA_signal_29097), .Q (new_AGEMA_signal_29098) ) ;
    buf_clk new_AGEMA_reg_buffer_8145 ( .C (clk), .D (new_AGEMA_signal_29100), .Q (new_AGEMA_signal_29101) ) ;
    buf_clk new_AGEMA_reg_buffer_8148 ( .C (clk), .D (new_AGEMA_signal_29103), .Q (new_AGEMA_signal_29104) ) ;
    buf_clk new_AGEMA_reg_buffer_8151 ( .C (clk), .D (new_AGEMA_signal_29106), .Q (new_AGEMA_signal_29107) ) ;
    buf_clk new_AGEMA_reg_buffer_8154 ( .C (clk), .D (new_AGEMA_signal_29109), .Q (new_AGEMA_signal_29110) ) ;
    buf_clk new_AGEMA_reg_buffer_8157 ( .C (clk), .D (new_AGEMA_signal_29112), .Q (new_AGEMA_signal_29113) ) ;
    buf_clk new_AGEMA_reg_buffer_8160 ( .C (clk), .D (new_AGEMA_signal_29115), .Q (new_AGEMA_signal_29116) ) ;
    buf_clk new_AGEMA_reg_buffer_8163 ( .C (clk), .D (new_AGEMA_signal_29118), .Q (new_AGEMA_signal_29119) ) ;
    buf_clk new_AGEMA_reg_buffer_8166 ( .C (clk), .D (new_AGEMA_signal_29121), .Q (new_AGEMA_signal_29122) ) ;
    buf_clk new_AGEMA_reg_buffer_8169 ( .C (clk), .D (new_AGEMA_signal_29124), .Q (new_AGEMA_signal_29125) ) ;
    buf_clk new_AGEMA_reg_buffer_8172 ( .C (clk), .D (new_AGEMA_signal_29127), .Q (new_AGEMA_signal_29128) ) ;
    buf_clk new_AGEMA_reg_buffer_8175 ( .C (clk), .D (new_AGEMA_signal_29130), .Q (new_AGEMA_signal_29131) ) ;
    buf_clk new_AGEMA_reg_buffer_8178 ( .C (clk), .D (new_AGEMA_signal_29133), .Q (new_AGEMA_signal_29134) ) ;
    buf_clk new_AGEMA_reg_buffer_8181 ( .C (clk), .D (new_AGEMA_signal_29136), .Q (new_AGEMA_signal_29137) ) ;
    buf_clk new_AGEMA_reg_buffer_8184 ( .C (clk), .D (new_AGEMA_signal_29139), .Q (new_AGEMA_signal_29140) ) ;
    buf_clk new_AGEMA_reg_buffer_8187 ( .C (clk), .D (new_AGEMA_signal_29142), .Q (new_AGEMA_signal_29143) ) ;
    buf_clk new_AGEMA_reg_buffer_8190 ( .C (clk), .D (new_AGEMA_signal_29145), .Q (new_AGEMA_signal_29146) ) ;
    buf_clk new_AGEMA_reg_buffer_8193 ( .C (clk), .D (new_AGEMA_signal_29148), .Q (new_AGEMA_signal_29149) ) ;
    buf_clk new_AGEMA_reg_buffer_8196 ( .C (clk), .D (new_AGEMA_signal_29151), .Q (new_AGEMA_signal_29152) ) ;
    buf_clk new_AGEMA_reg_buffer_8199 ( .C (clk), .D (new_AGEMA_signal_29154), .Q (new_AGEMA_signal_29155) ) ;
    buf_clk new_AGEMA_reg_buffer_8202 ( .C (clk), .D (new_AGEMA_signal_29157), .Q (new_AGEMA_signal_29158) ) ;
    buf_clk new_AGEMA_reg_buffer_8205 ( .C (clk), .D (new_AGEMA_signal_29160), .Q (new_AGEMA_signal_29161) ) ;
    buf_clk new_AGEMA_reg_buffer_8208 ( .C (clk), .D (new_AGEMA_signal_29163), .Q (new_AGEMA_signal_29164) ) ;
    buf_clk new_AGEMA_reg_buffer_8211 ( .C (clk), .D (new_AGEMA_signal_29166), .Q (new_AGEMA_signal_29167) ) ;
    buf_clk new_AGEMA_reg_buffer_8214 ( .C (clk), .D (new_AGEMA_signal_29169), .Q (new_AGEMA_signal_29170) ) ;
    buf_clk new_AGEMA_reg_buffer_8217 ( .C (clk), .D (new_AGEMA_signal_29172), .Q (new_AGEMA_signal_29173) ) ;
    buf_clk new_AGEMA_reg_buffer_8220 ( .C (clk), .D (new_AGEMA_signal_29175), .Q (new_AGEMA_signal_29176) ) ;
    buf_clk new_AGEMA_reg_buffer_8223 ( .C (clk), .D (new_AGEMA_signal_29178), .Q (new_AGEMA_signal_29179) ) ;
    buf_clk new_AGEMA_reg_buffer_8226 ( .C (clk), .D (new_AGEMA_signal_29181), .Q (new_AGEMA_signal_29182) ) ;
    buf_clk new_AGEMA_reg_buffer_8229 ( .C (clk), .D (new_AGEMA_signal_29184), .Q (new_AGEMA_signal_29185) ) ;
    buf_clk new_AGEMA_reg_buffer_8232 ( .C (clk), .D (new_AGEMA_signal_29187), .Q (new_AGEMA_signal_29188) ) ;
    buf_clk new_AGEMA_reg_buffer_8235 ( .C (clk), .D (new_AGEMA_signal_29190), .Q (new_AGEMA_signal_29191) ) ;
    buf_clk new_AGEMA_reg_buffer_8238 ( .C (clk), .D (new_AGEMA_signal_29193), .Q (new_AGEMA_signal_29194) ) ;
    buf_clk new_AGEMA_reg_buffer_8241 ( .C (clk), .D (new_AGEMA_signal_29196), .Q (new_AGEMA_signal_29197) ) ;
    buf_clk new_AGEMA_reg_buffer_8244 ( .C (clk), .D (new_AGEMA_signal_29199), .Q (new_AGEMA_signal_29200) ) ;
    buf_clk new_AGEMA_reg_buffer_8247 ( .C (clk), .D (new_AGEMA_signal_29202), .Q (new_AGEMA_signal_29203) ) ;
    buf_clk new_AGEMA_reg_buffer_8250 ( .C (clk), .D (new_AGEMA_signal_29205), .Q (new_AGEMA_signal_29206) ) ;
    buf_clk new_AGEMA_reg_buffer_8253 ( .C (clk), .D (new_AGEMA_signal_29208), .Q (new_AGEMA_signal_29209) ) ;
    buf_clk new_AGEMA_reg_buffer_8256 ( .C (clk), .D (new_AGEMA_signal_29211), .Q (new_AGEMA_signal_29212) ) ;
    buf_clk new_AGEMA_reg_buffer_8259 ( .C (clk), .D (new_AGEMA_signal_29214), .Q (new_AGEMA_signal_29215) ) ;
    buf_clk new_AGEMA_reg_buffer_8262 ( .C (clk), .D (new_AGEMA_signal_29217), .Q (new_AGEMA_signal_29218) ) ;
    buf_clk new_AGEMA_reg_buffer_8265 ( .C (clk), .D (new_AGEMA_signal_29220), .Q (new_AGEMA_signal_29221) ) ;
    buf_clk new_AGEMA_reg_buffer_8268 ( .C (clk), .D (new_AGEMA_signal_29223), .Q (new_AGEMA_signal_29224) ) ;
    buf_clk new_AGEMA_reg_buffer_8271 ( .C (clk), .D (new_AGEMA_signal_29226), .Q (new_AGEMA_signal_29227) ) ;
    buf_clk new_AGEMA_reg_buffer_8274 ( .C (clk), .D (new_AGEMA_signal_29229), .Q (new_AGEMA_signal_29230) ) ;
    buf_clk new_AGEMA_reg_buffer_8277 ( .C (clk), .D (new_AGEMA_signal_29232), .Q (new_AGEMA_signal_29233) ) ;
    buf_clk new_AGEMA_reg_buffer_8280 ( .C (clk), .D (new_AGEMA_signal_29235), .Q (new_AGEMA_signal_29236) ) ;
    buf_clk new_AGEMA_reg_buffer_8283 ( .C (clk), .D (new_AGEMA_signal_29238), .Q (new_AGEMA_signal_29239) ) ;
    buf_clk new_AGEMA_reg_buffer_8286 ( .C (clk), .D (new_AGEMA_signal_29241), .Q (new_AGEMA_signal_29242) ) ;
    buf_clk new_AGEMA_reg_buffer_8289 ( .C (clk), .D (new_AGEMA_signal_29244), .Q (new_AGEMA_signal_29245) ) ;
    buf_clk new_AGEMA_reg_buffer_8292 ( .C (clk), .D (new_AGEMA_signal_29247), .Q (new_AGEMA_signal_29248) ) ;
    buf_clk new_AGEMA_reg_buffer_8295 ( .C (clk), .D (new_AGEMA_signal_29250), .Q (new_AGEMA_signal_29251) ) ;
    buf_clk new_AGEMA_reg_buffer_8298 ( .C (clk), .D (new_AGEMA_signal_29253), .Q (new_AGEMA_signal_29254) ) ;
    buf_clk new_AGEMA_reg_buffer_8301 ( .C (clk), .D (new_AGEMA_signal_29256), .Q (new_AGEMA_signal_29257) ) ;
    buf_clk new_AGEMA_reg_buffer_8304 ( .C (clk), .D (new_AGEMA_signal_29259), .Q (new_AGEMA_signal_29260) ) ;
    buf_clk new_AGEMA_reg_buffer_8307 ( .C (clk), .D (new_AGEMA_signal_29262), .Q (new_AGEMA_signal_29263) ) ;
    buf_clk new_AGEMA_reg_buffer_8310 ( .C (clk), .D (new_AGEMA_signal_29265), .Q (new_AGEMA_signal_29266) ) ;
    buf_clk new_AGEMA_reg_buffer_8313 ( .C (clk), .D (new_AGEMA_signal_29268), .Q (new_AGEMA_signal_29269) ) ;
    buf_clk new_AGEMA_reg_buffer_8316 ( .C (clk), .D (new_AGEMA_signal_29271), .Q (new_AGEMA_signal_29272) ) ;
    buf_clk new_AGEMA_reg_buffer_8319 ( .C (clk), .D (new_AGEMA_signal_29274), .Q (new_AGEMA_signal_29275) ) ;
    buf_clk new_AGEMA_reg_buffer_8322 ( .C (clk), .D (new_AGEMA_signal_29277), .Q (new_AGEMA_signal_29278) ) ;
    buf_clk new_AGEMA_reg_buffer_8325 ( .C (clk), .D (new_AGEMA_signal_29280), .Q (new_AGEMA_signal_29281) ) ;
    buf_clk new_AGEMA_reg_buffer_8328 ( .C (clk), .D (new_AGEMA_signal_29283), .Q (new_AGEMA_signal_29284) ) ;
    buf_clk new_AGEMA_reg_buffer_8331 ( .C (clk), .D (new_AGEMA_signal_29286), .Q (new_AGEMA_signal_29287) ) ;
    buf_clk new_AGEMA_reg_buffer_8334 ( .C (clk), .D (new_AGEMA_signal_29289), .Q (new_AGEMA_signal_29290) ) ;
    buf_clk new_AGEMA_reg_buffer_8337 ( .C (clk), .D (new_AGEMA_signal_29292), .Q (new_AGEMA_signal_29293) ) ;
    buf_clk new_AGEMA_reg_buffer_8340 ( .C (clk), .D (new_AGEMA_signal_29295), .Q (new_AGEMA_signal_29296) ) ;
    buf_clk new_AGEMA_reg_buffer_8343 ( .C (clk), .D (new_AGEMA_signal_29298), .Q (new_AGEMA_signal_29299) ) ;
    buf_clk new_AGEMA_reg_buffer_8346 ( .C (clk), .D (new_AGEMA_signal_29301), .Q (new_AGEMA_signal_29302) ) ;
    buf_clk new_AGEMA_reg_buffer_8349 ( .C (clk), .D (new_AGEMA_signal_29304), .Q (new_AGEMA_signal_29305) ) ;
    buf_clk new_AGEMA_reg_buffer_8352 ( .C (clk), .D (new_AGEMA_signal_29307), .Q (new_AGEMA_signal_29308) ) ;
    buf_clk new_AGEMA_reg_buffer_8355 ( .C (clk), .D (new_AGEMA_signal_29310), .Q (new_AGEMA_signal_29311) ) ;
    buf_clk new_AGEMA_reg_buffer_8358 ( .C (clk), .D (new_AGEMA_signal_29313), .Q (new_AGEMA_signal_29314) ) ;
    buf_clk new_AGEMA_reg_buffer_8361 ( .C (clk), .D (new_AGEMA_signal_29316), .Q (new_AGEMA_signal_29317) ) ;
    buf_clk new_AGEMA_reg_buffer_8364 ( .C (clk), .D (new_AGEMA_signal_29319), .Q (new_AGEMA_signal_29320) ) ;
    buf_clk new_AGEMA_reg_buffer_8367 ( .C (clk), .D (new_AGEMA_signal_29322), .Q (new_AGEMA_signal_29323) ) ;
    buf_clk new_AGEMA_reg_buffer_8370 ( .C (clk), .D (new_AGEMA_signal_29325), .Q (new_AGEMA_signal_29326) ) ;
    buf_clk new_AGEMA_reg_buffer_8373 ( .C (clk), .D (new_AGEMA_signal_29328), .Q (new_AGEMA_signal_29329) ) ;
    buf_clk new_AGEMA_reg_buffer_8376 ( .C (clk), .D (new_AGEMA_signal_29331), .Q (new_AGEMA_signal_29332) ) ;
    buf_clk new_AGEMA_reg_buffer_8379 ( .C (clk), .D (new_AGEMA_signal_29334), .Q (new_AGEMA_signal_29335) ) ;
    buf_clk new_AGEMA_reg_buffer_8382 ( .C (clk), .D (new_AGEMA_signal_29337), .Q (new_AGEMA_signal_29338) ) ;
    buf_clk new_AGEMA_reg_buffer_8385 ( .C (clk), .D (new_AGEMA_signal_29340), .Q (new_AGEMA_signal_29341) ) ;
    buf_clk new_AGEMA_reg_buffer_8388 ( .C (clk), .D (new_AGEMA_signal_29343), .Q (new_AGEMA_signal_29344) ) ;
    buf_clk new_AGEMA_reg_buffer_8391 ( .C (clk), .D (new_AGEMA_signal_29346), .Q (new_AGEMA_signal_29347) ) ;
    buf_clk new_AGEMA_reg_buffer_8394 ( .C (clk), .D (new_AGEMA_signal_29349), .Q (new_AGEMA_signal_29350) ) ;
    buf_clk new_AGEMA_reg_buffer_8397 ( .C (clk), .D (new_AGEMA_signal_29352), .Q (new_AGEMA_signal_29353) ) ;
    buf_clk new_AGEMA_reg_buffer_8400 ( .C (clk), .D (new_AGEMA_signal_29355), .Q (new_AGEMA_signal_29356) ) ;
    buf_clk new_AGEMA_reg_buffer_8403 ( .C (clk), .D (new_AGEMA_signal_29358), .Q (new_AGEMA_signal_29359) ) ;
    buf_clk new_AGEMA_reg_buffer_8406 ( .C (clk), .D (new_AGEMA_signal_29361), .Q (new_AGEMA_signal_29362) ) ;
    buf_clk new_AGEMA_reg_buffer_8409 ( .C (clk), .D (new_AGEMA_signal_29364), .Q (new_AGEMA_signal_29365) ) ;
    buf_clk new_AGEMA_reg_buffer_8412 ( .C (clk), .D (new_AGEMA_signal_29367), .Q (new_AGEMA_signal_29368) ) ;
    buf_clk new_AGEMA_reg_buffer_8415 ( .C (clk), .D (new_AGEMA_signal_29370), .Q (new_AGEMA_signal_29371) ) ;
    buf_clk new_AGEMA_reg_buffer_8418 ( .C (clk), .D (new_AGEMA_signal_29373), .Q (new_AGEMA_signal_29374) ) ;
    buf_clk new_AGEMA_reg_buffer_8421 ( .C (clk), .D (new_AGEMA_signal_29376), .Q (new_AGEMA_signal_29377) ) ;
    buf_clk new_AGEMA_reg_buffer_8424 ( .C (clk), .D (new_AGEMA_signal_29379), .Q (new_AGEMA_signal_29380) ) ;
    buf_clk new_AGEMA_reg_buffer_8427 ( .C (clk), .D (new_AGEMA_signal_29382), .Q (new_AGEMA_signal_29383) ) ;
    buf_clk new_AGEMA_reg_buffer_8430 ( .C (clk), .D (new_AGEMA_signal_29385), .Q (new_AGEMA_signal_29386) ) ;
    buf_clk new_AGEMA_reg_buffer_8433 ( .C (clk), .D (new_AGEMA_signal_29388), .Q (new_AGEMA_signal_29389) ) ;
    buf_clk new_AGEMA_reg_buffer_8436 ( .C (clk), .D (new_AGEMA_signal_29391), .Q (new_AGEMA_signal_29392) ) ;
    buf_clk new_AGEMA_reg_buffer_8439 ( .C (clk), .D (new_AGEMA_signal_29394), .Q (new_AGEMA_signal_29395) ) ;
    buf_clk new_AGEMA_reg_buffer_8442 ( .C (clk), .D (new_AGEMA_signal_29397), .Q (new_AGEMA_signal_29398) ) ;
    buf_clk new_AGEMA_reg_buffer_8445 ( .C (clk), .D (new_AGEMA_signal_29400), .Q (new_AGEMA_signal_29401) ) ;
    buf_clk new_AGEMA_reg_buffer_8448 ( .C (clk), .D (new_AGEMA_signal_29403), .Q (new_AGEMA_signal_29404) ) ;
    buf_clk new_AGEMA_reg_buffer_8451 ( .C (clk), .D (new_AGEMA_signal_29406), .Q (new_AGEMA_signal_29407) ) ;
    buf_clk new_AGEMA_reg_buffer_8454 ( .C (clk), .D (new_AGEMA_signal_29409), .Q (new_AGEMA_signal_29410) ) ;
    buf_clk new_AGEMA_reg_buffer_8457 ( .C (clk), .D (new_AGEMA_signal_29412), .Q (new_AGEMA_signal_29413) ) ;
    buf_clk new_AGEMA_reg_buffer_8460 ( .C (clk), .D (new_AGEMA_signal_29415), .Q (new_AGEMA_signal_29416) ) ;
    buf_clk new_AGEMA_reg_buffer_8463 ( .C (clk), .D (new_AGEMA_signal_29418), .Q (new_AGEMA_signal_29419) ) ;
    buf_clk new_AGEMA_reg_buffer_8466 ( .C (clk), .D (new_AGEMA_signal_29421), .Q (new_AGEMA_signal_29422) ) ;
    buf_clk new_AGEMA_reg_buffer_8469 ( .C (clk), .D (new_AGEMA_signal_29424), .Q (new_AGEMA_signal_29425) ) ;
    buf_clk new_AGEMA_reg_buffer_8472 ( .C (clk), .D (new_AGEMA_signal_29427), .Q (new_AGEMA_signal_29428) ) ;
    buf_clk new_AGEMA_reg_buffer_8475 ( .C (clk), .D (new_AGEMA_signal_29430), .Q (new_AGEMA_signal_29431) ) ;
    buf_clk new_AGEMA_reg_buffer_8478 ( .C (clk), .D (new_AGEMA_signal_29433), .Q (new_AGEMA_signal_29434) ) ;
    buf_clk new_AGEMA_reg_buffer_8481 ( .C (clk), .D (new_AGEMA_signal_29436), .Q (new_AGEMA_signal_29437) ) ;
    buf_clk new_AGEMA_reg_buffer_8484 ( .C (clk), .D (new_AGEMA_signal_29439), .Q (new_AGEMA_signal_29440) ) ;
    buf_clk new_AGEMA_reg_buffer_8487 ( .C (clk), .D (new_AGEMA_signal_29442), .Q (new_AGEMA_signal_29443) ) ;
    buf_clk new_AGEMA_reg_buffer_8490 ( .C (clk), .D (new_AGEMA_signal_29445), .Q (new_AGEMA_signal_29446) ) ;
    buf_clk new_AGEMA_reg_buffer_8493 ( .C (clk), .D (new_AGEMA_signal_29448), .Q (new_AGEMA_signal_29449) ) ;
    buf_clk new_AGEMA_reg_buffer_8496 ( .C (clk), .D (new_AGEMA_signal_29451), .Q (new_AGEMA_signal_29452) ) ;
    buf_clk new_AGEMA_reg_buffer_8499 ( .C (clk), .D (new_AGEMA_signal_29454), .Q (new_AGEMA_signal_29455) ) ;
    buf_clk new_AGEMA_reg_buffer_8502 ( .C (clk), .D (new_AGEMA_signal_29457), .Q (new_AGEMA_signal_29458) ) ;
    buf_clk new_AGEMA_reg_buffer_8505 ( .C (clk), .D (new_AGEMA_signal_29460), .Q (new_AGEMA_signal_29461) ) ;
    buf_clk new_AGEMA_reg_buffer_8508 ( .C (clk), .D (new_AGEMA_signal_29463), .Q (new_AGEMA_signal_29464) ) ;
    buf_clk new_AGEMA_reg_buffer_8511 ( .C (clk), .D (new_AGEMA_signal_29466), .Q (new_AGEMA_signal_29467) ) ;
    buf_clk new_AGEMA_reg_buffer_8514 ( .C (clk), .D (new_AGEMA_signal_29469), .Q (new_AGEMA_signal_29470) ) ;
    buf_clk new_AGEMA_reg_buffer_8517 ( .C (clk), .D (new_AGEMA_signal_29472), .Q (new_AGEMA_signal_29473) ) ;
    buf_clk new_AGEMA_reg_buffer_8520 ( .C (clk), .D (new_AGEMA_signal_29475), .Q (new_AGEMA_signal_29476) ) ;
    buf_clk new_AGEMA_reg_buffer_8523 ( .C (clk), .D (new_AGEMA_signal_29478), .Q (new_AGEMA_signal_29479) ) ;
    buf_clk new_AGEMA_reg_buffer_8526 ( .C (clk), .D (new_AGEMA_signal_29481), .Q (new_AGEMA_signal_29482) ) ;
    buf_clk new_AGEMA_reg_buffer_8529 ( .C (clk), .D (new_AGEMA_signal_29484), .Q (new_AGEMA_signal_29485) ) ;
    buf_clk new_AGEMA_reg_buffer_8532 ( .C (clk), .D (new_AGEMA_signal_29487), .Q (new_AGEMA_signal_29488) ) ;
    buf_clk new_AGEMA_reg_buffer_8535 ( .C (clk), .D (new_AGEMA_signal_29490), .Q (new_AGEMA_signal_29491) ) ;
    buf_clk new_AGEMA_reg_buffer_8538 ( .C (clk), .D (new_AGEMA_signal_29493), .Q (new_AGEMA_signal_29494) ) ;
    buf_clk new_AGEMA_reg_buffer_8541 ( .C (clk), .D (new_AGEMA_signal_29496), .Q (new_AGEMA_signal_29497) ) ;
    buf_clk new_AGEMA_reg_buffer_8544 ( .C (clk), .D (new_AGEMA_signal_29499), .Q (new_AGEMA_signal_29500) ) ;
    buf_clk new_AGEMA_reg_buffer_8547 ( .C (clk), .D (new_AGEMA_signal_29502), .Q (new_AGEMA_signal_29503) ) ;
    buf_clk new_AGEMA_reg_buffer_8550 ( .C (clk), .D (new_AGEMA_signal_29505), .Q (new_AGEMA_signal_29506) ) ;
    buf_clk new_AGEMA_reg_buffer_8553 ( .C (clk), .D (new_AGEMA_signal_29508), .Q (new_AGEMA_signal_29509) ) ;
    buf_clk new_AGEMA_reg_buffer_8556 ( .C (clk), .D (new_AGEMA_signal_29511), .Q (new_AGEMA_signal_29512) ) ;
    buf_clk new_AGEMA_reg_buffer_8559 ( .C (clk), .D (new_AGEMA_signal_29514), .Q (new_AGEMA_signal_29515) ) ;
    buf_clk new_AGEMA_reg_buffer_8562 ( .C (clk), .D (new_AGEMA_signal_29517), .Q (new_AGEMA_signal_29518) ) ;
    buf_clk new_AGEMA_reg_buffer_8565 ( .C (clk), .D (new_AGEMA_signal_29520), .Q (new_AGEMA_signal_29521) ) ;
    buf_clk new_AGEMA_reg_buffer_8568 ( .C (clk), .D (new_AGEMA_signal_29523), .Q (new_AGEMA_signal_29524) ) ;
    buf_clk new_AGEMA_reg_buffer_8571 ( .C (clk), .D (new_AGEMA_signal_29526), .Q (new_AGEMA_signal_29527) ) ;
    buf_clk new_AGEMA_reg_buffer_8574 ( .C (clk), .D (new_AGEMA_signal_29529), .Q (new_AGEMA_signal_29530) ) ;
    buf_clk new_AGEMA_reg_buffer_8577 ( .C (clk), .D (new_AGEMA_signal_29532), .Q (new_AGEMA_signal_29533) ) ;
    buf_clk new_AGEMA_reg_buffer_8580 ( .C (clk), .D (new_AGEMA_signal_29535), .Q (new_AGEMA_signal_29536) ) ;
    buf_clk new_AGEMA_reg_buffer_8583 ( .C (clk), .D (new_AGEMA_signal_29538), .Q (new_AGEMA_signal_29539) ) ;
    buf_clk new_AGEMA_reg_buffer_8586 ( .C (clk), .D (new_AGEMA_signal_29541), .Q (new_AGEMA_signal_29542) ) ;
    buf_clk new_AGEMA_reg_buffer_8589 ( .C (clk), .D (new_AGEMA_signal_29544), .Q (new_AGEMA_signal_29545) ) ;
    buf_clk new_AGEMA_reg_buffer_8592 ( .C (clk), .D (new_AGEMA_signal_29547), .Q (new_AGEMA_signal_29548) ) ;
    buf_clk new_AGEMA_reg_buffer_8595 ( .C (clk), .D (new_AGEMA_signal_29550), .Q (new_AGEMA_signal_29551) ) ;
    buf_clk new_AGEMA_reg_buffer_8598 ( .C (clk), .D (new_AGEMA_signal_29553), .Q (new_AGEMA_signal_29554) ) ;
    buf_clk new_AGEMA_reg_buffer_8601 ( .C (clk), .D (new_AGEMA_signal_29556), .Q (new_AGEMA_signal_29557) ) ;
    buf_clk new_AGEMA_reg_buffer_8604 ( .C (clk), .D (new_AGEMA_signal_29559), .Q (new_AGEMA_signal_29560) ) ;
    buf_clk new_AGEMA_reg_buffer_8607 ( .C (clk), .D (new_AGEMA_signal_29562), .Q (new_AGEMA_signal_29563) ) ;
    buf_clk new_AGEMA_reg_buffer_8610 ( .C (clk), .D (new_AGEMA_signal_29565), .Q (new_AGEMA_signal_29566) ) ;
    buf_clk new_AGEMA_reg_buffer_8613 ( .C (clk), .D (new_AGEMA_signal_29568), .Q (new_AGEMA_signal_29569) ) ;
    buf_clk new_AGEMA_reg_buffer_8616 ( .C (clk), .D (new_AGEMA_signal_29571), .Q (new_AGEMA_signal_29572) ) ;
    buf_clk new_AGEMA_reg_buffer_8619 ( .C (clk), .D (new_AGEMA_signal_29574), .Q (new_AGEMA_signal_29575) ) ;
    buf_clk new_AGEMA_reg_buffer_8622 ( .C (clk), .D (new_AGEMA_signal_29577), .Q (new_AGEMA_signal_29578) ) ;
    buf_clk new_AGEMA_reg_buffer_8625 ( .C (clk), .D (new_AGEMA_signal_29580), .Q (new_AGEMA_signal_29581) ) ;
    buf_clk new_AGEMA_reg_buffer_8628 ( .C (clk), .D (new_AGEMA_signal_29583), .Q (new_AGEMA_signal_29584) ) ;
    buf_clk new_AGEMA_reg_buffer_8631 ( .C (clk), .D (new_AGEMA_signal_29586), .Q (new_AGEMA_signal_29587) ) ;
    buf_clk new_AGEMA_reg_buffer_8634 ( .C (clk), .D (new_AGEMA_signal_29589), .Q (new_AGEMA_signal_29590) ) ;
    buf_clk new_AGEMA_reg_buffer_8637 ( .C (clk), .D (new_AGEMA_signal_29592), .Q (new_AGEMA_signal_29593) ) ;
    buf_clk new_AGEMA_reg_buffer_8640 ( .C (clk), .D (new_AGEMA_signal_29595), .Q (new_AGEMA_signal_29596) ) ;
    buf_clk new_AGEMA_reg_buffer_8643 ( .C (clk), .D (new_AGEMA_signal_29598), .Q (new_AGEMA_signal_29599) ) ;
    buf_clk new_AGEMA_reg_buffer_8646 ( .C (clk), .D (new_AGEMA_signal_29601), .Q (new_AGEMA_signal_29602) ) ;
    buf_clk new_AGEMA_reg_buffer_8649 ( .C (clk), .D (new_AGEMA_signal_29604), .Q (new_AGEMA_signal_29605) ) ;
    buf_clk new_AGEMA_reg_buffer_8652 ( .C (clk), .D (new_AGEMA_signal_29607), .Q (new_AGEMA_signal_29608) ) ;
    buf_clk new_AGEMA_reg_buffer_8655 ( .C (clk), .D (new_AGEMA_signal_29610), .Q (new_AGEMA_signal_29611) ) ;
    buf_clk new_AGEMA_reg_buffer_8658 ( .C (clk), .D (new_AGEMA_signal_29613), .Q (new_AGEMA_signal_29614) ) ;
    buf_clk new_AGEMA_reg_buffer_8661 ( .C (clk), .D (new_AGEMA_signal_29616), .Q (new_AGEMA_signal_29617) ) ;
    buf_clk new_AGEMA_reg_buffer_8664 ( .C (clk), .D (new_AGEMA_signal_29619), .Q (new_AGEMA_signal_29620) ) ;
    buf_clk new_AGEMA_reg_buffer_8667 ( .C (clk), .D (new_AGEMA_signal_29622), .Q (new_AGEMA_signal_29623) ) ;
    buf_clk new_AGEMA_reg_buffer_8670 ( .C (clk), .D (new_AGEMA_signal_29625), .Q (new_AGEMA_signal_29626) ) ;
    buf_clk new_AGEMA_reg_buffer_8673 ( .C (clk), .D (new_AGEMA_signal_29628), .Q (new_AGEMA_signal_29629) ) ;
    buf_clk new_AGEMA_reg_buffer_8676 ( .C (clk), .D (new_AGEMA_signal_29631), .Q (new_AGEMA_signal_29632) ) ;
    buf_clk new_AGEMA_reg_buffer_8679 ( .C (clk), .D (new_AGEMA_signal_29634), .Q (new_AGEMA_signal_29635) ) ;
    buf_clk new_AGEMA_reg_buffer_8682 ( .C (clk), .D (new_AGEMA_signal_29637), .Q (new_AGEMA_signal_29638) ) ;
    buf_clk new_AGEMA_reg_buffer_8685 ( .C (clk), .D (new_AGEMA_signal_29640), .Q (new_AGEMA_signal_29641) ) ;
    buf_clk new_AGEMA_reg_buffer_8688 ( .C (clk), .D (new_AGEMA_signal_29643), .Q (new_AGEMA_signal_29644) ) ;
    buf_clk new_AGEMA_reg_buffer_8691 ( .C (clk), .D (new_AGEMA_signal_29646), .Q (new_AGEMA_signal_29647) ) ;
    buf_clk new_AGEMA_reg_buffer_8694 ( .C (clk), .D (new_AGEMA_signal_29649), .Q (new_AGEMA_signal_29650) ) ;
    buf_clk new_AGEMA_reg_buffer_8697 ( .C (clk), .D (new_AGEMA_signal_29652), .Q (new_AGEMA_signal_29653) ) ;
    buf_clk new_AGEMA_reg_buffer_8700 ( .C (clk), .D (new_AGEMA_signal_29655), .Q (new_AGEMA_signal_29656) ) ;
    buf_clk new_AGEMA_reg_buffer_8703 ( .C (clk), .D (new_AGEMA_signal_29658), .Q (new_AGEMA_signal_29659) ) ;
    buf_clk new_AGEMA_reg_buffer_8706 ( .C (clk), .D (new_AGEMA_signal_29661), .Q (new_AGEMA_signal_29662) ) ;
    buf_clk new_AGEMA_reg_buffer_8709 ( .C (clk), .D (new_AGEMA_signal_29664), .Q (new_AGEMA_signal_29665) ) ;
    buf_clk new_AGEMA_reg_buffer_8712 ( .C (clk), .D (new_AGEMA_signal_29667), .Q (new_AGEMA_signal_29668) ) ;
    buf_clk new_AGEMA_reg_buffer_8715 ( .C (clk), .D (new_AGEMA_signal_29670), .Q (new_AGEMA_signal_29671) ) ;
    buf_clk new_AGEMA_reg_buffer_8718 ( .C (clk), .D (new_AGEMA_signal_29673), .Q (new_AGEMA_signal_29674) ) ;
    buf_clk new_AGEMA_reg_buffer_8721 ( .C (clk), .D (new_AGEMA_signal_29676), .Q (new_AGEMA_signal_29677) ) ;
    buf_clk new_AGEMA_reg_buffer_8724 ( .C (clk), .D (new_AGEMA_signal_29679), .Q (new_AGEMA_signal_29680) ) ;
    buf_clk new_AGEMA_reg_buffer_8727 ( .C (clk), .D (new_AGEMA_signal_29682), .Q (new_AGEMA_signal_29683) ) ;
    buf_clk new_AGEMA_reg_buffer_8730 ( .C (clk), .D (new_AGEMA_signal_29685), .Q (new_AGEMA_signal_29686) ) ;
    buf_clk new_AGEMA_reg_buffer_8733 ( .C (clk), .D (new_AGEMA_signal_29688), .Q (new_AGEMA_signal_29689) ) ;
    buf_clk new_AGEMA_reg_buffer_8736 ( .C (clk), .D (new_AGEMA_signal_29691), .Q (new_AGEMA_signal_29692) ) ;
    buf_clk new_AGEMA_reg_buffer_8739 ( .C (clk), .D (new_AGEMA_signal_29694), .Q (new_AGEMA_signal_29695) ) ;
    buf_clk new_AGEMA_reg_buffer_8742 ( .C (clk), .D (new_AGEMA_signal_29697), .Q (new_AGEMA_signal_29698) ) ;
    buf_clk new_AGEMA_reg_buffer_8745 ( .C (clk), .D (new_AGEMA_signal_29700), .Q (new_AGEMA_signal_29701) ) ;
    buf_clk new_AGEMA_reg_buffer_8748 ( .C (clk), .D (new_AGEMA_signal_29703), .Q (new_AGEMA_signal_29704) ) ;
    buf_clk new_AGEMA_reg_buffer_8751 ( .C (clk), .D (new_AGEMA_signal_29706), .Q (new_AGEMA_signal_29707) ) ;
    buf_clk new_AGEMA_reg_buffer_8754 ( .C (clk), .D (new_AGEMA_signal_29709), .Q (new_AGEMA_signal_29710) ) ;
    buf_clk new_AGEMA_reg_buffer_8757 ( .C (clk), .D (new_AGEMA_signal_29712), .Q (new_AGEMA_signal_29713) ) ;
    buf_clk new_AGEMA_reg_buffer_8760 ( .C (clk), .D (new_AGEMA_signal_29715), .Q (new_AGEMA_signal_29716) ) ;
    buf_clk new_AGEMA_reg_buffer_8763 ( .C (clk), .D (new_AGEMA_signal_29718), .Q (new_AGEMA_signal_29719) ) ;
    buf_clk new_AGEMA_reg_buffer_8766 ( .C (clk), .D (new_AGEMA_signal_29721), .Q (new_AGEMA_signal_29722) ) ;
    buf_clk new_AGEMA_reg_buffer_8769 ( .C (clk), .D (new_AGEMA_signal_29724), .Q (new_AGEMA_signal_29725) ) ;
    buf_clk new_AGEMA_reg_buffer_8772 ( .C (clk), .D (new_AGEMA_signal_29727), .Q (new_AGEMA_signal_29728) ) ;
    buf_clk new_AGEMA_reg_buffer_8775 ( .C (clk), .D (new_AGEMA_signal_29730), .Q (new_AGEMA_signal_29731) ) ;
    buf_clk new_AGEMA_reg_buffer_8778 ( .C (clk), .D (new_AGEMA_signal_29733), .Q (new_AGEMA_signal_29734) ) ;
    buf_clk new_AGEMA_reg_buffer_8781 ( .C (clk), .D (new_AGEMA_signal_29736), .Q (new_AGEMA_signal_29737) ) ;
    buf_clk new_AGEMA_reg_buffer_8784 ( .C (clk), .D (new_AGEMA_signal_29739), .Q (new_AGEMA_signal_29740) ) ;
    buf_clk new_AGEMA_reg_buffer_8787 ( .C (clk), .D (new_AGEMA_signal_29742), .Q (new_AGEMA_signal_29743) ) ;
    buf_clk new_AGEMA_reg_buffer_8790 ( .C (clk), .D (new_AGEMA_signal_29745), .Q (new_AGEMA_signal_29746) ) ;
    buf_clk new_AGEMA_reg_buffer_8793 ( .C (clk), .D (new_AGEMA_signal_29748), .Q (new_AGEMA_signal_29749) ) ;
    buf_clk new_AGEMA_reg_buffer_8796 ( .C (clk), .D (new_AGEMA_signal_29751), .Q (new_AGEMA_signal_29752) ) ;
    buf_clk new_AGEMA_reg_buffer_8799 ( .C (clk), .D (new_AGEMA_signal_29754), .Q (new_AGEMA_signal_29755) ) ;
    buf_clk new_AGEMA_reg_buffer_8802 ( .C (clk), .D (new_AGEMA_signal_29757), .Q (new_AGEMA_signal_29758) ) ;
    buf_clk new_AGEMA_reg_buffer_8805 ( .C (clk), .D (new_AGEMA_signal_29760), .Q (new_AGEMA_signal_29761) ) ;
    buf_clk new_AGEMA_reg_buffer_8808 ( .C (clk), .D (new_AGEMA_signal_29763), .Q (new_AGEMA_signal_29764) ) ;
    buf_clk new_AGEMA_reg_buffer_8811 ( .C (clk), .D (new_AGEMA_signal_29766), .Q (new_AGEMA_signal_29767) ) ;
    buf_clk new_AGEMA_reg_buffer_8814 ( .C (clk), .D (new_AGEMA_signal_29769), .Q (new_AGEMA_signal_29770) ) ;
    buf_clk new_AGEMA_reg_buffer_8817 ( .C (clk), .D (new_AGEMA_signal_29772), .Q (new_AGEMA_signal_29773) ) ;
    buf_clk new_AGEMA_reg_buffer_8820 ( .C (clk), .D (new_AGEMA_signal_29775), .Q (new_AGEMA_signal_29776) ) ;
    buf_clk new_AGEMA_reg_buffer_8823 ( .C (clk), .D (new_AGEMA_signal_29778), .Q (new_AGEMA_signal_29779) ) ;
    buf_clk new_AGEMA_reg_buffer_8826 ( .C (clk), .D (new_AGEMA_signal_29781), .Q (new_AGEMA_signal_29782) ) ;
    buf_clk new_AGEMA_reg_buffer_8829 ( .C (clk), .D (new_AGEMA_signal_29784), .Q (new_AGEMA_signal_29785) ) ;
    buf_clk new_AGEMA_reg_buffer_8832 ( .C (clk), .D (new_AGEMA_signal_29787), .Q (new_AGEMA_signal_29788) ) ;
    buf_clk new_AGEMA_reg_buffer_8835 ( .C (clk), .D (new_AGEMA_signal_29790), .Q (new_AGEMA_signal_29791) ) ;
    buf_clk new_AGEMA_reg_buffer_8838 ( .C (clk), .D (new_AGEMA_signal_29793), .Q (new_AGEMA_signal_29794) ) ;
    buf_clk new_AGEMA_reg_buffer_8841 ( .C (clk), .D (new_AGEMA_signal_29796), .Q (new_AGEMA_signal_29797) ) ;
    buf_clk new_AGEMA_reg_buffer_8844 ( .C (clk), .D (new_AGEMA_signal_29799), .Q (new_AGEMA_signal_29800) ) ;
    buf_clk new_AGEMA_reg_buffer_8847 ( .C (clk), .D (new_AGEMA_signal_29802), .Q (new_AGEMA_signal_29803) ) ;
    buf_clk new_AGEMA_reg_buffer_8850 ( .C (clk), .D (new_AGEMA_signal_29805), .Q (new_AGEMA_signal_29806) ) ;
    buf_clk new_AGEMA_reg_buffer_8853 ( .C (clk), .D (new_AGEMA_signal_29808), .Q (new_AGEMA_signal_29809) ) ;
    buf_clk new_AGEMA_reg_buffer_8856 ( .C (clk), .D (new_AGEMA_signal_29811), .Q (new_AGEMA_signal_29812) ) ;
    buf_clk new_AGEMA_reg_buffer_8859 ( .C (clk), .D (new_AGEMA_signal_29814), .Q (new_AGEMA_signal_29815) ) ;
    buf_clk new_AGEMA_reg_buffer_8862 ( .C (clk), .D (new_AGEMA_signal_29817), .Q (new_AGEMA_signal_29818) ) ;
    buf_clk new_AGEMA_reg_buffer_8865 ( .C (clk), .D (new_AGEMA_signal_29820), .Q (new_AGEMA_signal_29821) ) ;
    buf_clk new_AGEMA_reg_buffer_8868 ( .C (clk), .D (new_AGEMA_signal_29823), .Q (new_AGEMA_signal_29824) ) ;
    buf_clk new_AGEMA_reg_buffer_8871 ( .C (clk), .D (new_AGEMA_signal_29826), .Q (new_AGEMA_signal_29827) ) ;
    buf_clk new_AGEMA_reg_buffer_8874 ( .C (clk), .D (new_AGEMA_signal_29829), .Q (new_AGEMA_signal_29830) ) ;
    buf_clk new_AGEMA_reg_buffer_8877 ( .C (clk), .D (new_AGEMA_signal_29832), .Q (new_AGEMA_signal_29833) ) ;
    buf_clk new_AGEMA_reg_buffer_8880 ( .C (clk), .D (new_AGEMA_signal_29835), .Q (new_AGEMA_signal_29836) ) ;
    buf_clk new_AGEMA_reg_buffer_8883 ( .C (clk), .D (new_AGEMA_signal_29838), .Q (new_AGEMA_signal_29839) ) ;
    buf_clk new_AGEMA_reg_buffer_8886 ( .C (clk), .D (new_AGEMA_signal_29841), .Q (new_AGEMA_signal_29842) ) ;
    buf_clk new_AGEMA_reg_buffer_8889 ( .C (clk), .D (new_AGEMA_signal_29844), .Q (new_AGEMA_signal_29845) ) ;
    buf_clk new_AGEMA_reg_buffer_8892 ( .C (clk), .D (new_AGEMA_signal_29847), .Q (new_AGEMA_signal_29848) ) ;
    buf_clk new_AGEMA_reg_buffer_8895 ( .C (clk), .D (new_AGEMA_signal_29850), .Q (new_AGEMA_signal_29851) ) ;
    buf_clk new_AGEMA_reg_buffer_8898 ( .C (clk), .D (new_AGEMA_signal_29853), .Q (new_AGEMA_signal_29854) ) ;
    buf_clk new_AGEMA_reg_buffer_8901 ( .C (clk), .D (new_AGEMA_signal_29856), .Q (new_AGEMA_signal_29857) ) ;
    buf_clk new_AGEMA_reg_buffer_8904 ( .C (clk), .D (new_AGEMA_signal_29859), .Q (new_AGEMA_signal_29860) ) ;
    buf_clk new_AGEMA_reg_buffer_8907 ( .C (clk), .D (new_AGEMA_signal_29862), .Q (new_AGEMA_signal_29863) ) ;
    buf_clk new_AGEMA_reg_buffer_8910 ( .C (clk), .D (new_AGEMA_signal_29865), .Q (new_AGEMA_signal_29866) ) ;
    buf_clk new_AGEMA_reg_buffer_8913 ( .C (clk), .D (new_AGEMA_signal_29868), .Q (new_AGEMA_signal_29869) ) ;
    buf_clk new_AGEMA_reg_buffer_8916 ( .C (clk), .D (new_AGEMA_signal_29871), .Q (new_AGEMA_signal_29872) ) ;
    buf_clk new_AGEMA_reg_buffer_8919 ( .C (clk), .D (new_AGEMA_signal_29874), .Q (new_AGEMA_signal_29875) ) ;
    buf_clk new_AGEMA_reg_buffer_8922 ( .C (clk), .D (new_AGEMA_signal_29877), .Q (new_AGEMA_signal_29878) ) ;
    buf_clk new_AGEMA_reg_buffer_8925 ( .C (clk), .D (new_AGEMA_signal_29880), .Q (new_AGEMA_signal_29881) ) ;
    buf_clk new_AGEMA_reg_buffer_8928 ( .C (clk), .D (new_AGEMA_signal_29883), .Q (new_AGEMA_signal_29884) ) ;
    buf_clk new_AGEMA_reg_buffer_8931 ( .C (clk), .D (new_AGEMA_signal_29886), .Q (new_AGEMA_signal_29887) ) ;
    buf_clk new_AGEMA_reg_buffer_8934 ( .C (clk), .D (new_AGEMA_signal_29889), .Q (new_AGEMA_signal_29890) ) ;
    buf_clk new_AGEMA_reg_buffer_8937 ( .C (clk), .D (new_AGEMA_signal_29892), .Q (new_AGEMA_signal_29893) ) ;
    buf_clk new_AGEMA_reg_buffer_8940 ( .C (clk), .D (new_AGEMA_signal_29895), .Q (new_AGEMA_signal_29896) ) ;
    buf_clk new_AGEMA_reg_buffer_8943 ( .C (clk), .D (new_AGEMA_signal_29898), .Q (new_AGEMA_signal_29899) ) ;
    buf_clk new_AGEMA_reg_buffer_8946 ( .C (clk), .D (new_AGEMA_signal_29901), .Q (new_AGEMA_signal_29902) ) ;
    buf_clk new_AGEMA_reg_buffer_8949 ( .C (clk), .D (new_AGEMA_signal_29904), .Q (new_AGEMA_signal_29905) ) ;
    buf_clk new_AGEMA_reg_buffer_8952 ( .C (clk), .D (new_AGEMA_signal_29907), .Q (new_AGEMA_signal_29908) ) ;
    buf_clk new_AGEMA_reg_buffer_8955 ( .C (clk), .D (new_AGEMA_signal_29910), .Q (new_AGEMA_signal_29911) ) ;
    buf_clk new_AGEMA_reg_buffer_8958 ( .C (clk), .D (new_AGEMA_signal_29913), .Q (new_AGEMA_signal_29914) ) ;
    buf_clk new_AGEMA_reg_buffer_8961 ( .C (clk), .D (new_AGEMA_signal_29916), .Q (new_AGEMA_signal_29917) ) ;
    buf_clk new_AGEMA_reg_buffer_8964 ( .C (clk), .D (new_AGEMA_signal_29919), .Q (new_AGEMA_signal_29920) ) ;
    buf_clk new_AGEMA_reg_buffer_8967 ( .C (clk), .D (new_AGEMA_signal_29922), .Q (new_AGEMA_signal_29923) ) ;
    buf_clk new_AGEMA_reg_buffer_8970 ( .C (clk), .D (new_AGEMA_signal_29925), .Q (new_AGEMA_signal_29926) ) ;
    buf_clk new_AGEMA_reg_buffer_8973 ( .C (clk), .D (new_AGEMA_signal_29928), .Q (new_AGEMA_signal_29929) ) ;
    buf_clk new_AGEMA_reg_buffer_8976 ( .C (clk), .D (new_AGEMA_signal_29931), .Q (new_AGEMA_signal_29932) ) ;
    buf_clk new_AGEMA_reg_buffer_8979 ( .C (clk), .D (new_AGEMA_signal_29934), .Q (new_AGEMA_signal_29935) ) ;
    buf_clk new_AGEMA_reg_buffer_8982 ( .C (clk), .D (new_AGEMA_signal_29937), .Q (new_AGEMA_signal_29938) ) ;
    buf_clk new_AGEMA_reg_buffer_8985 ( .C (clk), .D (new_AGEMA_signal_29940), .Q (new_AGEMA_signal_29941) ) ;
    buf_clk new_AGEMA_reg_buffer_8988 ( .C (clk), .D (new_AGEMA_signal_29943), .Q (new_AGEMA_signal_29944) ) ;
    buf_clk new_AGEMA_reg_buffer_8991 ( .C (clk), .D (new_AGEMA_signal_29946), .Q (new_AGEMA_signal_29947) ) ;
    buf_clk new_AGEMA_reg_buffer_8994 ( .C (clk), .D (new_AGEMA_signal_29949), .Q (new_AGEMA_signal_29950) ) ;
    buf_clk new_AGEMA_reg_buffer_8997 ( .C (clk), .D (new_AGEMA_signal_29952), .Q (new_AGEMA_signal_29953) ) ;
    buf_clk new_AGEMA_reg_buffer_9000 ( .C (clk), .D (new_AGEMA_signal_29955), .Q (new_AGEMA_signal_29956) ) ;
    buf_clk new_AGEMA_reg_buffer_9003 ( .C (clk), .D (new_AGEMA_signal_29958), .Q (new_AGEMA_signal_29959) ) ;
    buf_clk new_AGEMA_reg_buffer_9006 ( .C (clk), .D (new_AGEMA_signal_29961), .Q (new_AGEMA_signal_29962) ) ;
    buf_clk new_AGEMA_reg_buffer_9009 ( .C (clk), .D (new_AGEMA_signal_29964), .Q (new_AGEMA_signal_29965) ) ;
    buf_clk new_AGEMA_reg_buffer_9012 ( .C (clk), .D (new_AGEMA_signal_29967), .Q (new_AGEMA_signal_29968) ) ;
    buf_clk new_AGEMA_reg_buffer_9015 ( .C (clk), .D (new_AGEMA_signal_29970), .Q (new_AGEMA_signal_29971) ) ;
    buf_clk new_AGEMA_reg_buffer_9018 ( .C (clk), .D (new_AGEMA_signal_29973), .Q (new_AGEMA_signal_29974) ) ;
    buf_clk new_AGEMA_reg_buffer_9021 ( .C (clk), .D (new_AGEMA_signal_29976), .Q (new_AGEMA_signal_29977) ) ;
    buf_clk new_AGEMA_reg_buffer_9024 ( .C (clk), .D (new_AGEMA_signal_29979), .Q (new_AGEMA_signal_29980) ) ;
    buf_clk new_AGEMA_reg_buffer_9027 ( .C (clk), .D (new_AGEMA_signal_29982), .Q (new_AGEMA_signal_29983) ) ;
    buf_clk new_AGEMA_reg_buffer_9030 ( .C (clk), .D (new_AGEMA_signal_29985), .Q (new_AGEMA_signal_29986) ) ;
    buf_clk new_AGEMA_reg_buffer_9033 ( .C (clk), .D (new_AGEMA_signal_29988), .Q (new_AGEMA_signal_29989) ) ;
    buf_clk new_AGEMA_reg_buffer_9036 ( .C (clk), .D (new_AGEMA_signal_29991), .Q (new_AGEMA_signal_29992) ) ;
    buf_clk new_AGEMA_reg_buffer_9039 ( .C (clk), .D (new_AGEMA_signal_29994), .Q (new_AGEMA_signal_29995) ) ;
    buf_clk new_AGEMA_reg_buffer_9042 ( .C (clk), .D (new_AGEMA_signal_29997), .Q (new_AGEMA_signal_29998) ) ;
    buf_clk new_AGEMA_reg_buffer_9045 ( .C (clk), .D (new_AGEMA_signal_30000), .Q (new_AGEMA_signal_30001) ) ;
    buf_clk new_AGEMA_reg_buffer_9048 ( .C (clk), .D (new_AGEMA_signal_30003), .Q (new_AGEMA_signal_30004) ) ;
    buf_clk new_AGEMA_reg_buffer_9051 ( .C (clk), .D (new_AGEMA_signal_30006), .Q (new_AGEMA_signal_30007) ) ;
    buf_clk new_AGEMA_reg_buffer_9054 ( .C (clk), .D (new_AGEMA_signal_30009), .Q (new_AGEMA_signal_30010) ) ;
    buf_clk new_AGEMA_reg_buffer_9057 ( .C (clk), .D (new_AGEMA_signal_30012), .Q (new_AGEMA_signal_30013) ) ;
    buf_clk new_AGEMA_reg_buffer_9060 ( .C (clk), .D (new_AGEMA_signal_30015), .Q (new_AGEMA_signal_30016) ) ;
    buf_clk new_AGEMA_reg_buffer_9063 ( .C (clk), .D (new_AGEMA_signal_30018), .Q (new_AGEMA_signal_30019) ) ;
    buf_clk new_AGEMA_reg_buffer_9066 ( .C (clk), .D (new_AGEMA_signal_30021), .Q (new_AGEMA_signal_30022) ) ;
    buf_clk new_AGEMA_reg_buffer_9069 ( .C (clk), .D (new_AGEMA_signal_30024), .Q (new_AGEMA_signal_30025) ) ;
    buf_clk new_AGEMA_reg_buffer_9072 ( .C (clk), .D (new_AGEMA_signal_30027), .Q (new_AGEMA_signal_30028) ) ;
    buf_clk new_AGEMA_reg_buffer_9075 ( .C (clk), .D (new_AGEMA_signal_30030), .Q (new_AGEMA_signal_30031) ) ;
    buf_clk new_AGEMA_reg_buffer_9078 ( .C (clk), .D (new_AGEMA_signal_30033), .Q (new_AGEMA_signal_30034) ) ;
    buf_clk new_AGEMA_reg_buffer_9081 ( .C (clk), .D (new_AGEMA_signal_30036), .Q (new_AGEMA_signal_30037) ) ;
    buf_clk new_AGEMA_reg_buffer_9084 ( .C (clk), .D (new_AGEMA_signal_30039), .Q (new_AGEMA_signal_30040) ) ;
    buf_clk new_AGEMA_reg_buffer_9087 ( .C (clk), .D (new_AGEMA_signal_30042), .Q (new_AGEMA_signal_30043) ) ;
    buf_clk new_AGEMA_reg_buffer_9090 ( .C (clk), .D (new_AGEMA_signal_30045), .Q (new_AGEMA_signal_30046) ) ;
    buf_clk new_AGEMA_reg_buffer_9093 ( .C (clk), .D (new_AGEMA_signal_30048), .Q (new_AGEMA_signal_30049) ) ;
    buf_clk new_AGEMA_reg_buffer_9096 ( .C (clk), .D (new_AGEMA_signal_30051), .Q (new_AGEMA_signal_30052) ) ;
    buf_clk new_AGEMA_reg_buffer_9099 ( .C (clk), .D (new_AGEMA_signal_30054), .Q (new_AGEMA_signal_30055) ) ;
    buf_clk new_AGEMA_reg_buffer_9102 ( .C (clk), .D (new_AGEMA_signal_30057), .Q (new_AGEMA_signal_30058) ) ;
    buf_clk new_AGEMA_reg_buffer_9105 ( .C (clk), .D (new_AGEMA_signal_30060), .Q (new_AGEMA_signal_30061) ) ;
    buf_clk new_AGEMA_reg_buffer_9108 ( .C (clk), .D (new_AGEMA_signal_30063), .Q (new_AGEMA_signal_30064) ) ;
    buf_clk new_AGEMA_reg_buffer_9111 ( .C (clk), .D (new_AGEMA_signal_30066), .Q (new_AGEMA_signal_30067) ) ;
    buf_clk new_AGEMA_reg_buffer_9114 ( .C (clk), .D (new_AGEMA_signal_30069), .Q (new_AGEMA_signal_30070) ) ;
    buf_clk new_AGEMA_reg_buffer_9117 ( .C (clk), .D (new_AGEMA_signal_30072), .Q (new_AGEMA_signal_30073) ) ;
    buf_clk new_AGEMA_reg_buffer_9120 ( .C (clk), .D (new_AGEMA_signal_30075), .Q (new_AGEMA_signal_30076) ) ;
    buf_clk new_AGEMA_reg_buffer_9123 ( .C (clk), .D (new_AGEMA_signal_30078), .Q (new_AGEMA_signal_30079) ) ;
    buf_clk new_AGEMA_reg_buffer_9126 ( .C (clk), .D (new_AGEMA_signal_30081), .Q (new_AGEMA_signal_30082) ) ;
    buf_clk new_AGEMA_reg_buffer_9129 ( .C (clk), .D (new_AGEMA_signal_30084), .Q (new_AGEMA_signal_30085) ) ;
    buf_clk new_AGEMA_reg_buffer_9132 ( .C (clk), .D (new_AGEMA_signal_30087), .Q (new_AGEMA_signal_30088) ) ;
    buf_clk new_AGEMA_reg_buffer_9135 ( .C (clk), .D (new_AGEMA_signal_30090), .Q (new_AGEMA_signal_30091) ) ;
    buf_clk new_AGEMA_reg_buffer_9138 ( .C (clk), .D (new_AGEMA_signal_30093), .Q (new_AGEMA_signal_30094) ) ;
    buf_clk new_AGEMA_reg_buffer_9141 ( .C (clk), .D (new_AGEMA_signal_30096), .Q (new_AGEMA_signal_30097) ) ;
    buf_clk new_AGEMA_reg_buffer_9144 ( .C (clk), .D (new_AGEMA_signal_30099), .Q (new_AGEMA_signal_30100) ) ;
    buf_clk new_AGEMA_reg_buffer_9147 ( .C (clk), .D (new_AGEMA_signal_30102), .Q (new_AGEMA_signal_30103) ) ;
    buf_clk new_AGEMA_reg_buffer_9150 ( .C (clk), .D (new_AGEMA_signal_30105), .Q (new_AGEMA_signal_30106) ) ;
    buf_clk new_AGEMA_reg_buffer_9153 ( .C (clk), .D (new_AGEMA_signal_30108), .Q (new_AGEMA_signal_30109) ) ;
    buf_clk new_AGEMA_reg_buffer_9156 ( .C (clk), .D (new_AGEMA_signal_30111), .Q (new_AGEMA_signal_30112) ) ;
    buf_clk new_AGEMA_reg_buffer_9159 ( .C (clk), .D (new_AGEMA_signal_30114), .Q (new_AGEMA_signal_30115) ) ;
    buf_clk new_AGEMA_reg_buffer_9162 ( .C (clk), .D (new_AGEMA_signal_30117), .Q (new_AGEMA_signal_30118) ) ;
    buf_clk new_AGEMA_reg_buffer_9165 ( .C (clk), .D (new_AGEMA_signal_30120), .Q (new_AGEMA_signal_30121) ) ;
    buf_clk new_AGEMA_reg_buffer_9168 ( .C (clk), .D (new_AGEMA_signal_30123), .Q (new_AGEMA_signal_30124) ) ;
    buf_clk new_AGEMA_reg_buffer_9171 ( .C (clk), .D (new_AGEMA_signal_30126), .Q (new_AGEMA_signal_30127) ) ;
    buf_clk new_AGEMA_reg_buffer_9174 ( .C (clk), .D (new_AGEMA_signal_30129), .Q (new_AGEMA_signal_30130) ) ;
    buf_clk new_AGEMA_reg_buffer_9177 ( .C (clk), .D (new_AGEMA_signal_30132), .Q (new_AGEMA_signal_30133) ) ;
    buf_clk new_AGEMA_reg_buffer_9180 ( .C (clk), .D (new_AGEMA_signal_30135), .Q (new_AGEMA_signal_30136) ) ;
    buf_clk new_AGEMA_reg_buffer_9183 ( .C (clk), .D (new_AGEMA_signal_30138), .Q (new_AGEMA_signal_30139) ) ;
    buf_clk new_AGEMA_reg_buffer_9186 ( .C (clk), .D (new_AGEMA_signal_30141), .Q (new_AGEMA_signal_30142) ) ;
    buf_clk new_AGEMA_reg_buffer_9189 ( .C (clk), .D (new_AGEMA_signal_30144), .Q (new_AGEMA_signal_30145) ) ;
    buf_clk new_AGEMA_reg_buffer_9192 ( .C (clk), .D (new_AGEMA_signal_30147), .Q (new_AGEMA_signal_30148) ) ;
    buf_clk new_AGEMA_reg_buffer_9195 ( .C (clk), .D (new_AGEMA_signal_30150), .Q (new_AGEMA_signal_30151) ) ;
    buf_clk new_AGEMA_reg_buffer_9198 ( .C (clk), .D (new_AGEMA_signal_30153), .Q (new_AGEMA_signal_30154) ) ;
    buf_clk new_AGEMA_reg_buffer_9201 ( .C (clk), .D (new_AGEMA_signal_30156), .Q (new_AGEMA_signal_30157) ) ;
    buf_clk new_AGEMA_reg_buffer_9204 ( .C (clk), .D (new_AGEMA_signal_30159), .Q (new_AGEMA_signal_30160) ) ;
    buf_clk new_AGEMA_reg_buffer_9207 ( .C (clk), .D (new_AGEMA_signal_30162), .Q (new_AGEMA_signal_30163) ) ;
    buf_clk new_AGEMA_reg_buffer_9210 ( .C (clk), .D (new_AGEMA_signal_30165), .Q (new_AGEMA_signal_30166) ) ;
    buf_clk new_AGEMA_reg_buffer_9213 ( .C (clk), .D (new_AGEMA_signal_30168), .Q (new_AGEMA_signal_30169) ) ;
    buf_clk new_AGEMA_reg_buffer_9216 ( .C (clk), .D (new_AGEMA_signal_30171), .Q (new_AGEMA_signal_30172) ) ;
    buf_clk new_AGEMA_reg_buffer_9219 ( .C (clk), .D (new_AGEMA_signal_30174), .Q (new_AGEMA_signal_30175) ) ;
    buf_clk new_AGEMA_reg_buffer_9222 ( .C (clk), .D (new_AGEMA_signal_30177), .Q (new_AGEMA_signal_30178) ) ;
    buf_clk new_AGEMA_reg_buffer_9225 ( .C (clk), .D (new_AGEMA_signal_30180), .Q (new_AGEMA_signal_30181) ) ;
    buf_clk new_AGEMA_reg_buffer_9228 ( .C (clk), .D (new_AGEMA_signal_30183), .Q (new_AGEMA_signal_30184) ) ;
    buf_clk new_AGEMA_reg_buffer_9231 ( .C (clk), .D (new_AGEMA_signal_30186), .Q (new_AGEMA_signal_30187) ) ;
    buf_clk new_AGEMA_reg_buffer_9234 ( .C (clk), .D (new_AGEMA_signal_30189), .Q (new_AGEMA_signal_30190) ) ;
    buf_clk new_AGEMA_reg_buffer_9237 ( .C (clk), .D (new_AGEMA_signal_30192), .Q (new_AGEMA_signal_30193) ) ;
    buf_clk new_AGEMA_reg_buffer_9240 ( .C (clk), .D (new_AGEMA_signal_30195), .Q (new_AGEMA_signal_30196) ) ;
    buf_clk new_AGEMA_reg_buffer_9243 ( .C (clk), .D (new_AGEMA_signal_30198), .Q (new_AGEMA_signal_30199) ) ;
    buf_clk new_AGEMA_reg_buffer_9246 ( .C (clk), .D (new_AGEMA_signal_30201), .Q (new_AGEMA_signal_30202) ) ;
    buf_clk new_AGEMA_reg_buffer_9249 ( .C (clk), .D (new_AGEMA_signal_30204), .Q (new_AGEMA_signal_30205) ) ;
    buf_clk new_AGEMA_reg_buffer_9252 ( .C (clk), .D (new_AGEMA_signal_30207), .Q (new_AGEMA_signal_30208) ) ;
    buf_clk new_AGEMA_reg_buffer_9255 ( .C (clk), .D (new_AGEMA_signal_30210), .Q (new_AGEMA_signal_30211) ) ;
    buf_clk new_AGEMA_reg_buffer_9258 ( .C (clk), .D (new_AGEMA_signal_30213), .Q (new_AGEMA_signal_30214) ) ;
    buf_clk new_AGEMA_reg_buffer_9261 ( .C (clk), .D (new_AGEMA_signal_30216), .Q (new_AGEMA_signal_30217) ) ;
    buf_clk new_AGEMA_reg_buffer_9264 ( .C (clk), .D (new_AGEMA_signal_30219), .Q (new_AGEMA_signal_30220) ) ;
    buf_clk new_AGEMA_reg_buffer_9267 ( .C (clk), .D (new_AGEMA_signal_30222), .Q (new_AGEMA_signal_30223) ) ;
    buf_clk new_AGEMA_reg_buffer_9270 ( .C (clk), .D (new_AGEMA_signal_30225), .Q (new_AGEMA_signal_30226) ) ;
    buf_clk new_AGEMA_reg_buffer_9273 ( .C (clk), .D (new_AGEMA_signal_30228), .Q (new_AGEMA_signal_30229) ) ;
    buf_clk new_AGEMA_reg_buffer_9276 ( .C (clk), .D (new_AGEMA_signal_30231), .Q (new_AGEMA_signal_30232) ) ;
    buf_clk new_AGEMA_reg_buffer_9279 ( .C (clk), .D (new_AGEMA_signal_30234), .Q (new_AGEMA_signal_30235) ) ;
    buf_clk new_AGEMA_reg_buffer_9282 ( .C (clk), .D (new_AGEMA_signal_30237), .Q (new_AGEMA_signal_30238) ) ;
    buf_clk new_AGEMA_reg_buffer_9285 ( .C (clk), .D (new_AGEMA_signal_30240), .Q (new_AGEMA_signal_30241) ) ;
    buf_clk new_AGEMA_reg_buffer_9288 ( .C (clk), .D (new_AGEMA_signal_30243), .Q (new_AGEMA_signal_30244) ) ;
    buf_clk new_AGEMA_reg_buffer_9291 ( .C (clk), .D (new_AGEMA_signal_30246), .Q (new_AGEMA_signal_30247) ) ;
    buf_clk new_AGEMA_reg_buffer_9294 ( .C (clk), .D (new_AGEMA_signal_30249), .Q (new_AGEMA_signal_30250) ) ;
    buf_clk new_AGEMA_reg_buffer_9297 ( .C (clk), .D (new_AGEMA_signal_30252), .Q (new_AGEMA_signal_30253) ) ;
    buf_clk new_AGEMA_reg_buffer_9300 ( .C (clk), .D (new_AGEMA_signal_30255), .Q (new_AGEMA_signal_30256) ) ;
    buf_clk new_AGEMA_reg_buffer_9303 ( .C (clk), .D (new_AGEMA_signal_30258), .Q (new_AGEMA_signal_30259) ) ;
    buf_clk new_AGEMA_reg_buffer_9306 ( .C (clk), .D (new_AGEMA_signal_30261), .Q (new_AGEMA_signal_30262) ) ;
    buf_clk new_AGEMA_reg_buffer_9309 ( .C (clk), .D (new_AGEMA_signal_30264), .Q (new_AGEMA_signal_30265) ) ;
    buf_clk new_AGEMA_reg_buffer_9312 ( .C (clk), .D (new_AGEMA_signal_30267), .Q (new_AGEMA_signal_30268) ) ;
    buf_clk new_AGEMA_reg_buffer_9315 ( .C (clk), .D (new_AGEMA_signal_30270), .Q (new_AGEMA_signal_30271) ) ;
    buf_clk new_AGEMA_reg_buffer_9318 ( .C (clk), .D (new_AGEMA_signal_30273), .Q (new_AGEMA_signal_30274) ) ;
    buf_clk new_AGEMA_reg_buffer_9321 ( .C (clk), .D (new_AGEMA_signal_30276), .Q (new_AGEMA_signal_30277) ) ;
    buf_clk new_AGEMA_reg_buffer_9324 ( .C (clk), .D (new_AGEMA_signal_30279), .Q (new_AGEMA_signal_30280) ) ;
    buf_clk new_AGEMA_reg_buffer_9327 ( .C (clk), .D (new_AGEMA_signal_30282), .Q (new_AGEMA_signal_30283) ) ;
    buf_clk new_AGEMA_reg_buffer_9330 ( .C (clk), .D (new_AGEMA_signal_30285), .Q (new_AGEMA_signal_30286) ) ;
    buf_clk new_AGEMA_reg_buffer_9333 ( .C (clk), .D (new_AGEMA_signal_30288), .Q (new_AGEMA_signal_30289) ) ;
    buf_clk new_AGEMA_reg_buffer_9336 ( .C (clk), .D (new_AGEMA_signal_30291), .Q (new_AGEMA_signal_30292) ) ;
    buf_clk new_AGEMA_reg_buffer_9339 ( .C (clk), .D (new_AGEMA_signal_30294), .Q (new_AGEMA_signal_30295) ) ;
    buf_clk new_AGEMA_reg_buffer_9342 ( .C (clk), .D (new_AGEMA_signal_30297), .Q (new_AGEMA_signal_30298) ) ;
    buf_clk new_AGEMA_reg_buffer_9345 ( .C (clk), .D (new_AGEMA_signal_30300), .Q (new_AGEMA_signal_30301) ) ;
    buf_clk new_AGEMA_reg_buffer_9348 ( .C (clk), .D (new_AGEMA_signal_30303), .Q (new_AGEMA_signal_30304) ) ;
    buf_clk new_AGEMA_reg_buffer_9351 ( .C (clk), .D (new_AGEMA_signal_30306), .Q (new_AGEMA_signal_30307) ) ;
    buf_clk new_AGEMA_reg_buffer_9354 ( .C (clk), .D (new_AGEMA_signal_30309), .Q (new_AGEMA_signal_30310) ) ;
    buf_clk new_AGEMA_reg_buffer_9357 ( .C (clk), .D (new_AGEMA_signal_30312), .Q (new_AGEMA_signal_30313) ) ;
    buf_clk new_AGEMA_reg_buffer_9360 ( .C (clk), .D (new_AGEMA_signal_30315), .Q (new_AGEMA_signal_30316) ) ;
    buf_clk new_AGEMA_reg_buffer_9363 ( .C (clk), .D (new_AGEMA_signal_30318), .Q (new_AGEMA_signal_30319) ) ;
    buf_clk new_AGEMA_reg_buffer_9366 ( .C (clk), .D (new_AGEMA_signal_30321), .Q (new_AGEMA_signal_30322) ) ;
    buf_clk new_AGEMA_reg_buffer_9369 ( .C (clk), .D (new_AGEMA_signal_30324), .Q (new_AGEMA_signal_30325) ) ;
    buf_clk new_AGEMA_reg_buffer_9372 ( .C (clk), .D (new_AGEMA_signal_30327), .Q (new_AGEMA_signal_30328) ) ;
    buf_clk new_AGEMA_reg_buffer_9375 ( .C (clk), .D (new_AGEMA_signal_30330), .Q (new_AGEMA_signal_30331) ) ;
    buf_clk new_AGEMA_reg_buffer_9378 ( .C (clk), .D (new_AGEMA_signal_30333), .Q (new_AGEMA_signal_30334) ) ;
    buf_clk new_AGEMA_reg_buffer_9381 ( .C (clk), .D (new_AGEMA_signal_30336), .Q (new_AGEMA_signal_30337) ) ;
    buf_clk new_AGEMA_reg_buffer_9384 ( .C (clk), .D (new_AGEMA_signal_30339), .Q (new_AGEMA_signal_30340) ) ;
    buf_clk new_AGEMA_reg_buffer_9387 ( .C (clk), .D (new_AGEMA_signal_30342), .Q (new_AGEMA_signal_30343) ) ;
    buf_clk new_AGEMA_reg_buffer_9390 ( .C (clk), .D (new_AGEMA_signal_30345), .Q (new_AGEMA_signal_30346) ) ;
    buf_clk new_AGEMA_reg_buffer_9393 ( .C (clk), .D (new_AGEMA_signal_30348), .Q (new_AGEMA_signal_30349) ) ;
    buf_clk new_AGEMA_reg_buffer_9396 ( .C (clk), .D (new_AGEMA_signal_30351), .Q (new_AGEMA_signal_30352) ) ;
    buf_clk new_AGEMA_reg_buffer_9399 ( .C (clk), .D (new_AGEMA_signal_30354), .Q (new_AGEMA_signal_30355) ) ;
    buf_clk new_AGEMA_reg_buffer_9402 ( .C (clk), .D (new_AGEMA_signal_30357), .Q (new_AGEMA_signal_30358) ) ;
    buf_clk new_AGEMA_reg_buffer_9405 ( .C (clk), .D (new_AGEMA_signal_30360), .Q (new_AGEMA_signal_30361) ) ;
    buf_clk new_AGEMA_reg_buffer_9408 ( .C (clk), .D (new_AGEMA_signal_30363), .Q (new_AGEMA_signal_30364) ) ;
    buf_clk new_AGEMA_reg_buffer_9411 ( .C (clk), .D (new_AGEMA_signal_30366), .Q (new_AGEMA_signal_30367) ) ;
    buf_clk new_AGEMA_reg_buffer_9414 ( .C (clk), .D (new_AGEMA_signal_30369), .Q (new_AGEMA_signal_30370) ) ;
    buf_clk new_AGEMA_reg_buffer_9417 ( .C (clk), .D (new_AGEMA_signal_30372), .Q (new_AGEMA_signal_30373) ) ;
    buf_clk new_AGEMA_reg_buffer_9420 ( .C (clk), .D (new_AGEMA_signal_30375), .Q (new_AGEMA_signal_30376) ) ;
    buf_clk new_AGEMA_reg_buffer_9423 ( .C (clk), .D (new_AGEMA_signal_30378), .Q (new_AGEMA_signal_30379) ) ;
    buf_clk new_AGEMA_reg_buffer_9426 ( .C (clk), .D (new_AGEMA_signal_30381), .Q (new_AGEMA_signal_30382) ) ;
    buf_clk new_AGEMA_reg_buffer_9429 ( .C (clk), .D (new_AGEMA_signal_30384), .Q (new_AGEMA_signal_30385) ) ;
    buf_clk new_AGEMA_reg_buffer_9432 ( .C (clk), .D (new_AGEMA_signal_30387), .Q (new_AGEMA_signal_30388) ) ;
    buf_clk new_AGEMA_reg_buffer_9435 ( .C (clk), .D (new_AGEMA_signal_30390), .Q (new_AGEMA_signal_30391) ) ;
    buf_clk new_AGEMA_reg_buffer_9438 ( .C (clk), .D (new_AGEMA_signal_30393), .Q (new_AGEMA_signal_30394) ) ;
    buf_clk new_AGEMA_reg_buffer_9441 ( .C (clk), .D (new_AGEMA_signal_30396), .Q (new_AGEMA_signal_30397) ) ;
    buf_clk new_AGEMA_reg_buffer_9444 ( .C (clk), .D (new_AGEMA_signal_30399), .Q (new_AGEMA_signal_30400) ) ;
    buf_clk new_AGEMA_reg_buffer_9447 ( .C (clk), .D (new_AGEMA_signal_30402), .Q (new_AGEMA_signal_30403) ) ;
    buf_clk new_AGEMA_reg_buffer_9450 ( .C (clk), .D (new_AGEMA_signal_30405), .Q (new_AGEMA_signal_30406) ) ;
    buf_clk new_AGEMA_reg_buffer_9453 ( .C (clk), .D (new_AGEMA_signal_30408), .Q (new_AGEMA_signal_30409) ) ;
    buf_clk new_AGEMA_reg_buffer_9456 ( .C (clk), .D (new_AGEMA_signal_30411), .Q (new_AGEMA_signal_30412) ) ;
    buf_clk new_AGEMA_reg_buffer_9459 ( .C (clk), .D (new_AGEMA_signal_30414), .Q (new_AGEMA_signal_30415) ) ;
    buf_clk new_AGEMA_reg_buffer_9462 ( .C (clk), .D (new_AGEMA_signal_30417), .Q (new_AGEMA_signal_30418) ) ;
    buf_clk new_AGEMA_reg_buffer_9465 ( .C (clk), .D (new_AGEMA_signal_30420), .Q (new_AGEMA_signal_30421) ) ;
    buf_clk new_AGEMA_reg_buffer_9468 ( .C (clk), .D (new_AGEMA_signal_30423), .Q (new_AGEMA_signal_30424) ) ;
    buf_clk new_AGEMA_reg_buffer_9471 ( .C (clk), .D (new_AGEMA_signal_30426), .Q (new_AGEMA_signal_30427) ) ;
    buf_clk new_AGEMA_reg_buffer_9474 ( .C (clk), .D (new_AGEMA_signal_30429), .Q (new_AGEMA_signal_30430) ) ;
    buf_clk new_AGEMA_reg_buffer_9477 ( .C (clk), .D (new_AGEMA_signal_30432), .Q (new_AGEMA_signal_30433) ) ;
    buf_clk new_AGEMA_reg_buffer_9480 ( .C (clk), .D (new_AGEMA_signal_30435), .Q (new_AGEMA_signal_30436) ) ;
    buf_clk new_AGEMA_reg_buffer_9483 ( .C (clk), .D (new_AGEMA_signal_30438), .Q (new_AGEMA_signal_30439) ) ;
    buf_clk new_AGEMA_reg_buffer_9486 ( .C (clk), .D (new_AGEMA_signal_30441), .Q (new_AGEMA_signal_30442) ) ;
    buf_clk new_AGEMA_reg_buffer_9489 ( .C (clk), .D (new_AGEMA_signal_30444), .Q (new_AGEMA_signal_30445) ) ;
    buf_clk new_AGEMA_reg_buffer_9492 ( .C (clk), .D (new_AGEMA_signal_30447), .Q (new_AGEMA_signal_30448) ) ;
    buf_clk new_AGEMA_reg_buffer_9495 ( .C (clk), .D (new_AGEMA_signal_30450), .Q (new_AGEMA_signal_30451) ) ;
    buf_clk new_AGEMA_reg_buffer_9498 ( .C (clk), .D (new_AGEMA_signal_30453), .Q (new_AGEMA_signal_30454) ) ;
    buf_clk new_AGEMA_reg_buffer_9501 ( .C (clk), .D (new_AGEMA_signal_30456), .Q (new_AGEMA_signal_30457) ) ;
    buf_clk new_AGEMA_reg_buffer_9504 ( .C (clk), .D (new_AGEMA_signal_30459), .Q (new_AGEMA_signal_30460) ) ;
    buf_clk new_AGEMA_reg_buffer_9507 ( .C (clk), .D (new_AGEMA_signal_30462), .Q (new_AGEMA_signal_30463) ) ;
    buf_clk new_AGEMA_reg_buffer_9510 ( .C (clk), .D (new_AGEMA_signal_30465), .Q (new_AGEMA_signal_30466) ) ;
    buf_clk new_AGEMA_reg_buffer_9513 ( .C (clk), .D (new_AGEMA_signal_30468), .Q (new_AGEMA_signal_30469) ) ;
    buf_clk new_AGEMA_reg_buffer_9516 ( .C (clk), .D (new_AGEMA_signal_30471), .Q (new_AGEMA_signal_30472) ) ;
    buf_clk new_AGEMA_reg_buffer_9519 ( .C (clk), .D (new_AGEMA_signal_30474), .Q (new_AGEMA_signal_30475) ) ;
    buf_clk new_AGEMA_reg_buffer_9522 ( .C (clk), .D (new_AGEMA_signal_30477), .Q (new_AGEMA_signal_30478) ) ;
    buf_clk new_AGEMA_reg_buffer_9525 ( .C (clk), .D (new_AGEMA_signal_30480), .Q (new_AGEMA_signal_30481) ) ;
    buf_clk new_AGEMA_reg_buffer_9528 ( .C (clk), .D (new_AGEMA_signal_30483), .Q (new_AGEMA_signal_30484) ) ;
    buf_clk new_AGEMA_reg_buffer_9531 ( .C (clk), .D (new_AGEMA_signal_30486), .Q (new_AGEMA_signal_30487) ) ;
    buf_clk new_AGEMA_reg_buffer_9534 ( .C (clk), .D (new_AGEMA_signal_30489), .Q (new_AGEMA_signal_30490) ) ;
    buf_clk new_AGEMA_reg_buffer_9537 ( .C (clk), .D (new_AGEMA_signal_30492), .Q (new_AGEMA_signal_30493) ) ;
    buf_clk new_AGEMA_reg_buffer_9540 ( .C (clk), .D (new_AGEMA_signal_30495), .Q (new_AGEMA_signal_30496) ) ;
    buf_clk new_AGEMA_reg_buffer_9543 ( .C (clk), .D (new_AGEMA_signal_30498), .Q (new_AGEMA_signal_30499) ) ;
    buf_clk new_AGEMA_reg_buffer_9546 ( .C (clk), .D (new_AGEMA_signal_30501), .Q (new_AGEMA_signal_30502) ) ;
    buf_clk new_AGEMA_reg_buffer_9549 ( .C (clk), .D (new_AGEMA_signal_30504), .Q (new_AGEMA_signal_30505) ) ;
    buf_clk new_AGEMA_reg_buffer_9552 ( .C (clk), .D (new_AGEMA_signal_30507), .Q (new_AGEMA_signal_30508) ) ;
    buf_clk new_AGEMA_reg_buffer_9555 ( .C (clk), .D (new_AGEMA_signal_30510), .Q (new_AGEMA_signal_30511) ) ;
    buf_clk new_AGEMA_reg_buffer_9558 ( .C (clk), .D (new_AGEMA_signal_30513), .Q (new_AGEMA_signal_30514) ) ;
    buf_clk new_AGEMA_reg_buffer_9561 ( .C (clk), .D (new_AGEMA_signal_30516), .Q (new_AGEMA_signal_30517) ) ;
    buf_clk new_AGEMA_reg_buffer_9564 ( .C (clk), .D (new_AGEMA_signal_30519), .Q (new_AGEMA_signal_30520) ) ;
    buf_clk new_AGEMA_reg_buffer_9567 ( .C (clk), .D (new_AGEMA_signal_30522), .Q (new_AGEMA_signal_30523) ) ;
    buf_clk new_AGEMA_reg_buffer_9570 ( .C (clk), .D (new_AGEMA_signal_30525), .Q (new_AGEMA_signal_30526) ) ;
    buf_clk new_AGEMA_reg_buffer_9573 ( .C (clk), .D (new_AGEMA_signal_30528), .Q (new_AGEMA_signal_30529) ) ;
    buf_clk new_AGEMA_reg_buffer_9576 ( .C (clk), .D (new_AGEMA_signal_30531), .Q (new_AGEMA_signal_30532) ) ;
    buf_clk new_AGEMA_reg_buffer_9579 ( .C (clk), .D (new_AGEMA_signal_30534), .Q (new_AGEMA_signal_30535) ) ;
    buf_clk new_AGEMA_reg_buffer_9582 ( .C (clk), .D (new_AGEMA_signal_30537), .Q (new_AGEMA_signal_30538) ) ;
    buf_clk new_AGEMA_reg_buffer_9585 ( .C (clk), .D (new_AGEMA_signal_30540), .Q (new_AGEMA_signal_30541) ) ;
    buf_clk new_AGEMA_reg_buffer_9588 ( .C (clk), .D (new_AGEMA_signal_30543), .Q (new_AGEMA_signal_30544) ) ;
    buf_clk new_AGEMA_reg_buffer_9591 ( .C (clk), .D (new_AGEMA_signal_30546), .Q (new_AGEMA_signal_30547) ) ;
    buf_clk new_AGEMA_reg_buffer_9594 ( .C (clk), .D (new_AGEMA_signal_30549), .Q (new_AGEMA_signal_30550) ) ;
    buf_clk new_AGEMA_reg_buffer_9597 ( .C (clk), .D (new_AGEMA_signal_30552), .Q (new_AGEMA_signal_30553) ) ;
    buf_clk new_AGEMA_reg_buffer_9600 ( .C (clk), .D (new_AGEMA_signal_30555), .Q (new_AGEMA_signal_30556) ) ;
    buf_clk new_AGEMA_reg_buffer_9603 ( .C (clk), .D (new_AGEMA_signal_30558), .Q (new_AGEMA_signal_30559) ) ;
    buf_clk new_AGEMA_reg_buffer_9606 ( .C (clk), .D (new_AGEMA_signal_30561), .Q (new_AGEMA_signal_30562) ) ;
    buf_clk new_AGEMA_reg_buffer_9609 ( .C (clk), .D (new_AGEMA_signal_30564), .Q (new_AGEMA_signal_30565) ) ;
    buf_clk new_AGEMA_reg_buffer_9612 ( .C (clk), .D (new_AGEMA_signal_30567), .Q (new_AGEMA_signal_30568) ) ;
    buf_clk new_AGEMA_reg_buffer_9615 ( .C (clk), .D (new_AGEMA_signal_30570), .Q (new_AGEMA_signal_30571) ) ;
    buf_clk new_AGEMA_reg_buffer_9618 ( .C (clk), .D (new_AGEMA_signal_30573), .Q (new_AGEMA_signal_30574) ) ;
    buf_clk new_AGEMA_reg_buffer_9621 ( .C (clk), .D (new_AGEMA_signal_30576), .Q (new_AGEMA_signal_30577) ) ;
    buf_clk new_AGEMA_reg_buffer_9624 ( .C (clk), .D (new_AGEMA_signal_30579), .Q (new_AGEMA_signal_30580) ) ;
    buf_clk new_AGEMA_reg_buffer_9627 ( .C (clk), .D (new_AGEMA_signal_30582), .Q (new_AGEMA_signal_30583) ) ;
    buf_clk new_AGEMA_reg_buffer_9630 ( .C (clk), .D (new_AGEMA_signal_30585), .Q (new_AGEMA_signal_30586) ) ;
    buf_clk new_AGEMA_reg_buffer_9633 ( .C (clk), .D (new_AGEMA_signal_30588), .Q (new_AGEMA_signal_30589) ) ;
    buf_clk new_AGEMA_reg_buffer_9636 ( .C (clk), .D (new_AGEMA_signal_30591), .Q (new_AGEMA_signal_30592) ) ;
    buf_clk new_AGEMA_reg_buffer_9639 ( .C (clk), .D (new_AGEMA_signal_30594), .Q (new_AGEMA_signal_30595) ) ;
    buf_clk new_AGEMA_reg_buffer_9642 ( .C (clk), .D (new_AGEMA_signal_30597), .Q (new_AGEMA_signal_30598) ) ;
    buf_clk new_AGEMA_reg_buffer_9645 ( .C (clk), .D (new_AGEMA_signal_30600), .Q (new_AGEMA_signal_30601) ) ;
    buf_clk new_AGEMA_reg_buffer_9648 ( .C (clk), .D (new_AGEMA_signal_30603), .Q (new_AGEMA_signal_30604) ) ;
    buf_clk new_AGEMA_reg_buffer_9651 ( .C (clk), .D (new_AGEMA_signal_30606), .Q (new_AGEMA_signal_30607) ) ;
    buf_clk new_AGEMA_reg_buffer_9654 ( .C (clk), .D (new_AGEMA_signal_30609), .Q (new_AGEMA_signal_30610) ) ;
    buf_clk new_AGEMA_reg_buffer_9657 ( .C (clk), .D (new_AGEMA_signal_30612), .Q (new_AGEMA_signal_30613) ) ;
    buf_clk new_AGEMA_reg_buffer_9660 ( .C (clk), .D (new_AGEMA_signal_30615), .Q (new_AGEMA_signal_30616) ) ;
    buf_clk new_AGEMA_reg_buffer_9663 ( .C (clk), .D (new_AGEMA_signal_30618), .Q (new_AGEMA_signal_30619) ) ;
    buf_clk new_AGEMA_reg_buffer_9666 ( .C (clk), .D (new_AGEMA_signal_30621), .Q (new_AGEMA_signal_30622) ) ;
    buf_clk new_AGEMA_reg_buffer_9669 ( .C (clk), .D (new_AGEMA_signal_30624), .Q (new_AGEMA_signal_30625) ) ;
    buf_clk new_AGEMA_reg_buffer_9672 ( .C (clk), .D (new_AGEMA_signal_30627), .Q (new_AGEMA_signal_30628) ) ;
    buf_clk new_AGEMA_reg_buffer_9675 ( .C (clk), .D (new_AGEMA_signal_30630), .Q (new_AGEMA_signal_30631) ) ;
    buf_clk new_AGEMA_reg_buffer_9678 ( .C (clk), .D (new_AGEMA_signal_30633), .Q (new_AGEMA_signal_30634) ) ;
    buf_clk new_AGEMA_reg_buffer_9681 ( .C (clk), .D (new_AGEMA_signal_30636), .Q (new_AGEMA_signal_30637) ) ;
    buf_clk new_AGEMA_reg_buffer_9684 ( .C (clk), .D (new_AGEMA_signal_30639), .Q (new_AGEMA_signal_30640) ) ;
    buf_clk new_AGEMA_reg_buffer_9687 ( .C (clk), .D (new_AGEMA_signal_30642), .Q (new_AGEMA_signal_30643) ) ;
    buf_clk new_AGEMA_reg_buffer_9690 ( .C (clk), .D (new_AGEMA_signal_30645), .Q (new_AGEMA_signal_30646) ) ;
    buf_clk new_AGEMA_reg_buffer_9693 ( .C (clk), .D (new_AGEMA_signal_30648), .Q (new_AGEMA_signal_30649) ) ;
    buf_clk new_AGEMA_reg_buffer_9696 ( .C (clk), .D (new_AGEMA_signal_30651), .Q (new_AGEMA_signal_30652) ) ;
    buf_clk new_AGEMA_reg_buffer_9699 ( .C (clk), .D (new_AGEMA_signal_30654), .Q (new_AGEMA_signal_30655) ) ;
    buf_clk new_AGEMA_reg_buffer_9702 ( .C (clk), .D (new_AGEMA_signal_30657), .Q (new_AGEMA_signal_30658) ) ;
    buf_clk new_AGEMA_reg_buffer_9705 ( .C (clk), .D (new_AGEMA_signal_30660), .Q (new_AGEMA_signal_30661) ) ;
    buf_clk new_AGEMA_reg_buffer_9708 ( .C (clk), .D (new_AGEMA_signal_30663), .Q (new_AGEMA_signal_30664) ) ;
    buf_clk new_AGEMA_reg_buffer_9711 ( .C (clk), .D (new_AGEMA_signal_30666), .Q (new_AGEMA_signal_30667) ) ;
    buf_clk new_AGEMA_reg_buffer_9714 ( .C (clk), .D (new_AGEMA_signal_30669), .Q (new_AGEMA_signal_30670) ) ;
    buf_clk new_AGEMA_reg_buffer_9717 ( .C (clk), .D (new_AGEMA_signal_30672), .Q (new_AGEMA_signal_30673) ) ;
    buf_clk new_AGEMA_reg_buffer_9720 ( .C (clk), .D (new_AGEMA_signal_30675), .Q (new_AGEMA_signal_30676) ) ;
    buf_clk new_AGEMA_reg_buffer_9723 ( .C (clk), .D (new_AGEMA_signal_30678), .Q (new_AGEMA_signal_30679) ) ;
    buf_clk new_AGEMA_reg_buffer_9726 ( .C (clk), .D (new_AGEMA_signal_30681), .Q (new_AGEMA_signal_30682) ) ;
    buf_clk new_AGEMA_reg_buffer_9729 ( .C (clk), .D (new_AGEMA_signal_30684), .Q (new_AGEMA_signal_30685) ) ;
    buf_clk new_AGEMA_reg_buffer_9732 ( .C (clk), .D (new_AGEMA_signal_30687), .Q (new_AGEMA_signal_30688) ) ;
    buf_clk new_AGEMA_reg_buffer_9735 ( .C (clk), .D (new_AGEMA_signal_30690), .Q (new_AGEMA_signal_30691) ) ;
    buf_clk new_AGEMA_reg_buffer_9738 ( .C (clk), .D (new_AGEMA_signal_30693), .Q (new_AGEMA_signal_30694) ) ;
    buf_clk new_AGEMA_reg_buffer_9741 ( .C (clk), .D (new_AGEMA_signal_30696), .Q (new_AGEMA_signal_30697) ) ;
    buf_clk new_AGEMA_reg_buffer_9744 ( .C (clk), .D (new_AGEMA_signal_30699), .Q (new_AGEMA_signal_30700) ) ;
    buf_clk new_AGEMA_reg_buffer_9747 ( .C (clk), .D (new_AGEMA_signal_30702), .Q (new_AGEMA_signal_30703) ) ;
    buf_clk new_AGEMA_reg_buffer_9750 ( .C (clk), .D (new_AGEMA_signal_30705), .Q (new_AGEMA_signal_30706) ) ;
    buf_clk new_AGEMA_reg_buffer_9753 ( .C (clk), .D (new_AGEMA_signal_30708), .Q (new_AGEMA_signal_30709) ) ;
    buf_clk new_AGEMA_reg_buffer_9756 ( .C (clk), .D (new_AGEMA_signal_30711), .Q (new_AGEMA_signal_30712) ) ;
    buf_clk new_AGEMA_reg_buffer_9759 ( .C (clk), .D (new_AGEMA_signal_30714), .Q (new_AGEMA_signal_30715) ) ;
    buf_clk new_AGEMA_reg_buffer_9762 ( .C (clk), .D (new_AGEMA_signal_30717), .Q (new_AGEMA_signal_30718) ) ;
    buf_clk new_AGEMA_reg_buffer_9765 ( .C (clk), .D (new_AGEMA_signal_30720), .Q (new_AGEMA_signal_30721) ) ;
    buf_clk new_AGEMA_reg_buffer_9768 ( .C (clk), .D (new_AGEMA_signal_30723), .Q (new_AGEMA_signal_30724) ) ;
    buf_clk new_AGEMA_reg_buffer_9771 ( .C (clk), .D (new_AGEMA_signal_30726), .Q (new_AGEMA_signal_30727) ) ;
    buf_clk new_AGEMA_reg_buffer_9774 ( .C (clk), .D (new_AGEMA_signal_30729), .Q (new_AGEMA_signal_30730) ) ;
    buf_clk new_AGEMA_reg_buffer_9777 ( .C (clk), .D (new_AGEMA_signal_30732), .Q (new_AGEMA_signal_30733) ) ;
    buf_clk new_AGEMA_reg_buffer_9780 ( .C (clk), .D (new_AGEMA_signal_30735), .Q (new_AGEMA_signal_30736) ) ;
    buf_clk new_AGEMA_reg_buffer_9783 ( .C (clk), .D (new_AGEMA_signal_30738), .Q (new_AGEMA_signal_30739) ) ;
    buf_clk new_AGEMA_reg_buffer_9786 ( .C (clk), .D (new_AGEMA_signal_30741), .Q (new_AGEMA_signal_30742) ) ;
    buf_clk new_AGEMA_reg_buffer_9789 ( .C (clk), .D (new_AGEMA_signal_30744), .Q (new_AGEMA_signal_30745) ) ;
    buf_clk new_AGEMA_reg_buffer_9792 ( .C (clk), .D (new_AGEMA_signal_30747), .Q (new_AGEMA_signal_30748) ) ;
    buf_clk new_AGEMA_reg_buffer_9795 ( .C (clk), .D (new_AGEMA_signal_30750), .Q (new_AGEMA_signal_30751) ) ;
    buf_clk new_AGEMA_reg_buffer_9798 ( .C (clk), .D (new_AGEMA_signal_30753), .Q (new_AGEMA_signal_30754) ) ;
    buf_clk new_AGEMA_reg_buffer_9801 ( .C (clk), .D (new_AGEMA_signal_30756), .Q (new_AGEMA_signal_30757) ) ;
    buf_clk new_AGEMA_reg_buffer_9804 ( .C (clk), .D (new_AGEMA_signal_30759), .Q (new_AGEMA_signal_30760) ) ;
    buf_clk new_AGEMA_reg_buffer_9807 ( .C (clk), .D (new_AGEMA_signal_30762), .Q (new_AGEMA_signal_30763) ) ;
    buf_clk new_AGEMA_reg_buffer_9810 ( .C (clk), .D (new_AGEMA_signal_30765), .Q (new_AGEMA_signal_30766) ) ;
    buf_clk new_AGEMA_reg_buffer_9813 ( .C (clk), .D (new_AGEMA_signal_30768), .Q (new_AGEMA_signal_30769) ) ;
    buf_clk new_AGEMA_reg_buffer_9816 ( .C (clk), .D (new_AGEMA_signal_30771), .Q (new_AGEMA_signal_30772) ) ;
    buf_clk new_AGEMA_reg_buffer_9819 ( .C (clk), .D (new_AGEMA_signal_30774), .Q (new_AGEMA_signal_30775) ) ;
    buf_clk new_AGEMA_reg_buffer_9822 ( .C (clk), .D (new_AGEMA_signal_30777), .Q (new_AGEMA_signal_30778) ) ;
    buf_clk new_AGEMA_reg_buffer_9825 ( .C (clk), .D (new_AGEMA_signal_30780), .Q (new_AGEMA_signal_30781) ) ;
    buf_clk new_AGEMA_reg_buffer_9828 ( .C (clk), .D (new_AGEMA_signal_30783), .Q (new_AGEMA_signal_30784) ) ;
    buf_clk new_AGEMA_reg_buffer_9831 ( .C (clk), .D (new_AGEMA_signal_30786), .Q (new_AGEMA_signal_30787) ) ;
    buf_clk new_AGEMA_reg_buffer_9834 ( .C (clk), .D (new_AGEMA_signal_30789), .Q (new_AGEMA_signal_30790) ) ;
    buf_clk new_AGEMA_reg_buffer_9837 ( .C (clk), .D (new_AGEMA_signal_30792), .Q (new_AGEMA_signal_30793) ) ;
    buf_clk new_AGEMA_reg_buffer_9840 ( .C (clk), .D (new_AGEMA_signal_30795), .Q (new_AGEMA_signal_30796) ) ;
    buf_clk new_AGEMA_reg_buffer_9843 ( .C (clk), .D (new_AGEMA_signal_30798), .Q (new_AGEMA_signal_30799) ) ;
    buf_clk new_AGEMA_reg_buffer_9846 ( .C (clk), .D (new_AGEMA_signal_30801), .Q (new_AGEMA_signal_30802) ) ;
    buf_clk new_AGEMA_reg_buffer_9849 ( .C (clk), .D (new_AGEMA_signal_30804), .Q (new_AGEMA_signal_30805) ) ;
    buf_clk new_AGEMA_reg_buffer_9852 ( .C (clk), .D (new_AGEMA_signal_30807), .Q (new_AGEMA_signal_30808) ) ;
    buf_clk new_AGEMA_reg_buffer_9855 ( .C (clk), .D (new_AGEMA_signal_30810), .Q (new_AGEMA_signal_30811) ) ;
    buf_clk new_AGEMA_reg_buffer_9858 ( .C (clk), .D (new_AGEMA_signal_30813), .Q (new_AGEMA_signal_30814) ) ;
    buf_clk new_AGEMA_reg_buffer_9861 ( .C (clk), .D (new_AGEMA_signal_30816), .Q (new_AGEMA_signal_30817) ) ;
    buf_clk new_AGEMA_reg_buffer_9864 ( .C (clk), .D (new_AGEMA_signal_30819), .Q (new_AGEMA_signal_30820) ) ;
    buf_clk new_AGEMA_reg_buffer_9867 ( .C (clk), .D (new_AGEMA_signal_30822), .Q (new_AGEMA_signal_30823) ) ;
    buf_clk new_AGEMA_reg_buffer_9870 ( .C (clk), .D (new_AGEMA_signal_30825), .Q (new_AGEMA_signal_30826) ) ;
    buf_clk new_AGEMA_reg_buffer_9873 ( .C (clk), .D (new_AGEMA_signal_30828), .Q (new_AGEMA_signal_30829) ) ;
    buf_clk new_AGEMA_reg_buffer_9876 ( .C (clk), .D (new_AGEMA_signal_30831), .Q (new_AGEMA_signal_30832) ) ;
    buf_clk new_AGEMA_reg_buffer_9879 ( .C (clk), .D (new_AGEMA_signal_30834), .Q (new_AGEMA_signal_30835) ) ;
    buf_clk new_AGEMA_reg_buffer_9882 ( .C (clk), .D (new_AGEMA_signal_30837), .Q (new_AGEMA_signal_30838) ) ;
    buf_clk new_AGEMA_reg_buffer_9885 ( .C (clk), .D (new_AGEMA_signal_30840), .Q (new_AGEMA_signal_30841) ) ;
    buf_clk new_AGEMA_reg_buffer_9888 ( .C (clk), .D (new_AGEMA_signal_30843), .Q (new_AGEMA_signal_30844) ) ;
    buf_clk new_AGEMA_reg_buffer_9891 ( .C (clk), .D (new_AGEMA_signal_30846), .Q (new_AGEMA_signal_30847) ) ;
    buf_clk new_AGEMA_reg_buffer_9894 ( .C (clk), .D (new_AGEMA_signal_30849), .Q (new_AGEMA_signal_30850) ) ;
    buf_clk new_AGEMA_reg_buffer_9897 ( .C (clk), .D (new_AGEMA_signal_30852), .Q (new_AGEMA_signal_30853) ) ;
    buf_clk new_AGEMA_reg_buffer_9900 ( .C (clk), .D (new_AGEMA_signal_30855), .Q (new_AGEMA_signal_30856) ) ;
    buf_clk new_AGEMA_reg_buffer_9903 ( .C (clk), .D (new_AGEMA_signal_30858), .Q (new_AGEMA_signal_30859) ) ;
    buf_clk new_AGEMA_reg_buffer_9906 ( .C (clk), .D (new_AGEMA_signal_30861), .Q (new_AGEMA_signal_30862) ) ;
    buf_clk new_AGEMA_reg_buffer_9909 ( .C (clk), .D (new_AGEMA_signal_30864), .Q (new_AGEMA_signal_30865) ) ;
    buf_clk new_AGEMA_reg_buffer_9912 ( .C (clk), .D (new_AGEMA_signal_30867), .Q (new_AGEMA_signal_30868) ) ;
    buf_clk new_AGEMA_reg_buffer_9915 ( .C (clk), .D (new_AGEMA_signal_30870), .Q (new_AGEMA_signal_30871) ) ;
    buf_clk new_AGEMA_reg_buffer_9918 ( .C (clk), .D (new_AGEMA_signal_30873), .Q (new_AGEMA_signal_30874) ) ;
    buf_clk new_AGEMA_reg_buffer_9921 ( .C (clk), .D (new_AGEMA_signal_30876), .Q (new_AGEMA_signal_30877) ) ;
    buf_clk new_AGEMA_reg_buffer_9924 ( .C (clk), .D (new_AGEMA_signal_30879), .Q (new_AGEMA_signal_30880) ) ;
    buf_clk new_AGEMA_reg_buffer_9927 ( .C (clk), .D (new_AGEMA_signal_30882), .Q (new_AGEMA_signal_30883) ) ;
    buf_clk new_AGEMA_reg_buffer_9930 ( .C (clk), .D (new_AGEMA_signal_30885), .Q (new_AGEMA_signal_30886) ) ;
    buf_clk new_AGEMA_reg_buffer_9933 ( .C (clk), .D (new_AGEMA_signal_30888), .Q (new_AGEMA_signal_30889) ) ;
    buf_clk new_AGEMA_reg_buffer_9936 ( .C (clk), .D (new_AGEMA_signal_30891), .Q (new_AGEMA_signal_30892) ) ;
    buf_clk new_AGEMA_reg_buffer_9939 ( .C (clk), .D (new_AGEMA_signal_30894), .Q (new_AGEMA_signal_30895) ) ;
    buf_clk new_AGEMA_reg_buffer_9942 ( .C (clk), .D (new_AGEMA_signal_30897), .Q (new_AGEMA_signal_30898) ) ;
    buf_clk new_AGEMA_reg_buffer_9945 ( .C (clk), .D (new_AGEMA_signal_30900), .Q (new_AGEMA_signal_30901) ) ;
    buf_clk new_AGEMA_reg_buffer_9948 ( .C (clk), .D (new_AGEMA_signal_30903), .Q (new_AGEMA_signal_30904) ) ;
    buf_clk new_AGEMA_reg_buffer_9951 ( .C (clk), .D (new_AGEMA_signal_30906), .Q (new_AGEMA_signal_30907) ) ;
    buf_clk new_AGEMA_reg_buffer_9954 ( .C (clk), .D (new_AGEMA_signal_30909), .Q (new_AGEMA_signal_30910) ) ;
    buf_clk new_AGEMA_reg_buffer_9957 ( .C (clk), .D (new_AGEMA_signal_30912), .Q (new_AGEMA_signal_30913) ) ;
    buf_clk new_AGEMA_reg_buffer_9960 ( .C (clk), .D (new_AGEMA_signal_30915), .Q (new_AGEMA_signal_30916) ) ;
    buf_clk new_AGEMA_reg_buffer_9963 ( .C (clk), .D (new_AGEMA_signal_30918), .Q (new_AGEMA_signal_30919) ) ;
    buf_clk new_AGEMA_reg_buffer_9966 ( .C (clk), .D (new_AGEMA_signal_30921), .Q (new_AGEMA_signal_30922) ) ;
    buf_clk new_AGEMA_reg_buffer_9969 ( .C (clk), .D (new_AGEMA_signal_30924), .Q (new_AGEMA_signal_30925) ) ;
    buf_clk new_AGEMA_reg_buffer_9972 ( .C (clk), .D (new_AGEMA_signal_30927), .Q (new_AGEMA_signal_30928) ) ;
    buf_clk new_AGEMA_reg_buffer_9975 ( .C (clk), .D (new_AGEMA_signal_30930), .Q (new_AGEMA_signal_30931) ) ;
    buf_clk new_AGEMA_reg_buffer_9978 ( .C (clk), .D (new_AGEMA_signal_30933), .Q (new_AGEMA_signal_30934) ) ;
    buf_clk new_AGEMA_reg_buffer_9981 ( .C (clk), .D (new_AGEMA_signal_30936), .Q (new_AGEMA_signal_30937) ) ;
    buf_clk new_AGEMA_reg_buffer_9984 ( .C (clk), .D (new_AGEMA_signal_30939), .Q (new_AGEMA_signal_30940) ) ;
    buf_clk new_AGEMA_reg_buffer_9987 ( .C (clk), .D (new_AGEMA_signal_30942), .Q (new_AGEMA_signal_30943) ) ;
    buf_clk new_AGEMA_reg_buffer_9990 ( .C (clk), .D (new_AGEMA_signal_30945), .Q (new_AGEMA_signal_30946) ) ;
    buf_clk new_AGEMA_reg_buffer_9993 ( .C (clk), .D (new_AGEMA_signal_30948), .Q (new_AGEMA_signal_30949) ) ;
    buf_clk new_AGEMA_reg_buffer_9996 ( .C (clk), .D (new_AGEMA_signal_30951), .Q (new_AGEMA_signal_30952) ) ;
    buf_clk new_AGEMA_reg_buffer_9999 ( .C (clk), .D (new_AGEMA_signal_30954), .Q (new_AGEMA_signal_30955) ) ;
    buf_clk new_AGEMA_reg_buffer_10002 ( .C (clk), .D (new_AGEMA_signal_30957), .Q (new_AGEMA_signal_30958) ) ;
    buf_clk new_AGEMA_reg_buffer_10005 ( .C (clk), .D (new_AGEMA_signal_30960), .Q (new_AGEMA_signal_30961) ) ;
    buf_clk new_AGEMA_reg_buffer_10008 ( .C (clk), .D (new_AGEMA_signal_30963), .Q (new_AGEMA_signal_30964) ) ;
    buf_clk new_AGEMA_reg_buffer_10011 ( .C (clk), .D (new_AGEMA_signal_30966), .Q (new_AGEMA_signal_30967) ) ;
    buf_clk new_AGEMA_reg_buffer_10014 ( .C (clk), .D (new_AGEMA_signal_30969), .Q (new_AGEMA_signal_30970) ) ;
    buf_clk new_AGEMA_reg_buffer_10017 ( .C (clk), .D (new_AGEMA_signal_30972), .Q (new_AGEMA_signal_30973) ) ;
    buf_clk new_AGEMA_reg_buffer_10020 ( .C (clk), .D (new_AGEMA_signal_30975), .Q (new_AGEMA_signal_30976) ) ;
    buf_clk new_AGEMA_reg_buffer_10023 ( .C (clk), .D (new_AGEMA_signal_30978), .Q (new_AGEMA_signal_30979) ) ;
    buf_clk new_AGEMA_reg_buffer_10026 ( .C (clk), .D (new_AGEMA_signal_30981), .Q (new_AGEMA_signal_30982) ) ;
    buf_clk new_AGEMA_reg_buffer_10029 ( .C (clk), .D (new_AGEMA_signal_30984), .Q (new_AGEMA_signal_30985) ) ;
    buf_clk new_AGEMA_reg_buffer_10032 ( .C (clk), .D (new_AGEMA_signal_30987), .Q (new_AGEMA_signal_30988) ) ;
    buf_clk new_AGEMA_reg_buffer_10035 ( .C (clk), .D (new_AGEMA_signal_30990), .Q (new_AGEMA_signal_30991) ) ;
    buf_clk new_AGEMA_reg_buffer_10038 ( .C (clk), .D (new_AGEMA_signal_30993), .Q (new_AGEMA_signal_30994) ) ;
    buf_clk new_AGEMA_reg_buffer_10041 ( .C (clk), .D (new_AGEMA_signal_30996), .Q (new_AGEMA_signal_30997) ) ;
    buf_clk new_AGEMA_reg_buffer_10044 ( .C (clk), .D (new_AGEMA_signal_30999), .Q (new_AGEMA_signal_31000) ) ;
    buf_clk new_AGEMA_reg_buffer_10047 ( .C (clk), .D (new_AGEMA_signal_31002), .Q (new_AGEMA_signal_31003) ) ;
    buf_clk new_AGEMA_reg_buffer_10050 ( .C (clk), .D (new_AGEMA_signal_31005), .Q (new_AGEMA_signal_31006) ) ;
    buf_clk new_AGEMA_reg_buffer_10053 ( .C (clk), .D (new_AGEMA_signal_31008), .Q (new_AGEMA_signal_31009) ) ;
    buf_clk new_AGEMA_reg_buffer_10056 ( .C (clk), .D (new_AGEMA_signal_31011), .Q (new_AGEMA_signal_31012) ) ;
    buf_clk new_AGEMA_reg_buffer_10059 ( .C (clk), .D (new_AGEMA_signal_31014), .Q (new_AGEMA_signal_31015) ) ;
    buf_clk new_AGEMA_reg_buffer_10062 ( .C (clk), .D (new_AGEMA_signal_31017), .Q (new_AGEMA_signal_31018) ) ;
    buf_clk new_AGEMA_reg_buffer_10065 ( .C (clk), .D (new_AGEMA_signal_31020), .Q (new_AGEMA_signal_31021) ) ;
    buf_clk new_AGEMA_reg_buffer_10068 ( .C (clk), .D (new_AGEMA_signal_31023), .Q (new_AGEMA_signal_31024) ) ;
    buf_clk new_AGEMA_reg_buffer_10071 ( .C (clk), .D (new_AGEMA_signal_31026), .Q (new_AGEMA_signal_31027) ) ;
    buf_clk new_AGEMA_reg_buffer_10074 ( .C (clk), .D (new_AGEMA_signal_31029), .Q (new_AGEMA_signal_31030) ) ;
    buf_clk new_AGEMA_reg_buffer_10077 ( .C (clk), .D (new_AGEMA_signal_31032), .Q (new_AGEMA_signal_31033) ) ;
    buf_clk new_AGEMA_reg_buffer_10080 ( .C (clk), .D (new_AGEMA_signal_31035), .Q (new_AGEMA_signal_31036) ) ;
    buf_clk new_AGEMA_reg_buffer_10083 ( .C (clk), .D (new_AGEMA_signal_31038), .Q (new_AGEMA_signal_31039) ) ;
    buf_clk new_AGEMA_reg_buffer_10086 ( .C (clk), .D (new_AGEMA_signal_31041), .Q (new_AGEMA_signal_31042) ) ;
    buf_clk new_AGEMA_reg_buffer_10089 ( .C (clk), .D (new_AGEMA_signal_31044), .Q (new_AGEMA_signal_31045) ) ;
    buf_clk new_AGEMA_reg_buffer_10092 ( .C (clk), .D (new_AGEMA_signal_31047), .Q (new_AGEMA_signal_31048) ) ;
    buf_clk new_AGEMA_reg_buffer_10095 ( .C (clk), .D (new_AGEMA_signal_31050), .Q (new_AGEMA_signal_31051) ) ;
    buf_clk new_AGEMA_reg_buffer_10098 ( .C (clk), .D (new_AGEMA_signal_31053), .Q (new_AGEMA_signal_31054) ) ;
    buf_clk new_AGEMA_reg_buffer_10101 ( .C (clk), .D (new_AGEMA_signal_31056), .Q (new_AGEMA_signal_31057) ) ;
    buf_clk new_AGEMA_reg_buffer_10104 ( .C (clk), .D (new_AGEMA_signal_31059), .Q (new_AGEMA_signal_31060) ) ;
    buf_clk new_AGEMA_reg_buffer_10107 ( .C (clk), .D (new_AGEMA_signal_31062), .Q (new_AGEMA_signal_31063) ) ;
    buf_clk new_AGEMA_reg_buffer_10110 ( .C (clk), .D (new_AGEMA_signal_31065), .Q (new_AGEMA_signal_31066) ) ;
    buf_clk new_AGEMA_reg_buffer_10113 ( .C (clk), .D (new_AGEMA_signal_31068), .Q (new_AGEMA_signal_31069) ) ;
    buf_clk new_AGEMA_reg_buffer_10116 ( .C (clk), .D (new_AGEMA_signal_31071), .Q (new_AGEMA_signal_31072) ) ;
    buf_clk new_AGEMA_reg_buffer_10119 ( .C (clk), .D (new_AGEMA_signal_31074), .Q (new_AGEMA_signal_31075) ) ;
    buf_clk new_AGEMA_reg_buffer_10122 ( .C (clk), .D (new_AGEMA_signal_31077), .Q (new_AGEMA_signal_31078) ) ;
    buf_clk new_AGEMA_reg_buffer_10125 ( .C (clk), .D (new_AGEMA_signal_31080), .Q (new_AGEMA_signal_31081) ) ;
    buf_clk new_AGEMA_reg_buffer_10128 ( .C (clk), .D (new_AGEMA_signal_31083), .Q (new_AGEMA_signal_31084) ) ;
    buf_clk new_AGEMA_reg_buffer_10131 ( .C (clk), .D (new_AGEMA_signal_31086), .Q (new_AGEMA_signal_31087) ) ;
    buf_clk new_AGEMA_reg_buffer_10134 ( .C (clk), .D (new_AGEMA_signal_31089), .Q (new_AGEMA_signal_31090) ) ;
    buf_clk new_AGEMA_reg_buffer_10137 ( .C (clk), .D (new_AGEMA_signal_31092), .Q (new_AGEMA_signal_31093) ) ;
    buf_clk new_AGEMA_reg_buffer_10140 ( .C (clk), .D (new_AGEMA_signal_31095), .Q (new_AGEMA_signal_31096) ) ;
    buf_clk new_AGEMA_reg_buffer_10143 ( .C (clk), .D (new_AGEMA_signal_31098), .Q (new_AGEMA_signal_31099) ) ;
    buf_clk new_AGEMA_reg_buffer_10146 ( .C (clk), .D (new_AGEMA_signal_31101), .Q (new_AGEMA_signal_31102) ) ;
    buf_clk new_AGEMA_reg_buffer_10149 ( .C (clk), .D (new_AGEMA_signal_31104), .Q (new_AGEMA_signal_31105) ) ;
    buf_clk new_AGEMA_reg_buffer_10152 ( .C (clk), .D (new_AGEMA_signal_31107), .Q (new_AGEMA_signal_31108) ) ;
    buf_clk new_AGEMA_reg_buffer_10155 ( .C (clk), .D (new_AGEMA_signal_31110), .Q (new_AGEMA_signal_31111) ) ;
    buf_clk new_AGEMA_reg_buffer_10158 ( .C (clk), .D (new_AGEMA_signal_31113), .Q (new_AGEMA_signal_31114) ) ;
    buf_clk new_AGEMA_reg_buffer_10161 ( .C (clk), .D (new_AGEMA_signal_31116), .Q (new_AGEMA_signal_31117) ) ;
    buf_clk new_AGEMA_reg_buffer_10164 ( .C (clk), .D (new_AGEMA_signal_31119), .Q (new_AGEMA_signal_31120) ) ;
    buf_clk new_AGEMA_reg_buffer_10167 ( .C (clk), .D (new_AGEMA_signal_31122), .Q (new_AGEMA_signal_31123) ) ;
    buf_clk new_AGEMA_reg_buffer_10170 ( .C (clk), .D (new_AGEMA_signal_31125), .Q (new_AGEMA_signal_31126) ) ;
    buf_clk new_AGEMA_reg_buffer_10173 ( .C (clk), .D (new_AGEMA_signal_31128), .Q (new_AGEMA_signal_31129) ) ;
    buf_clk new_AGEMA_reg_buffer_10176 ( .C (clk), .D (new_AGEMA_signal_31131), .Q (new_AGEMA_signal_31132) ) ;
    buf_clk new_AGEMA_reg_buffer_10179 ( .C (clk), .D (new_AGEMA_signal_31134), .Q (new_AGEMA_signal_31135) ) ;
    buf_clk new_AGEMA_reg_buffer_10182 ( .C (clk), .D (new_AGEMA_signal_31137), .Q (new_AGEMA_signal_31138) ) ;
    buf_clk new_AGEMA_reg_buffer_10185 ( .C (clk), .D (new_AGEMA_signal_31140), .Q (new_AGEMA_signal_31141) ) ;
    buf_clk new_AGEMA_reg_buffer_10188 ( .C (clk), .D (new_AGEMA_signal_31143), .Q (new_AGEMA_signal_31144) ) ;
    buf_clk new_AGEMA_reg_buffer_10191 ( .C (clk), .D (new_AGEMA_signal_31146), .Q (new_AGEMA_signal_31147) ) ;
    buf_clk new_AGEMA_reg_buffer_10194 ( .C (clk), .D (new_AGEMA_signal_31149), .Q (new_AGEMA_signal_31150) ) ;
    buf_clk new_AGEMA_reg_buffer_10197 ( .C (clk), .D (new_AGEMA_signal_31152), .Q (new_AGEMA_signal_31153) ) ;
    buf_clk new_AGEMA_reg_buffer_10200 ( .C (clk), .D (new_AGEMA_signal_31155), .Q (new_AGEMA_signal_31156) ) ;
    buf_clk new_AGEMA_reg_buffer_10203 ( .C (clk), .D (new_AGEMA_signal_31158), .Q (new_AGEMA_signal_31159) ) ;
    buf_clk new_AGEMA_reg_buffer_10206 ( .C (clk), .D (new_AGEMA_signal_31161), .Q (new_AGEMA_signal_31162) ) ;
    buf_clk new_AGEMA_reg_buffer_10209 ( .C (clk), .D (new_AGEMA_signal_31164), .Q (new_AGEMA_signal_31165) ) ;
    buf_clk new_AGEMA_reg_buffer_10212 ( .C (clk), .D (new_AGEMA_signal_31167), .Q (new_AGEMA_signal_31168) ) ;
    buf_clk new_AGEMA_reg_buffer_10215 ( .C (clk), .D (new_AGEMA_signal_31170), .Q (new_AGEMA_signal_31171) ) ;
    buf_clk new_AGEMA_reg_buffer_10218 ( .C (clk), .D (new_AGEMA_signal_31173), .Q (new_AGEMA_signal_31174) ) ;
    buf_clk new_AGEMA_reg_buffer_10221 ( .C (clk), .D (new_AGEMA_signal_31176), .Q (new_AGEMA_signal_31177) ) ;
    buf_clk new_AGEMA_reg_buffer_10224 ( .C (clk), .D (new_AGEMA_signal_31179), .Q (new_AGEMA_signal_31180) ) ;
    buf_clk new_AGEMA_reg_buffer_10227 ( .C (clk), .D (new_AGEMA_signal_31182), .Q (new_AGEMA_signal_31183) ) ;
    buf_clk new_AGEMA_reg_buffer_10230 ( .C (clk), .D (new_AGEMA_signal_31185), .Q (new_AGEMA_signal_31186) ) ;
    buf_clk new_AGEMA_reg_buffer_10233 ( .C (clk), .D (new_AGEMA_signal_31188), .Q (new_AGEMA_signal_31189) ) ;
    buf_clk new_AGEMA_reg_buffer_10236 ( .C (clk), .D (new_AGEMA_signal_31191), .Q (new_AGEMA_signal_31192) ) ;
    buf_clk new_AGEMA_reg_buffer_10239 ( .C (clk), .D (new_AGEMA_signal_31194), .Q (new_AGEMA_signal_31195) ) ;
    buf_clk new_AGEMA_reg_buffer_10242 ( .C (clk), .D (new_AGEMA_signal_31197), .Q (new_AGEMA_signal_31198) ) ;
    buf_clk new_AGEMA_reg_buffer_10245 ( .C (clk), .D (new_AGEMA_signal_31200), .Q (new_AGEMA_signal_31201) ) ;
    buf_clk new_AGEMA_reg_buffer_10248 ( .C (clk), .D (new_AGEMA_signal_31203), .Q (new_AGEMA_signal_31204) ) ;
    buf_clk new_AGEMA_reg_buffer_10251 ( .C (clk), .D (new_AGEMA_signal_31206), .Q (new_AGEMA_signal_31207) ) ;
    buf_clk new_AGEMA_reg_buffer_10254 ( .C (clk), .D (new_AGEMA_signal_31209), .Q (new_AGEMA_signal_31210) ) ;
    buf_clk new_AGEMA_reg_buffer_10257 ( .C (clk), .D (new_AGEMA_signal_31212), .Q (new_AGEMA_signal_31213) ) ;
    buf_clk new_AGEMA_reg_buffer_10260 ( .C (clk), .D (new_AGEMA_signal_31215), .Q (new_AGEMA_signal_31216) ) ;
    buf_clk new_AGEMA_reg_buffer_10263 ( .C (clk), .D (new_AGEMA_signal_31218), .Q (new_AGEMA_signal_31219) ) ;
    buf_clk new_AGEMA_reg_buffer_10266 ( .C (clk), .D (new_AGEMA_signal_31221), .Q (new_AGEMA_signal_31222) ) ;
    buf_clk new_AGEMA_reg_buffer_10269 ( .C (clk), .D (new_AGEMA_signal_31224), .Q (new_AGEMA_signal_31225) ) ;
    buf_clk new_AGEMA_reg_buffer_10272 ( .C (clk), .D (new_AGEMA_signal_31227), .Q (new_AGEMA_signal_31228) ) ;
    buf_clk new_AGEMA_reg_buffer_10275 ( .C (clk), .D (new_AGEMA_signal_31230), .Q (new_AGEMA_signal_31231) ) ;
    buf_clk new_AGEMA_reg_buffer_10278 ( .C (clk), .D (new_AGEMA_signal_31233), .Q (new_AGEMA_signal_31234) ) ;
    buf_clk new_AGEMA_reg_buffer_10281 ( .C (clk), .D (new_AGEMA_signal_31236), .Q (new_AGEMA_signal_31237) ) ;
    buf_clk new_AGEMA_reg_buffer_10284 ( .C (clk), .D (new_AGEMA_signal_31239), .Q (new_AGEMA_signal_31240) ) ;
    buf_clk new_AGEMA_reg_buffer_10287 ( .C (clk), .D (new_AGEMA_signal_31242), .Q (new_AGEMA_signal_31243) ) ;
    buf_clk new_AGEMA_reg_buffer_10290 ( .C (clk), .D (new_AGEMA_signal_31245), .Q (new_AGEMA_signal_31246) ) ;
    buf_clk new_AGEMA_reg_buffer_10293 ( .C (clk), .D (new_AGEMA_signal_31248), .Q (new_AGEMA_signal_31249) ) ;
    buf_clk new_AGEMA_reg_buffer_10296 ( .C (clk), .D (new_AGEMA_signal_31251), .Q (new_AGEMA_signal_31252) ) ;
    buf_clk new_AGEMA_reg_buffer_10299 ( .C (clk), .D (new_AGEMA_signal_31254), .Q (new_AGEMA_signal_31255) ) ;
    buf_clk new_AGEMA_reg_buffer_10302 ( .C (clk), .D (new_AGEMA_signal_31257), .Q (new_AGEMA_signal_31258) ) ;
    buf_clk new_AGEMA_reg_buffer_10305 ( .C (clk), .D (new_AGEMA_signal_31260), .Q (new_AGEMA_signal_31261) ) ;
    buf_clk new_AGEMA_reg_buffer_10308 ( .C (clk), .D (new_AGEMA_signal_31263), .Q (new_AGEMA_signal_31264) ) ;
    buf_clk new_AGEMA_reg_buffer_10311 ( .C (clk), .D (new_AGEMA_signal_31266), .Q (new_AGEMA_signal_31267) ) ;
    buf_clk new_AGEMA_reg_buffer_10314 ( .C (clk), .D (new_AGEMA_signal_31269), .Q (new_AGEMA_signal_31270) ) ;
    buf_clk new_AGEMA_reg_buffer_10317 ( .C (clk), .D (new_AGEMA_signal_31272), .Q (new_AGEMA_signal_31273) ) ;
    buf_clk new_AGEMA_reg_buffer_10320 ( .C (clk), .D (new_AGEMA_signal_31275), .Q (new_AGEMA_signal_31276) ) ;
    buf_clk new_AGEMA_reg_buffer_10323 ( .C (clk), .D (new_AGEMA_signal_31278), .Q (new_AGEMA_signal_31279) ) ;
    buf_clk new_AGEMA_reg_buffer_10326 ( .C (clk), .D (new_AGEMA_signal_31281), .Q (new_AGEMA_signal_31282) ) ;
    buf_clk new_AGEMA_reg_buffer_10329 ( .C (clk), .D (new_AGEMA_signal_31284), .Q (new_AGEMA_signal_31285) ) ;
    buf_clk new_AGEMA_reg_buffer_10332 ( .C (clk), .D (new_AGEMA_signal_31287), .Q (new_AGEMA_signal_31288) ) ;
    buf_clk new_AGEMA_reg_buffer_10335 ( .C (clk), .D (new_AGEMA_signal_31290), .Q (new_AGEMA_signal_31291) ) ;
    buf_clk new_AGEMA_reg_buffer_10338 ( .C (clk), .D (new_AGEMA_signal_31293), .Q (new_AGEMA_signal_31294) ) ;
    buf_clk new_AGEMA_reg_buffer_10341 ( .C (clk), .D (new_AGEMA_signal_31296), .Q (new_AGEMA_signal_31297) ) ;
    buf_clk new_AGEMA_reg_buffer_10344 ( .C (clk), .D (new_AGEMA_signal_31299), .Q (new_AGEMA_signal_31300) ) ;
    buf_clk new_AGEMA_reg_buffer_10347 ( .C (clk), .D (new_AGEMA_signal_31302), .Q (new_AGEMA_signal_31303) ) ;
    buf_clk new_AGEMA_reg_buffer_10350 ( .C (clk), .D (new_AGEMA_signal_31305), .Q (new_AGEMA_signal_31306) ) ;
    buf_clk new_AGEMA_reg_buffer_10353 ( .C (clk), .D (new_AGEMA_signal_31308), .Q (new_AGEMA_signal_31309) ) ;
    buf_clk new_AGEMA_reg_buffer_10356 ( .C (clk), .D (new_AGEMA_signal_31311), .Q (new_AGEMA_signal_31312) ) ;
    buf_clk new_AGEMA_reg_buffer_10359 ( .C (clk), .D (new_AGEMA_signal_31314), .Q (new_AGEMA_signal_31315) ) ;
    buf_clk new_AGEMA_reg_buffer_10362 ( .C (clk), .D (new_AGEMA_signal_31317), .Q (new_AGEMA_signal_31318) ) ;
    buf_clk new_AGEMA_reg_buffer_10365 ( .C (clk), .D (new_AGEMA_signal_31320), .Q (new_AGEMA_signal_31321) ) ;
    buf_clk new_AGEMA_reg_buffer_10368 ( .C (clk), .D (new_AGEMA_signal_31323), .Q (new_AGEMA_signal_31324) ) ;
    buf_clk new_AGEMA_reg_buffer_10371 ( .C (clk), .D (new_AGEMA_signal_31326), .Q (new_AGEMA_signal_31327) ) ;
    buf_clk new_AGEMA_reg_buffer_10374 ( .C (clk), .D (new_AGEMA_signal_31329), .Q (new_AGEMA_signal_31330) ) ;
    buf_clk new_AGEMA_reg_buffer_10377 ( .C (clk), .D (new_AGEMA_signal_31332), .Q (new_AGEMA_signal_31333) ) ;
    buf_clk new_AGEMA_reg_buffer_10380 ( .C (clk), .D (new_AGEMA_signal_31335), .Q (new_AGEMA_signal_31336) ) ;
    buf_clk new_AGEMA_reg_buffer_10383 ( .C (clk), .D (new_AGEMA_signal_31338), .Q (new_AGEMA_signal_31339) ) ;
    buf_clk new_AGEMA_reg_buffer_10386 ( .C (clk), .D (new_AGEMA_signal_31341), .Q (new_AGEMA_signal_31342) ) ;
    buf_clk new_AGEMA_reg_buffer_10389 ( .C (clk), .D (new_AGEMA_signal_31344), .Q (new_AGEMA_signal_31345) ) ;
    buf_clk new_AGEMA_reg_buffer_10392 ( .C (clk), .D (new_AGEMA_signal_31347), .Q (new_AGEMA_signal_31348) ) ;
    buf_clk new_AGEMA_reg_buffer_10395 ( .C (clk), .D (new_AGEMA_signal_31350), .Q (new_AGEMA_signal_31351) ) ;
    buf_clk new_AGEMA_reg_buffer_10398 ( .C (clk), .D (new_AGEMA_signal_31353), .Q (new_AGEMA_signal_31354) ) ;
    buf_clk new_AGEMA_reg_buffer_10401 ( .C (clk), .D (new_AGEMA_signal_31356), .Q (new_AGEMA_signal_31357) ) ;
    buf_clk new_AGEMA_reg_buffer_10404 ( .C (clk), .D (new_AGEMA_signal_31359), .Q (new_AGEMA_signal_31360) ) ;
    buf_clk new_AGEMA_reg_buffer_10407 ( .C (clk), .D (new_AGEMA_signal_31362), .Q (new_AGEMA_signal_31363) ) ;
    buf_clk new_AGEMA_reg_buffer_10410 ( .C (clk), .D (new_AGEMA_signal_31365), .Q (new_AGEMA_signal_31366) ) ;
    buf_clk new_AGEMA_reg_buffer_10413 ( .C (clk), .D (new_AGEMA_signal_31368), .Q (new_AGEMA_signal_31369) ) ;
    buf_clk new_AGEMA_reg_buffer_10416 ( .C (clk), .D (new_AGEMA_signal_31371), .Q (new_AGEMA_signal_31372) ) ;
    buf_clk new_AGEMA_reg_buffer_10419 ( .C (clk), .D (new_AGEMA_signal_31374), .Q (new_AGEMA_signal_31375) ) ;
    buf_clk new_AGEMA_reg_buffer_10422 ( .C (clk), .D (new_AGEMA_signal_31377), .Q (new_AGEMA_signal_31378) ) ;
    buf_clk new_AGEMA_reg_buffer_10425 ( .C (clk), .D (new_AGEMA_signal_31380), .Q (new_AGEMA_signal_31381) ) ;
    buf_clk new_AGEMA_reg_buffer_10428 ( .C (clk), .D (new_AGEMA_signal_31383), .Q (new_AGEMA_signal_31384) ) ;
    buf_clk new_AGEMA_reg_buffer_10431 ( .C (clk), .D (new_AGEMA_signal_31386), .Q (new_AGEMA_signal_31387) ) ;
    buf_clk new_AGEMA_reg_buffer_10434 ( .C (clk), .D (new_AGEMA_signal_31389), .Q (new_AGEMA_signal_31390) ) ;
    buf_clk new_AGEMA_reg_buffer_10437 ( .C (clk), .D (new_AGEMA_signal_31392), .Q (new_AGEMA_signal_31393) ) ;
    buf_clk new_AGEMA_reg_buffer_10440 ( .C (clk), .D (new_AGEMA_signal_31395), .Q (new_AGEMA_signal_31396) ) ;
    buf_clk new_AGEMA_reg_buffer_10443 ( .C (clk), .D (new_AGEMA_signal_31398), .Q (new_AGEMA_signal_31399) ) ;
    buf_clk new_AGEMA_reg_buffer_10446 ( .C (clk), .D (new_AGEMA_signal_31401), .Q (new_AGEMA_signal_31402) ) ;
    buf_clk new_AGEMA_reg_buffer_10449 ( .C (clk), .D (new_AGEMA_signal_31404), .Q (new_AGEMA_signal_31405) ) ;
    buf_clk new_AGEMA_reg_buffer_10452 ( .C (clk), .D (new_AGEMA_signal_31407), .Q (new_AGEMA_signal_31408) ) ;
    buf_clk new_AGEMA_reg_buffer_10455 ( .C (clk), .D (new_AGEMA_signal_31410), .Q (new_AGEMA_signal_31411) ) ;
    buf_clk new_AGEMA_reg_buffer_10458 ( .C (clk), .D (new_AGEMA_signal_31413), .Q (new_AGEMA_signal_31414) ) ;
    buf_clk new_AGEMA_reg_buffer_10461 ( .C (clk), .D (new_AGEMA_signal_31416), .Q (new_AGEMA_signal_31417) ) ;
    buf_clk new_AGEMA_reg_buffer_10464 ( .C (clk), .D (new_AGEMA_signal_31419), .Q (new_AGEMA_signal_31420) ) ;
    buf_clk new_AGEMA_reg_buffer_10467 ( .C (clk), .D (new_AGEMA_signal_31422), .Q (new_AGEMA_signal_31423) ) ;
    buf_clk new_AGEMA_reg_buffer_10470 ( .C (clk), .D (new_AGEMA_signal_31425), .Q (new_AGEMA_signal_31426) ) ;
    buf_clk new_AGEMA_reg_buffer_10473 ( .C (clk), .D (new_AGEMA_signal_31428), .Q (new_AGEMA_signal_31429) ) ;
    buf_clk new_AGEMA_reg_buffer_10476 ( .C (clk), .D (new_AGEMA_signal_31431), .Q (new_AGEMA_signal_31432) ) ;
    buf_clk new_AGEMA_reg_buffer_10479 ( .C (clk), .D (new_AGEMA_signal_31434), .Q (new_AGEMA_signal_31435) ) ;
    buf_clk new_AGEMA_reg_buffer_10482 ( .C (clk), .D (new_AGEMA_signal_31437), .Q (new_AGEMA_signal_31438) ) ;
    buf_clk new_AGEMA_reg_buffer_10485 ( .C (clk), .D (new_AGEMA_signal_31440), .Q (new_AGEMA_signal_31441) ) ;
    buf_clk new_AGEMA_reg_buffer_10488 ( .C (clk), .D (new_AGEMA_signal_31443), .Q (new_AGEMA_signal_31444) ) ;
    buf_clk new_AGEMA_reg_buffer_10491 ( .C (clk), .D (new_AGEMA_signal_31446), .Q (new_AGEMA_signal_31447) ) ;
    buf_clk new_AGEMA_reg_buffer_10494 ( .C (clk), .D (new_AGEMA_signal_31449), .Q (new_AGEMA_signal_31450) ) ;
    buf_clk new_AGEMA_reg_buffer_10497 ( .C (clk), .D (new_AGEMA_signal_31452), .Q (new_AGEMA_signal_31453) ) ;
    buf_clk new_AGEMA_reg_buffer_10500 ( .C (clk), .D (new_AGEMA_signal_31455), .Q (new_AGEMA_signal_31456) ) ;
    buf_clk new_AGEMA_reg_buffer_10503 ( .C (clk), .D (new_AGEMA_signal_31458), .Q (new_AGEMA_signal_31459) ) ;
    buf_clk new_AGEMA_reg_buffer_10506 ( .C (clk), .D (new_AGEMA_signal_31461), .Q (new_AGEMA_signal_31462) ) ;
    buf_clk new_AGEMA_reg_buffer_10509 ( .C (clk), .D (new_AGEMA_signal_31464), .Q (new_AGEMA_signal_31465) ) ;
    buf_clk new_AGEMA_reg_buffer_10512 ( .C (clk), .D (new_AGEMA_signal_31467), .Q (new_AGEMA_signal_31468) ) ;
    buf_clk new_AGEMA_reg_buffer_10515 ( .C (clk), .D (new_AGEMA_signal_31470), .Q (new_AGEMA_signal_31471) ) ;
    buf_clk new_AGEMA_reg_buffer_10518 ( .C (clk), .D (new_AGEMA_signal_31473), .Q (new_AGEMA_signal_31474) ) ;
    buf_clk new_AGEMA_reg_buffer_10521 ( .C (clk), .D (new_AGEMA_signal_31476), .Q (new_AGEMA_signal_31477) ) ;
    buf_clk new_AGEMA_reg_buffer_10524 ( .C (clk), .D (new_AGEMA_signal_31479), .Q (new_AGEMA_signal_31480) ) ;
    buf_clk new_AGEMA_reg_buffer_10527 ( .C (clk), .D (new_AGEMA_signal_31482), .Q (new_AGEMA_signal_31483) ) ;
    buf_clk new_AGEMA_reg_buffer_10530 ( .C (clk), .D (new_AGEMA_signal_31485), .Q (new_AGEMA_signal_31486) ) ;
    buf_clk new_AGEMA_reg_buffer_10533 ( .C (clk), .D (new_AGEMA_signal_31488), .Q (new_AGEMA_signal_31489) ) ;
    buf_clk new_AGEMA_reg_buffer_10536 ( .C (clk), .D (new_AGEMA_signal_31491), .Q (new_AGEMA_signal_31492) ) ;
    buf_clk new_AGEMA_reg_buffer_10539 ( .C (clk), .D (new_AGEMA_signal_31494), .Q (new_AGEMA_signal_31495) ) ;
    buf_clk new_AGEMA_reg_buffer_10542 ( .C (clk), .D (new_AGEMA_signal_31497), .Q (new_AGEMA_signal_31498) ) ;
    buf_clk new_AGEMA_reg_buffer_10545 ( .C (clk), .D (new_AGEMA_signal_31500), .Q (new_AGEMA_signal_31501) ) ;
    buf_clk new_AGEMA_reg_buffer_10548 ( .C (clk), .D (new_AGEMA_signal_31503), .Q (new_AGEMA_signal_31504) ) ;
    buf_clk new_AGEMA_reg_buffer_10551 ( .C (clk), .D (new_AGEMA_signal_31506), .Q (new_AGEMA_signal_31507) ) ;
    buf_clk new_AGEMA_reg_buffer_10554 ( .C (clk), .D (new_AGEMA_signal_31509), .Q (new_AGEMA_signal_31510) ) ;
    buf_clk new_AGEMA_reg_buffer_10557 ( .C (clk), .D (new_AGEMA_signal_31512), .Q (new_AGEMA_signal_31513) ) ;
    buf_clk new_AGEMA_reg_buffer_10560 ( .C (clk), .D (new_AGEMA_signal_31515), .Q (new_AGEMA_signal_31516) ) ;
    buf_clk new_AGEMA_reg_buffer_10563 ( .C (clk), .D (new_AGEMA_signal_31518), .Q (new_AGEMA_signal_31519) ) ;
    buf_clk new_AGEMA_reg_buffer_10566 ( .C (clk), .D (new_AGEMA_signal_31521), .Q (new_AGEMA_signal_31522) ) ;
    buf_clk new_AGEMA_reg_buffer_10569 ( .C (clk), .D (new_AGEMA_signal_31524), .Q (new_AGEMA_signal_31525) ) ;
    buf_clk new_AGEMA_reg_buffer_10572 ( .C (clk), .D (new_AGEMA_signal_31527), .Q (new_AGEMA_signal_31528) ) ;
    buf_clk new_AGEMA_reg_buffer_10575 ( .C (clk), .D (new_AGEMA_signal_31530), .Q (new_AGEMA_signal_31531) ) ;
    buf_clk new_AGEMA_reg_buffer_10578 ( .C (clk), .D (new_AGEMA_signal_31533), .Q (new_AGEMA_signal_31534) ) ;
    buf_clk new_AGEMA_reg_buffer_10581 ( .C (clk), .D (new_AGEMA_signal_31536), .Q (new_AGEMA_signal_31537) ) ;
    buf_clk new_AGEMA_reg_buffer_10584 ( .C (clk), .D (new_AGEMA_signal_31539), .Q (new_AGEMA_signal_31540) ) ;
    buf_clk new_AGEMA_reg_buffer_10587 ( .C (clk), .D (new_AGEMA_signal_31542), .Q (new_AGEMA_signal_31543) ) ;
    buf_clk new_AGEMA_reg_buffer_10590 ( .C (clk), .D (new_AGEMA_signal_31545), .Q (new_AGEMA_signal_31546) ) ;
    buf_clk new_AGEMA_reg_buffer_10593 ( .C (clk), .D (new_AGEMA_signal_31548), .Q (new_AGEMA_signal_31549) ) ;
    buf_clk new_AGEMA_reg_buffer_10596 ( .C (clk), .D (new_AGEMA_signal_31551), .Q (new_AGEMA_signal_31552) ) ;
    buf_clk new_AGEMA_reg_buffer_10599 ( .C (clk), .D (new_AGEMA_signal_31554), .Q (new_AGEMA_signal_31555) ) ;
    buf_clk new_AGEMA_reg_buffer_10602 ( .C (clk), .D (new_AGEMA_signal_31557), .Q (new_AGEMA_signal_31558) ) ;
    buf_clk new_AGEMA_reg_buffer_10605 ( .C (clk), .D (new_AGEMA_signal_31560), .Q (new_AGEMA_signal_31561) ) ;
    buf_clk new_AGEMA_reg_buffer_10608 ( .C (clk), .D (new_AGEMA_signal_31563), .Q (new_AGEMA_signal_31564) ) ;
    buf_clk new_AGEMA_reg_buffer_10611 ( .C (clk), .D (new_AGEMA_signal_31566), .Q (new_AGEMA_signal_31567) ) ;
    buf_clk new_AGEMA_reg_buffer_10614 ( .C (clk), .D (new_AGEMA_signal_31569), .Q (new_AGEMA_signal_31570) ) ;
    buf_clk new_AGEMA_reg_buffer_10617 ( .C (clk), .D (new_AGEMA_signal_31572), .Q (new_AGEMA_signal_31573) ) ;
    buf_clk new_AGEMA_reg_buffer_10620 ( .C (clk), .D (new_AGEMA_signal_31575), .Q (new_AGEMA_signal_31576) ) ;
    buf_clk new_AGEMA_reg_buffer_10623 ( .C (clk), .D (new_AGEMA_signal_31578), .Q (new_AGEMA_signal_31579) ) ;
    buf_clk new_AGEMA_reg_buffer_10626 ( .C (clk), .D (new_AGEMA_signal_31581), .Q (new_AGEMA_signal_31582) ) ;
    buf_clk new_AGEMA_reg_buffer_10629 ( .C (clk), .D (new_AGEMA_signal_31584), .Q (new_AGEMA_signal_31585) ) ;
    buf_clk new_AGEMA_reg_buffer_10632 ( .C (clk), .D (new_AGEMA_signal_31587), .Q (new_AGEMA_signal_31588) ) ;
    buf_clk new_AGEMA_reg_buffer_10635 ( .C (clk), .D (new_AGEMA_signal_31590), .Q (new_AGEMA_signal_31591) ) ;
    buf_clk new_AGEMA_reg_buffer_10638 ( .C (clk), .D (new_AGEMA_signal_31593), .Q (new_AGEMA_signal_31594) ) ;
    buf_clk new_AGEMA_reg_buffer_10641 ( .C (clk), .D (new_AGEMA_signal_31596), .Q (new_AGEMA_signal_31597) ) ;
    buf_clk new_AGEMA_reg_buffer_10644 ( .C (clk), .D (new_AGEMA_signal_31599), .Q (new_AGEMA_signal_31600) ) ;
    buf_clk new_AGEMA_reg_buffer_10647 ( .C (clk), .D (new_AGEMA_signal_31602), .Q (new_AGEMA_signal_31603) ) ;
    buf_clk new_AGEMA_reg_buffer_10650 ( .C (clk), .D (new_AGEMA_signal_31605), .Q (new_AGEMA_signal_31606) ) ;
    buf_clk new_AGEMA_reg_buffer_10653 ( .C (clk), .D (new_AGEMA_signal_31608), .Q (new_AGEMA_signal_31609) ) ;
    buf_clk new_AGEMA_reg_buffer_10656 ( .C (clk), .D (new_AGEMA_signal_31611), .Q (new_AGEMA_signal_31612) ) ;
    buf_clk new_AGEMA_reg_buffer_10659 ( .C (clk), .D (new_AGEMA_signal_31614), .Q (new_AGEMA_signal_31615) ) ;
    buf_clk new_AGEMA_reg_buffer_10662 ( .C (clk), .D (new_AGEMA_signal_31617), .Q (new_AGEMA_signal_31618) ) ;
    buf_clk new_AGEMA_reg_buffer_10665 ( .C (clk), .D (new_AGEMA_signal_31620), .Q (new_AGEMA_signal_31621) ) ;
    buf_clk new_AGEMA_reg_buffer_10668 ( .C (clk), .D (new_AGEMA_signal_31623), .Q (new_AGEMA_signal_31624) ) ;
    buf_clk new_AGEMA_reg_buffer_10671 ( .C (clk), .D (new_AGEMA_signal_31626), .Q (new_AGEMA_signal_31627) ) ;
    buf_clk new_AGEMA_reg_buffer_10674 ( .C (clk), .D (new_AGEMA_signal_31629), .Q (new_AGEMA_signal_31630) ) ;
    buf_clk new_AGEMA_reg_buffer_10677 ( .C (clk), .D (new_AGEMA_signal_31632), .Q (new_AGEMA_signal_31633) ) ;
    buf_clk new_AGEMA_reg_buffer_10680 ( .C (clk), .D (new_AGEMA_signal_31635), .Q (new_AGEMA_signal_31636) ) ;
    buf_clk new_AGEMA_reg_buffer_10683 ( .C (clk), .D (new_AGEMA_signal_31638), .Q (new_AGEMA_signal_31639) ) ;
    buf_clk new_AGEMA_reg_buffer_10686 ( .C (clk), .D (new_AGEMA_signal_31641), .Q (new_AGEMA_signal_31642) ) ;
    buf_clk new_AGEMA_reg_buffer_10689 ( .C (clk), .D (new_AGEMA_signal_31644), .Q (new_AGEMA_signal_31645) ) ;
    buf_clk new_AGEMA_reg_buffer_10692 ( .C (clk), .D (new_AGEMA_signal_31647), .Q (new_AGEMA_signal_31648) ) ;
    buf_clk new_AGEMA_reg_buffer_10695 ( .C (clk), .D (new_AGEMA_signal_31650), .Q (new_AGEMA_signal_31651) ) ;
    buf_clk new_AGEMA_reg_buffer_10698 ( .C (clk), .D (new_AGEMA_signal_31653), .Q (new_AGEMA_signal_31654) ) ;
    buf_clk new_AGEMA_reg_buffer_10701 ( .C (clk), .D (new_AGEMA_signal_31656), .Q (new_AGEMA_signal_31657) ) ;
    buf_clk new_AGEMA_reg_buffer_10704 ( .C (clk), .D (new_AGEMA_signal_31659), .Q (new_AGEMA_signal_31660) ) ;
    buf_clk new_AGEMA_reg_buffer_10707 ( .C (clk), .D (new_AGEMA_signal_31662), .Q (new_AGEMA_signal_31663) ) ;
    buf_clk new_AGEMA_reg_buffer_10711 ( .C (clk), .D (new_AGEMA_signal_31666), .Q (new_AGEMA_signal_31667) ) ;
    buf_clk new_AGEMA_reg_buffer_10715 ( .C (clk), .D (new_AGEMA_signal_31670), .Q (new_AGEMA_signal_31671) ) ;
    buf_clk new_AGEMA_reg_buffer_10719 ( .C (clk), .D (new_AGEMA_signal_31674), .Q (new_AGEMA_signal_31675) ) ;
    buf_clk new_AGEMA_reg_buffer_10723 ( .C (clk), .D (new_AGEMA_signal_31678), .Q (new_AGEMA_signal_31679) ) ;
    buf_clk new_AGEMA_reg_buffer_10727 ( .C (clk), .D (new_AGEMA_signal_31682), .Q (new_AGEMA_signal_31683) ) ;
    buf_clk new_AGEMA_reg_buffer_10731 ( .C (clk), .D (new_AGEMA_signal_31686), .Q (new_AGEMA_signal_31687) ) ;
    buf_clk new_AGEMA_reg_buffer_10735 ( .C (clk), .D (new_AGEMA_signal_31690), .Q (new_AGEMA_signal_31691) ) ;
    buf_clk new_AGEMA_reg_buffer_10739 ( .C (clk), .D (new_AGEMA_signal_31694), .Q (new_AGEMA_signal_31695) ) ;
    buf_clk new_AGEMA_reg_buffer_10743 ( .C (clk), .D (new_AGEMA_signal_31698), .Q (new_AGEMA_signal_31699) ) ;
    buf_clk new_AGEMA_reg_buffer_10747 ( .C (clk), .D (new_AGEMA_signal_31702), .Q (new_AGEMA_signal_31703) ) ;
    buf_clk new_AGEMA_reg_buffer_10751 ( .C (clk), .D (new_AGEMA_signal_31706), .Q (new_AGEMA_signal_31707) ) ;
    buf_clk new_AGEMA_reg_buffer_10755 ( .C (clk), .D (new_AGEMA_signal_31710), .Q (new_AGEMA_signal_31711) ) ;
    buf_clk new_AGEMA_reg_buffer_10759 ( .C (clk), .D (new_AGEMA_signal_31714), .Q (new_AGEMA_signal_31715) ) ;
    buf_clk new_AGEMA_reg_buffer_10763 ( .C (clk), .D (new_AGEMA_signal_31718), .Q (new_AGEMA_signal_31719) ) ;
    buf_clk new_AGEMA_reg_buffer_10767 ( .C (clk), .D (new_AGEMA_signal_31722), .Q (new_AGEMA_signal_31723) ) ;
    buf_clk new_AGEMA_reg_buffer_10771 ( .C (clk), .D (new_AGEMA_signal_31726), .Q (new_AGEMA_signal_31727) ) ;
    buf_clk new_AGEMA_reg_buffer_10775 ( .C (clk), .D (new_AGEMA_signal_31730), .Q (new_AGEMA_signal_31731) ) ;
    buf_clk new_AGEMA_reg_buffer_10779 ( .C (clk), .D (new_AGEMA_signal_31734), .Q (new_AGEMA_signal_31735) ) ;
    buf_clk new_AGEMA_reg_buffer_10783 ( .C (clk), .D (new_AGEMA_signal_31738), .Q (new_AGEMA_signal_31739) ) ;
    buf_clk new_AGEMA_reg_buffer_10787 ( .C (clk), .D (new_AGEMA_signal_31742), .Q (new_AGEMA_signal_31743) ) ;
    buf_clk new_AGEMA_reg_buffer_10791 ( .C (clk), .D (new_AGEMA_signal_31746), .Q (new_AGEMA_signal_31747) ) ;
    buf_clk new_AGEMA_reg_buffer_10795 ( .C (clk), .D (new_AGEMA_signal_31750), .Q (new_AGEMA_signal_31751) ) ;
    buf_clk new_AGEMA_reg_buffer_10799 ( .C (clk), .D (new_AGEMA_signal_31754), .Q (new_AGEMA_signal_31755) ) ;
    buf_clk new_AGEMA_reg_buffer_10803 ( .C (clk), .D (new_AGEMA_signal_31758), .Q (new_AGEMA_signal_31759) ) ;
    buf_clk new_AGEMA_reg_buffer_10807 ( .C (clk), .D (new_AGEMA_signal_31762), .Q (new_AGEMA_signal_31763) ) ;
    buf_clk new_AGEMA_reg_buffer_10811 ( .C (clk), .D (new_AGEMA_signal_31766), .Q (new_AGEMA_signal_31767) ) ;
    buf_clk new_AGEMA_reg_buffer_10815 ( .C (clk), .D (new_AGEMA_signal_31770), .Q (new_AGEMA_signal_31771) ) ;
    buf_clk new_AGEMA_reg_buffer_10819 ( .C (clk), .D (new_AGEMA_signal_31774), .Q (new_AGEMA_signal_31775) ) ;
    buf_clk new_AGEMA_reg_buffer_10823 ( .C (clk), .D (new_AGEMA_signal_31778), .Q (new_AGEMA_signal_31779) ) ;
    buf_clk new_AGEMA_reg_buffer_10827 ( .C (clk), .D (new_AGEMA_signal_31782), .Q (new_AGEMA_signal_31783) ) ;
    buf_clk new_AGEMA_reg_buffer_10831 ( .C (clk), .D (new_AGEMA_signal_31786), .Q (new_AGEMA_signal_31787) ) ;
    buf_clk new_AGEMA_reg_buffer_10835 ( .C (clk), .D (new_AGEMA_signal_31790), .Q (new_AGEMA_signal_31791) ) ;
    buf_clk new_AGEMA_reg_buffer_10839 ( .C (clk), .D (new_AGEMA_signal_31794), .Q (new_AGEMA_signal_31795) ) ;
    buf_clk new_AGEMA_reg_buffer_10843 ( .C (clk), .D (new_AGEMA_signal_31798), .Q (new_AGEMA_signal_31799) ) ;
    buf_clk new_AGEMA_reg_buffer_10847 ( .C (clk), .D (new_AGEMA_signal_31802), .Q (new_AGEMA_signal_31803) ) ;
    buf_clk new_AGEMA_reg_buffer_10851 ( .C (clk), .D (new_AGEMA_signal_31806), .Q (new_AGEMA_signal_31807) ) ;
    buf_clk new_AGEMA_reg_buffer_10855 ( .C (clk), .D (new_AGEMA_signal_31810), .Q (new_AGEMA_signal_31811) ) ;
    buf_clk new_AGEMA_reg_buffer_10859 ( .C (clk), .D (new_AGEMA_signal_31814), .Q (new_AGEMA_signal_31815) ) ;
    buf_clk new_AGEMA_reg_buffer_10863 ( .C (clk), .D (new_AGEMA_signal_31818), .Q (new_AGEMA_signal_31819) ) ;
    buf_clk new_AGEMA_reg_buffer_10867 ( .C (clk), .D (new_AGEMA_signal_31822), .Q (new_AGEMA_signal_31823) ) ;
    buf_clk new_AGEMA_reg_buffer_10871 ( .C (clk), .D (new_AGEMA_signal_31826), .Q (new_AGEMA_signal_31827) ) ;
    buf_clk new_AGEMA_reg_buffer_10875 ( .C (clk), .D (new_AGEMA_signal_31830), .Q (new_AGEMA_signal_31831) ) ;
    buf_clk new_AGEMA_reg_buffer_10879 ( .C (clk), .D (new_AGEMA_signal_31834), .Q (new_AGEMA_signal_31835) ) ;
    buf_clk new_AGEMA_reg_buffer_10883 ( .C (clk), .D (new_AGEMA_signal_31838), .Q (new_AGEMA_signal_31839) ) ;
    buf_clk new_AGEMA_reg_buffer_10887 ( .C (clk), .D (new_AGEMA_signal_31842), .Q (new_AGEMA_signal_31843) ) ;
    buf_clk new_AGEMA_reg_buffer_10891 ( .C (clk), .D (new_AGEMA_signal_31846), .Q (new_AGEMA_signal_31847) ) ;
    buf_clk new_AGEMA_reg_buffer_10895 ( .C (clk), .D (new_AGEMA_signal_31850), .Q (new_AGEMA_signal_31851) ) ;
    buf_clk new_AGEMA_reg_buffer_10899 ( .C (clk), .D (new_AGEMA_signal_31854), .Q (new_AGEMA_signal_31855) ) ;
    buf_clk new_AGEMA_reg_buffer_10903 ( .C (clk), .D (new_AGEMA_signal_31858), .Q (new_AGEMA_signal_31859) ) ;
    buf_clk new_AGEMA_reg_buffer_10907 ( .C (clk), .D (new_AGEMA_signal_31862), .Q (new_AGEMA_signal_31863) ) ;
    buf_clk new_AGEMA_reg_buffer_10911 ( .C (clk), .D (new_AGEMA_signal_31866), .Q (new_AGEMA_signal_31867) ) ;
    buf_clk new_AGEMA_reg_buffer_10915 ( .C (clk), .D (new_AGEMA_signal_31870), .Q (new_AGEMA_signal_31871) ) ;
    buf_clk new_AGEMA_reg_buffer_10919 ( .C (clk), .D (new_AGEMA_signal_31874), .Q (new_AGEMA_signal_31875) ) ;
    buf_clk new_AGEMA_reg_buffer_10923 ( .C (clk), .D (new_AGEMA_signal_31878), .Q (new_AGEMA_signal_31879) ) ;
    buf_clk new_AGEMA_reg_buffer_10927 ( .C (clk), .D (new_AGEMA_signal_31882), .Q (new_AGEMA_signal_31883) ) ;
    buf_clk new_AGEMA_reg_buffer_10931 ( .C (clk), .D (new_AGEMA_signal_31886), .Q (new_AGEMA_signal_31887) ) ;
    buf_clk new_AGEMA_reg_buffer_10935 ( .C (clk), .D (new_AGEMA_signal_31890), .Q (new_AGEMA_signal_31891) ) ;
    buf_clk new_AGEMA_reg_buffer_10939 ( .C (clk), .D (new_AGEMA_signal_31894), .Q (new_AGEMA_signal_31895) ) ;
    buf_clk new_AGEMA_reg_buffer_10943 ( .C (clk), .D (new_AGEMA_signal_31898), .Q (new_AGEMA_signal_31899) ) ;
    buf_clk new_AGEMA_reg_buffer_10947 ( .C (clk), .D (new_AGEMA_signal_31902), .Q (new_AGEMA_signal_31903) ) ;
    buf_clk new_AGEMA_reg_buffer_10951 ( .C (clk), .D (new_AGEMA_signal_31906), .Q (new_AGEMA_signal_31907) ) ;
    buf_clk new_AGEMA_reg_buffer_10955 ( .C (clk), .D (new_AGEMA_signal_31910), .Q (new_AGEMA_signal_31911) ) ;
    buf_clk new_AGEMA_reg_buffer_10959 ( .C (clk), .D (new_AGEMA_signal_31914), .Q (new_AGEMA_signal_31915) ) ;
    buf_clk new_AGEMA_reg_buffer_10963 ( .C (clk), .D (new_AGEMA_signal_31918), .Q (new_AGEMA_signal_31919) ) ;
    buf_clk new_AGEMA_reg_buffer_10967 ( .C (clk), .D (new_AGEMA_signal_31922), .Q (new_AGEMA_signal_31923) ) ;
    buf_clk new_AGEMA_reg_buffer_10971 ( .C (clk), .D (new_AGEMA_signal_31926), .Q (new_AGEMA_signal_31927) ) ;
    buf_clk new_AGEMA_reg_buffer_10975 ( .C (clk), .D (new_AGEMA_signal_31930), .Q (new_AGEMA_signal_31931) ) ;
    buf_clk new_AGEMA_reg_buffer_10979 ( .C (clk), .D (new_AGEMA_signal_31934), .Q (new_AGEMA_signal_31935) ) ;
    buf_clk new_AGEMA_reg_buffer_10983 ( .C (clk), .D (new_AGEMA_signal_31938), .Q (new_AGEMA_signal_31939) ) ;
    buf_clk new_AGEMA_reg_buffer_10987 ( .C (clk), .D (new_AGEMA_signal_31942), .Q (new_AGEMA_signal_31943) ) ;
    buf_clk new_AGEMA_reg_buffer_10991 ( .C (clk), .D (new_AGEMA_signal_31946), .Q (new_AGEMA_signal_31947) ) ;
    buf_clk new_AGEMA_reg_buffer_10995 ( .C (clk), .D (new_AGEMA_signal_31950), .Q (new_AGEMA_signal_31951) ) ;
    buf_clk new_AGEMA_reg_buffer_10999 ( .C (clk), .D (new_AGEMA_signal_31954), .Q (new_AGEMA_signal_31955) ) ;
    buf_clk new_AGEMA_reg_buffer_11003 ( .C (clk), .D (new_AGEMA_signal_31958), .Q (new_AGEMA_signal_31959) ) ;
    buf_clk new_AGEMA_reg_buffer_11007 ( .C (clk), .D (new_AGEMA_signal_31962), .Q (new_AGEMA_signal_31963) ) ;
    buf_clk new_AGEMA_reg_buffer_11011 ( .C (clk), .D (new_AGEMA_signal_31966), .Q (new_AGEMA_signal_31967) ) ;
    buf_clk new_AGEMA_reg_buffer_11015 ( .C (clk), .D (new_AGEMA_signal_31970), .Q (new_AGEMA_signal_31971) ) ;
    buf_clk new_AGEMA_reg_buffer_11019 ( .C (clk), .D (new_AGEMA_signal_31974), .Q (new_AGEMA_signal_31975) ) ;
    buf_clk new_AGEMA_reg_buffer_11023 ( .C (clk), .D (new_AGEMA_signal_31978), .Q (new_AGEMA_signal_31979) ) ;
    buf_clk new_AGEMA_reg_buffer_11027 ( .C (clk), .D (new_AGEMA_signal_31982), .Q (new_AGEMA_signal_31983) ) ;
    buf_clk new_AGEMA_reg_buffer_11031 ( .C (clk), .D (new_AGEMA_signal_31986), .Q (new_AGEMA_signal_31987) ) ;
    buf_clk new_AGEMA_reg_buffer_11035 ( .C (clk), .D (new_AGEMA_signal_31990), .Q (new_AGEMA_signal_31991) ) ;
    buf_clk new_AGEMA_reg_buffer_11039 ( .C (clk), .D (new_AGEMA_signal_31994), .Q (new_AGEMA_signal_31995) ) ;
    buf_clk new_AGEMA_reg_buffer_11043 ( .C (clk), .D (new_AGEMA_signal_31998), .Q (new_AGEMA_signal_31999) ) ;
    buf_clk new_AGEMA_reg_buffer_11047 ( .C (clk), .D (new_AGEMA_signal_32002), .Q (new_AGEMA_signal_32003) ) ;
    buf_clk new_AGEMA_reg_buffer_11051 ( .C (clk), .D (new_AGEMA_signal_32006), .Q (new_AGEMA_signal_32007) ) ;
    buf_clk new_AGEMA_reg_buffer_11055 ( .C (clk), .D (new_AGEMA_signal_32010), .Q (new_AGEMA_signal_32011) ) ;
    buf_clk new_AGEMA_reg_buffer_11059 ( .C (clk), .D (new_AGEMA_signal_32014), .Q (new_AGEMA_signal_32015) ) ;
    buf_clk new_AGEMA_reg_buffer_11063 ( .C (clk), .D (new_AGEMA_signal_32018), .Q (new_AGEMA_signal_32019) ) ;
    buf_clk new_AGEMA_reg_buffer_11067 ( .C (clk), .D (new_AGEMA_signal_32022), .Q (new_AGEMA_signal_32023) ) ;
    buf_clk new_AGEMA_reg_buffer_11071 ( .C (clk), .D (new_AGEMA_signal_32026), .Q (new_AGEMA_signal_32027) ) ;
    buf_clk new_AGEMA_reg_buffer_11075 ( .C (clk), .D (new_AGEMA_signal_32030), .Q (new_AGEMA_signal_32031) ) ;
    buf_clk new_AGEMA_reg_buffer_11079 ( .C (clk), .D (new_AGEMA_signal_32034), .Q (new_AGEMA_signal_32035) ) ;
    buf_clk new_AGEMA_reg_buffer_11083 ( .C (clk), .D (new_AGEMA_signal_32038), .Q (new_AGEMA_signal_32039) ) ;
    buf_clk new_AGEMA_reg_buffer_11087 ( .C (clk), .D (new_AGEMA_signal_32042), .Q (new_AGEMA_signal_32043) ) ;
    buf_clk new_AGEMA_reg_buffer_11091 ( .C (clk), .D (new_AGEMA_signal_32046), .Q (new_AGEMA_signal_32047) ) ;
    buf_clk new_AGEMA_reg_buffer_11095 ( .C (clk), .D (new_AGEMA_signal_32050), .Q (new_AGEMA_signal_32051) ) ;
    buf_clk new_AGEMA_reg_buffer_11099 ( .C (clk), .D (new_AGEMA_signal_32054), .Q (new_AGEMA_signal_32055) ) ;
    buf_clk new_AGEMA_reg_buffer_11103 ( .C (clk), .D (new_AGEMA_signal_32058), .Q (new_AGEMA_signal_32059) ) ;
    buf_clk new_AGEMA_reg_buffer_11107 ( .C (clk), .D (new_AGEMA_signal_32062), .Q (new_AGEMA_signal_32063) ) ;
    buf_clk new_AGEMA_reg_buffer_11111 ( .C (clk), .D (new_AGEMA_signal_32066), .Q (new_AGEMA_signal_32067) ) ;
    buf_clk new_AGEMA_reg_buffer_11115 ( .C (clk), .D (new_AGEMA_signal_32070), .Q (new_AGEMA_signal_32071) ) ;
    buf_clk new_AGEMA_reg_buffer_11119 ( .C (clk), .D (new_AGEMA_signal_32074), .Q (new_AGEMA_signal_32075) ) ;
    buf_clk new_AGEMA_reg_buffer_11123 ( .C (clk), .D (new_AGEMA_signal_32078), .Q (new_AGEMA_signal_32079) ) ;
    buf_clk new_AGEMA_reg_buffer_11127 ( .C (clk), .D (new_AGEMA_signal_32082), .Q (new_AGEMA_signal_32083) ) ;
    buf_clk new_AGEMA_reg_buffer_11131 ( .C (clk), .D (new_AGEMA_signal_32086), .Q (new_AGEMA_signal_32087) ) ;
    buf_clk new_AGEMA_reg_buffer_11135 ( .C (clk), .D (new_AGEMA_signal_32090), .Q (new_AGEMA_signal_32091) ) ;
    buf_clk new_AGEMA_reg_buffer_11139 ( .C (clk), .D (new_AGEMA_signal_32094), .Q (new_AGEMA_signal_32095) ) ;
    buf_clk new_AGEMA_reg_buffer_11143 ( .C (clk), .D (new_AGEMA_signal_32098), .Q (new_AGEMA_signal_32099) ) ;
    buf_clk new_AGEMA_reg_buffer_11147 ( .C (clk), .D (new_AGEMA_signal_32102), .Q (new_AGEMA_signal_32103) ) ;
    buf_clk new_AGEMA_reg_buffer_11151 ( .C (clk), .D (new_AGEMA_signal_32106), .Q (new_AGEMA_signal_32107) ) ;
    buf_clk new_AGEMA_reg_buffer_11155 ( .C (clk), .D (new_AGEMA_signal_32110), .Q (new_AGEMA_signal_32111) ) ;
    buf_clk new_AGEMA_reg_buffer_11159 ( .C (clk), .D (new_AGEMA_signal_32114), .Q (new_AGEMA_signal_32115) ) ;
    buf_clk new_AGEMA_reg_buffer_11163 ( .C (clk), .D (new_AGEMA_signal_32118), .Q (new_AGEMA_signal_32119) ) ;
    buf_clk new_AGEMA_reg_buffer_11167 ( .C (clk), .D (new_AGEMA_signal_32122), .Q (new_AGEMA_signal_32123) ) ;
    buf_clk new_AGEMA_reg_buffer_11171 ( .C (clk), .D (new_AGEMA_signal_32126), .Q (new_AGEMA_signal_32127) ) ;
    buf_clk new_AGEMA_reg_buffer_11175 ( .C (clk), .D (new_AGEMA_signal_32130), .Q (new_AGEMA_signal_32131) ) ;
    buf_clk new_AGEMA_reg_buffer_11179 ( .C (clk), .D (new_AGEMA_signal_32134), .Q (new_AGEMA_signal_32135) ) ;
    buf_clk new_AGEMA_reg_buffer_11183 ( .C (clk), .D (new_AGEMA_signal_32138), .Q (new_AGEMA_signal_32139) ) ;
    buf_clk new_AGEMA_reg_buffer_11187 ( .C (clk), .D (new_AGEMA_signal_32142), .Q (new_AGEMA_signal_32143) ) ;
    buf_clk new_AGEMA_reg_buffer_11191 ( .C (clk), .D (new_AGEMA_signal_32146), .Q (new_AGEMA_signal_32147) ) ;
    buf_clk new_AGEMA_reg_buffer_11195 ( .C (clk), .D (new_AGEMA_signal_32150), .Q (new_AGEMA_signal_32151) ) ;
    buf_clk new_AGEMA_reg_buffer_11199 ( .C (clk), .D (new_AGEMA_signal_32154), .Q (new_AGEMA_signal_32155) ) ;
    buf_clk new_AGEMA_reg_buffer_11203 ( .C (clk), .D (new_AGEMA_signal_32158), .Q (new_AGEMA_signal_32159) ) ;
    buf_clk new_AGEMA_reg_buffer_11207 ( .C (clk), .D (new_AGEMA_signal_32162), .Q (new_AGEMA_signal_32163) ) ;
    buf_clk new_AGEMA_reg_buffer_11211 ( .C (clk), .D (new_AGEMA_signal_32166), .Q (new_AGEMA_signal_32167) ) ;
    buf_clk new_AGEMA_reg_buffer_11215 ( .C (clk), .D (new_AGEMA_signal_32170), .Q (new_AGEMA_signal_32171) ) ;
    buf_clk new_AGEMA_reg_buffer_11219 ( .C (clk), .D (new_AGEMA_signal_32174), .Q (new_AGEMA_signal_32175) ) ;
    buf_clk new_AGEMA_reg_buffer_11223 ( .C (clk), .D (new_AGEMA_signal_32178), .Q (new_AGEMA_signal_32179) ) ;
    buf_clk new_AGEMA_reg_buffer_11227 ( .C (clk), .D (new_AGEMA_signal_32182), .Q (new_AGEMA_signal_32183) ) ;
    buf_clk new_AGEMA_reg_buffer_11231 ( .C (clk), .D (new_AGEMA_signal_32186), .Q (new_AGEMA_signal_32187) ) ;
    buf_clk new_AGEMA_reg_buffer_11235 ( .C (clk), .D (new_AGEMA_signal_32190), .Q (new_AGEMA_signal_32191) ) ;
    buf_clk new_AGEMA_reg_buffer_11239 ( .C (clk), .D (new_AGEMA_signal_32194), .Q (new_AGEMA_signal_32195) ) ;
    buf_clk new_AGEMA_reg_buffer_11243 ( .C (clk), .D (new_AGEMA_signal_32198), .Q (new_AGEMA_signal_32199) ) ;
    buf_clk new_AGEMA_reg_buffer_11247 ( .C (clk), .D (new_AGEMA_signal_32202), .Q (new_AGEMA_signal_32203) ) ;
    buf_clk new_AGEMA_reg_buffer_11251 ( .C (clk), .D (new_AGEMA_signal_32206), .Q (new_AGEMA_signal_32207) ) ;
    buf_clk new_AGEMA_reg_buffer_11255 ( .C (clk), .D (new_AGEMA_signal_32210), .Q (new_AGEMA_signal_32211) ) ;
    buf_clk new_AGEMA_reg_buffer_11259 ( .C (clk), .D (new_AGEMA_signal_32214), .Q (new_AGEMA_signal_32215) ) ;
    buf_clk new_AGEMA_reg_buffer_11263 ( .C (clk), .D (new_AGEMA_signal_32218), .Q (new_AGEMA_signal_32219) ) ;
    buf_clk new_AGEMA_reg_buffer_11267 ( .C (clk), .D (new_AGEMA_signal_32222), .Q (new_AGEMA_signal_32223) ) ;
    buf_clk new_AGEMA_reg_buffer_11271 ( .C (clk), .D (new_AGEMA_signal_32226), .Q (new_AGEMA_signal_32227) ) ;
    buf_clk new_AGEMA_reg_buffer_11275 ( .C (clk), .D (new_AGEMA_signal_32230), .Q (new_AGEMA_signal_32231) ) ;
    buf_clk new_AGEMA_reg_buffer_11279 ( .C (clk), .D (new_AGEMA_signal_32234), .Q (new_AGEMA_signal_32235) ) ;
    buf_clk new_AGEMA_reg_buffer_11283 ( .C (clk), .D (new_AGEMA_signal_32238), .Q (new_AGEMA_signal_32239) ) ;
    buf_clk new_AGEMA_reg_buffer_11287 ( .C (clk), .D (new_AGEMA_signal_32242), .Q (new_AGEMA_signal_32243) ) ;
    buf_clk new_AGEMA_reg_buffer_11291 ( .C (clk), .D (new_AGEMA_signal_32246), .Q (new_AGEMA_signal_32247) ) ;
    buf_clk new_AGEMA_reg_buffer_11295 ( .C (clk), .D (new_AGEMA_signal_32250), .Q (new_AGEMA_signal_32251) ) ;
    buf_clk new_AGEMA_reg_buffer_11299 ( .C (clk), .D (new_AGEMA_signal_32254), .Q (new_AGEMA_signal_32255) ) ;
    buf_clk new_AGEMA_reg_buffer_11303 ( .C (clk), .D (new_AGEMA_signal_32258), .Q (new_AGEMA_signal_32259) ) ;
    buf_clk new_AGEMA_reg_buffer_11307 ( .C (clk), .D (new_AGEMA_signal_32262), .Q (new_AGEMA_signal_32263) ) ;
    buf_clk new_AGEMA_reg_buffer_11311 ( .C (clk), .D (new_AGEMA_signal_32266), .Q (new_AGEMA_signal_32267) ) ;
    buf_clk new_AGEMA_reg_buffer_11315 ( .C (clk), .D (new_AGEMA_signal_32270), .Q (new_AGEMA_signal_32271) ) ;
    buf_clk new_AGEMA_reg_buffer_11319 ( .C (clk), .D (new_AGEMA_signal_32274), .Q (new_AGEMA_signal_32275) ) ;
    buf_clk new_AGEMA_reg_buffer_11323 ( .C (clk), .D (new_AGEMA_signal_32278), .Q (new_AGEMA_signal_32279) ) ;
    buf_clk new_AGEMA_reg_buffer_11327 ( .C (clk), .D (new_AGEMA_signal_32282), .Q (new_AGEMA_signal_32283) ) ;
    buf_clk new_AGEMA_reg_buffer_11331 ( .C (clk), .D (new_AGEMA_signal_32286), .Q (new_AGEMA_signal_32287) ) ;
    buf_clk new_AGEMA_reg_buffer_11335 ( .C (clk), .D (new_AGEMA_signal_32290), .Q (new_AGEMA_signal_32291) ) ;
    buf_clk new_AGEMA_reg_buffer_11339 ( .C (clk), .D (new_AGEMA_signal_32294), .Q (new_AGEMA_signal_32295) ) ;
    buf_clk new_AGEMA_reg_buffer_11343 ( .C (clk), .D (new_AGEMA_signal_32298), .Q (new_AGEMA_signal_32299) ) ;
    buf_clk new_AGEMA_reg_buffer_11347 ( .C (clk), .D (new_AGEMA_signal_32302), .Q (new_AGEMA_signal_32303) ) ;
    buf_clk new_AGEMA_reg_buffer_11351 ( .C (clk), .D (new_AGEMA_signal_32306), .Q (new_AGEMA_signal_32307) ) ;
    buf_clk new_AGEMA_reg_buffer_11355 ( .C (clk), .D (new_AGEMA_signal_32310), .Q (new_AGEMA_signal_32311) ) ;
    buf_clk new_AGEMA_reg_buffer_11359 ( .C (clk), .D (new_AGEMA_signal_32314), .Q (new_AGEMA_signal_32315) ) ;
    buf_clk new_AGEMA_reg_buffer_11363 ( .C (clk), .D (new_AGEMA_signal_32318), .Q (new_AGEMA_signal_32319) ) ;
    buf_clk new_AGEMA_reg_buffer_11367 ( .C (clk), .D (new_AGEMA_signal_32322), .Q (new_AGEMA_signal_32323) ) ;
    buf_clk new_AGEMA_reg_buffer_11371 ( .C (clk), .D (new_AGEMA_signal_32326), .Q (new_AGEMA_signal_32327) ) ;
    buf_clk new_AGEMA_reg_buffer_11375 ( .C (clk), .D (new_AGEMA_signal_32330), .Q (new_AGEMA_signal_32331) ) ;
    buf_clk new_AGEMA_reg_buffer_11379 ( .C (clk), .D (new_AGEMA_signal_32334), .Q (new_AGEMA_signal_32335) ) ;
    buf_clk new_AGEMA_reg_buffer_11383 ( .C (clk), .D (new_AGEMA_signal_32338), .Q (new_AGEMA_signal_32339) ) ;
    buf_clk new_AGEMA_reg_buffer_11387 ( .C (clk), .D (new_AGEMA_signal_32342), .Q (new_AGEMA_signal_32343) ) ;
    buf_clk new_AGEMA_reg_buffer_11391 ( .C (clk), .D (new_AGEMA_signal_32346), .Q (new_AGEMA_signal_32347) ) ;
    buf_clk new_AGEMA_reg_buffer_11395 ( .C (clk), .D (new_AGEMA_signal_32350), .Q (new_AGEMA_signal_32351) ) ;
    buf_clk new_AGEMA_reg_buffer_11399 ( .C (clk), .D (new_AGEMA_signal_32354), .Q (new_AGEMA_signal_32355) ) ;
    buf_clk new_AGEMA_reg_buffer_11403 ( .C (clk), .D (new_AGEMA_signal_32358), .Q (new_AGEMA_signal_32359) ) ;
    buf_clk new_AGEMA_reg_buffer_11407 ( .C (clk), .D (new_AGEMA_signal_32362), .Q (new_AGEMA_signal_32363) ) ;
    buf_clk new_AGEMA_reg_buffer_11411 ( .C (clk), .D (new_AGEMA_signal_32366), .Q (new_AGEMA_signal_32367) ) ;
    buf_clk new_AGEMA_reg_buffer_11415 ( .C (clk), .D (new_AGEMA_signal_32370), .Q (new_AGEMA_signal_32371) ) ;
    buf_clk new_AGEMA_reg_buffer_11419 ( .C (clk), .D (new_AGEMA_signal_32374), .Q (new_AGEMA_signal_32375) ) ;
    buf_clk new_AGEMA_reg_buffer_11423 ( .C (clk), .D (new_AGEMA_signal_32378), .Q (new_AGEMA_signal_32379) ) ;
    buf_clk new_AGEMA_reg_buffer_11427 ( .C (clk), .D (new_AGEMA_signal_32382), .Q (new_AGEMA_signal_32383) ) ;
    buf_clk new_AGEMA_reg_buffer_11431 ( .C (clk), .D (new_AGEMA_signal_32386), .Q (new_AGEMA_signal_32387) ) ;
    buf_clk new_AGEMA_reg_buffer_11435 ( .C (clk), .D (new_AGEMA_signal_32390), .Q (new_AGEMA_signal_32391) ) ;
    buf_clk new_AGEMA_reg_buffer_11439 ( .C (clk), .D (new_AGEMA_signal_32394), .Q (new_AGEMA_signal_32395) ) ;
    buf_clk new_AGEMA_reg_buffer_11443 ( .C (clk), .D (new_AGEMA_signal_32398), .Q (new_AGEMA_signal_32399) ) ;
    buf_clk new_AGEMA_reg_buffer_11447 ( .C (clk), .D (new_AGEMA_signal_32402), .Q (new_AGEMA_signal_32403) ) ;
    buf_clk new_AGEMA_reg_buffer_11451 ( .C (clk), .D (new_AGEMA_signal_32406), .Q (new_AGEMA_signal_32407) ) ;
    buf_clk new_AGEMA_reg_buffer_11455 ( .C (clk), .D (new_AGEMA_signal_32410), .Q (new_AGEMA_signal_32411) ) ;
    buf_clk new_AGEMA_reg_buffer_11459 ( .C (clk), .D (new_AGEMA_signal_32414), .Q (new_AGEMA_signal_32415) ) ;
    buf_clk new_AGEMA_reg_buffer_11463 ( .C (clk), .D (new_AGEMA_signal_32418), .Q (new_AGEMA_signal_32419) ) ;
    buf_clk new_AGEMA_reg_buffer_11467 ( .C (clk), .D (new_AGEMA_signal_32422), .Q (new_AGEMA_signal_32423) ) ;
    buf_clk new_AGEMA_reg_buffer_11471 ( .C (clk), .D (new_AGEMA_signal_32426), .Q (new_AGEMA_signal_32427) ) ;
    buf_clk new_AGEMA_reg_buffer_11475 ( .C (clk), .D (new_AGEMA_signal_32430), .Q (new_AGEMA_signal_32431) ) ;
    buf_clk new_AGEMA_reg_buffer_11479 ( .C (clk), .D (new_AGEMA_signal_32434), .Q (new_AGEMA_signal_32435) ) ;
    buf_clk new_AGEMA_reg_buffer_11483 ( .C (clk), .D (new_AGEMA_signal_32438), .Q (new_AGEMA_signal_32439) ) ;
    buf_clk new_AGEMA_reg_buffer_11487 ( .C (clk), .D (new_AGEMA_signal_32442), .Q (new_AGEMA_signal_32443) ) ;
    buf_clk new_AGEMA_reg_buffer_11491 ( .C (clk), .D (new_AGEMA_signal_32446), .Q (new_AGEMA_signal_32447) ) ;
    buf_clk new_AGEMA_reg_buffer_11495 ( .C (clk), .D (new_AGEMA_signal_32450), .Q (new_AGEMA_signal_32451) ) ;
    buf_clk new_AGEMA_reg_buffer_11499 ( .C (clk), .D (new_AGEMA_signal_32454), .Q (new_AGEMA_signal_32455) ) ;
    buf_clk new_AGEMA_reg_buffer_11503 ( .C (clk), .D (new_AGEMA_signal_32458), .Q (new_AGEMA_signal_32459) ) ;
    buf_clk new_AGEMA_reg_buffer_11507 ( .C (clk), .D (new_AGEMA_signal_32462), .Q (new_AGEMA_signal_32463) ) ;
    buf_clk new_AGEMA_reg_buffer_11511 ( .C (clk), .D (new_AGEMA_signal_32466), .Q (new_AGEMA_signal_32467) ) ;
    buf_clk new_AGEMA_reg_buffer_11515 ( .C (clk), .D (new_AGEMA_signal_32470), .Q (new_AGEMA_signal_32471) ) ;
    buf_clk new_AGEMA_reg_buffer_11519 ( .C (clk), .D (new_AGEMA_signal_32474), .Q (new_AGEMA_signal_32475) ) ;
    buf_clk new_AGEMA_reg_buffer_11523 ( .C (clk), .D (new_AGEMA_signal_32478), .Q (new_AGEMA_signal_32479) ) ;
    buf_clk new_AGEMA_reg_buffer_11527 ( .C (clk), .D (new_AGEMA_signal_32482), .Q (new_AGEMA_signal_32483) ) ;
    buf_clk new_AGEMA_reg_buffer_11531 ( .C (clk), .D (new_AGEMA_signal_32486), .Q (new_AGEMA_signal_32487) ) ;
    buf_clk new_AGEMA_reg_buffer_11535 ( .C (clk), .D (new_AGEMA_signal_32490), .Q (new_AGEMA_signal_32491) ) ;
    buf_clk new_AGEMA_reg_buffer_11539 ( .C (clk), .D (new_AGEMA_signal_32494), .Q (new_AGEMA_signal_32495) ) ;
    buf_clk new_AGEMA_reg_buffer_11543 ( .C (clk), .D (new_AGEMA_signal_32498), .Q (new_AGEMA_signal_32499) ) ;
    buf_clk new_AGEMA_reg_buffer_11547 ( .C (clk), .D (new_AGEMA_signal_32502), .Q (new_AGEMA_signal_32503) ) ;
    buf_clk new_AGEMA_reg_buffer_11551 ( .C (clk), .D (new_AGEMA_signal_32506), .Q (new_AGEMA_signal_32507) ) ;
    buf_clk new_AGEMA_reg_buffer_11555 ( .C (clk), .D (new_AGEMA_signal_32510), .Q (new_AGEMA_signal_32511) ) ;
    buf_clk new_AGEMA_reg_buffer_11559 ( .C (clk), .D (new_AGEMA_signal_32514), .Q (new_AGEMA_signal_32515) ) ;
    buf_clk new_AGEMA_reg_buffer_11563 ( .C (clk), .D (new_AGEMA_signal_32518), .Q (new_AGEMA_signal_32519) ) ;
    buf_clk new_AGEMA_reg_buffer_11567 ( .C (clk), .D (new_AGEMA_signal_32522), .Q (new_AGEMA_signal_32523) ) ;
    buf_clk new_AGEMA_reg_buffer_11571 ( .C (clk), .D (new_AGEMA_signal_32526), .Q (new_AGEMA_signal_32527) ) ;
    buf_clk new_AGEMA_reg_buffer_11575 ( .C (clk), .D (new_AGEMA_signal_32530), .Q (new_AGEMA_signal_32531) ) ;
    buf_clk new_AGEMA_reg_buffer_11579 ( .C (clk), .D (new_AGEMA_signal_32534), .Q (new_AGEMA_signal_32535) ) ;
    buf_clk new_AGEMA_reg_buffer_11583 ( .C (clk), .D (new_AGEMA_signal_32538), .Q (new_AGEMA_signal_32539) ) ;
    buf_clk new_AGEMA_reg_buffer_11587 ( .C (clk), .D (new_AGEMA_signal_32542), .Q (new_AGEMA_signal_32543) ) ;
    buf_clk new_AGEMA_reg_buffer_11591 ( .C (clk), .D (new_AGEMA_signal_32546), .Q (new_AGEMA_signal_32547) ) ;
    buf_clk new_AGEMA_reg_buffer_11595 ( .C (clk), .D (new_AGEMA_signal_32550), .Q (new_AGEMA_signal_32551) ) ;
    buf_clk new_AGEMA_reg_buffer_11599 ( .C (clk), .D (new_AGEMA_signal_32554), .Q (new_AGEMA_signal_32555) ) ;
    buf_clk new_AGEMA_reg_buffer_11603 ( .C (clk), .D (new_AGEMA_signal_32558), .Q (new_AGEMA_signal_32559) ) ;
    buf_clk new_AGEMA_reg_buffer_11607 ( .C (clk), .D (new_AGEMA_signal_32562), .Q (new_AGEMA_signal_32563) ) ;
    buf_clk new_AGEMA_reg_buffer_11611 ( .C (clk), .D (new_AGEMA_signal_32566), .Q (new_AGEMA_signal_32567) ) ;
    buf_clk new_AGEMA_reg_buffer_11615 ( .C (clk), .D (new_AGEMA_signal_32570), .Q (new_AGEMA_signal_32571) ) ;
    buf_clk new_AGEMA_reg_buffer_11619 ( .C (clk), .D (new_AGEMA_signal_32574), .Q (new_AGEMA_signal_32575) ) ;
    buf_clk new_AGEMA_reg_buffer_11623 ( .C (clk), .D (new_AGEMA_signal_32578), .Q (new_AGEMA_signal_32579) ) ;
    buf_clk new_AGEMA_reg_buffer_11627 ( .C (clk), .D (new_AGEMA_signal_32582), .Q (new_AGEMA_signal_32583) ) ;
    buf_clk new_AGEMA_reg_buffer_11631 ( .C (clk), .D (new_AGEMA_signal_32586), .Q (new_AGEMA_signal_32587) ) ;
    buf_clk new_AGEMA_reg_buffer_11635 ( .C (clk), .D (new_AGEMA_signal_32590), .Q (new_AGEMA_signal_32591) ) ;
    buf_clk new_AGEMA_reg_buffer_11639 ( .C (clk), .D (new_AGEMA_signal_32594), .Q (new_AGEMA_signal_32595) ) ;
    buf_clk new_AGEMA_reg_buffer_11643 ( .C (clk), .D (new_AGEMA_signal_32598), .Q (new_AGEMA_signal_32599) ) ;
    buf_clk new_AGEMA_reg_buffer_11647 ( .C (clk), .D (new_AGEMA_signal_32602), .Q (new_AGEMA_signal_32603) ) ;
    buf_clk new_AGEMA_reg_buffer_11651 ( .C (clk), .D (new_AGEMA_signal_32606), .Q (new_AGEMA_signal_32607) ) ;
    buf_clk new_AGEMA_reg_buffer_11655 ( .C (clk), .D (new_AGEMA_signal_32610), .Q (new_AGEMA_signal_32611) ) ;
    buf_clk new_AGEMA_reg_buffer_11659 ( .C (clk), .D (new_AGEMA_signal_32614), .Q (new_AGEMA_signal_32615) ) ;
    buf_clk new_AGEMA_reg_buffer_11663 ( .C (clk), .D (new_AGEMA_signal_32618), .Q (new_AGEMA_signal_32619) ) ;
    buf_clk new_AGEMA_reg_buffer_11667 ( .C (clk), .D (new_AGEMA_signal_32622), .Q (new_AGEMA_signal_32623) ) ;
    buf_clk new_AGEMA_reg_buffer_11671 ( .C (clk), .D (new_AGEMA_signal_32626), .Q (new_AGEMA_signal_32627) ) ;
    buf_clk new_AGEMA_reg_buffer_11675 ( .C (clk), .D (new_AGEMA_signal_32630), .Q (new_AGEMA_signal_32631) ) ;
    buf_clk new_AGEMA_reg_buffer_11679 ( .C (clk), .D (new_AGEMA_signal_32634), .Q (new_AGEMA_signal_32635) ) ;
    buf_clk new_AGEMA_reg_buffer_11683 ( .C (clk), .D (new_AGEMA_signal_32638), .Q (new_AGEMA_signal_32639) ) ;
    buf_clk new_AGEMA_reg_buffer_11687 ( .C (clk), .D (new_AGEMA_signal_32642), .Q (new_AGEMA_signal_32643) ) ;
    buf_clk new_AGEMA_reg_buffer_11691 ( .C (clk), .D (new_AGEMA_signal_32646), .Q (new_AGEMA_signal_32647) ) ;
    buf_clk new_AGEMA_reg_buffer_11695 ( .C (clk), .D (new_AGEMA_signal_32650), .Q (new_AGEMA_signal_32651) ) ;
    buf_clk new_AGEMA_reg_buffer_11699 ( .C (clk), .D (new_AGEMA_signal_32654), .Q (new_AGEMA_signal_32655) ) ;
    buf_clk new_AGEMA_reg_buffer_11703 ( .C (clk), .D (new_AGEMA_signal_32658), .Q (new_AGEMA_signal_32659) ) ;
    buf_clk new_AGEMA_reg_buffer_11707 ( .C (clk), .D (new_AGEMA_signal_32662), .Q (new_AGEMA_signal_32663) ) ;
    buf_clk new_AGEMA_reg_buffer_11711 ( .C (clk), .D (new_AGEMA_signal_32666), .Q (new_AGEMA_signal_32667) ) ;
    buf_clk new_AGEMA_reg_buffer_11715 ( .C (clk), .D (new_AGEMA_signal_32670), .Q (new_AGEMA_signal_32671) ) ;
    buf_clk new_AGEMA_reg_buffer_11719 ( .C (clk), .D (new_AGEMA_signal_32674), .Q (new_AGEMA_signal_32675) ) ;
    buf_clk new_AGEMA_reg_buffer_11723 ( .C (clk), .D (new_AGEMA_signal_32678), .Q (new_AGEMA_signal_32679) ) ;
    buf_clk new_AGEMA_reg_buffer_11727 ( .C (clk), .D (new_AGEMA_signal_32682), .Q (new_AGEMA_signal_32683) ) ;
    buf_clk new_AGEMA_reg_buffer_11731 ( .C (clk), .D (new_AGEMA_signal_32686), .Q (new_AGEMA_signal_32687) ) ;
    buf_clk new_AGEMA_reg_buffer_11735 ( .C (clk), .D (new_AGEMA_signal_32690), .Q (new_AGEMA_signal_32691) ) ;
    buf_clk new_AGEMA_reg_buffer_11739 ( .C (clk), .D (new_AGEMA_signal_32694), .Q (new_AGEMA_signal_32695) ) ;
    buf_clk new_AGEMA_reg_buffer_11743 ( .C (clk), .D (new_AGEMA_signal_32698), .Q (new_AGEMA_signal_32699) ) ;
    buf_clk new_AGEMA_reg_buffer_11747 ( .C (clk), .D (new_AGEMA_signal_32702), .Q (new_AGEMA_signal_32703) ) ;
    buf_clk new_AGEMA_reg_buffer_11751 ( .C (clk), .D (new_AGEMA_signal_32706), .Q (new_AGEMA_signal_32707) ) ;
    buf_clk new_AGEMA_reg_buffer_11755 ( .C (clk), .D (new_AGEMA_signal_32710), .Q (new_AGEMA_signal_32711) ) ;
    buf_clk new_AGEMA_reg_buffer_11759 ( .C (clk), .D (new_AGEMA_signal_32714), .Q (new_AGEMA_signal_32715) ) ;
    buf_clk new_AGEMA_reg_buffer_11763 ( .C (clk), .D (new_AGEMA_signal_32718), .Q (new_AGEMA_signal_32719) ) ;
    buf_clk new_AGEMA_reg_buffer_11767 ( .C (clk), .D (new_AGEMA_signal_32722), .Q (new_AGEMA_signal_32723) ) ;
    buf_clk new_AGEMA_reg_buffer_11771 ( .C (clk), .D (new_AGEMA_signal_32726), .Q (new_AGEMA_signal_32727) ) ;
    buf_clk new_AGEMA_reg_buffer_11775 ( .C (clk), .D (new_AGEMA_signal_32730), .Q (new_AGEMA_signal_32731) ) ;
    buf_clk new_AGEMA_reg_buffer_11779 ( .C (clk), .D (new_AGEMA_signal_32734), .Q (new_AGEMA_signal_32735) ) ;
    buf_clk new_AGEMA_reg_buffer_11783 ( .C (clk), .D (new_AGEMA_signal_32738), .Q (new_AGEMA_signal_32739) ) ;
    buf_clk new_AGEMA_reg_buffer_11787 ( .C (clk), .D (new_AGEMA_signal_32742), .Q (new_AGEMA_signal_32743) ) ;
    buf_clk new_AGEMA_reg_buffer_11791 ( .C (clk), .D (new_AGEMA_signal_32746), .Q (new_AGEMA_signal_32747) ) ;
    buf_clk new_AGEMA_reg_buffer_11795 ( .C (clk), .D (new_AGEMA_signal_32750), .Q (new_AGEMA_signal_32751) ) ;
    buf_clk new_AGEMA_reg_buffer_11799 ( .C (clk), .D (new_AGEMA_signal_32754), .Q (new_AGEMA_signal_32755) ) ;
    buf_clk new_AGEMA_reg_buffer_11803 ( .C (clk), .D (new_AGEMA_signal_32758), .Q (new_AGEMA_signal_32759) ) ;
    buf_clk new_AGEMA_reg_buffer_11807 ( .C (clk), .D (new_AGEMA_signal_32762), .Q (new_AGEMA_signal_32763) ) ;
    buf_clk new_AGEMA_reg_buffer_11811 ( .C (clk), .D (new_AGEMA_signal_32766), .Q (new_AGEMA_signal_32767) ) ;
    buf_clk new_AGEMA_reg_buffer_11815 ( .C (clk), .D (new_AGEMA_signal_32770), .Q (new_AGEMA_signal_32771) ) ;
    buf_clk new_AGEMA_reg_buffer_11819 ( .C (clk), .D (new_AGEMA_signal_32774), .Q (new_AGEMA_signal_32775) ) ;
    buf_clk new_AGEMA_reg_buffer_11823 ( .C (clk), .D (new_AGEMA_signal_32778), .Q (new_AGEMA_signal_32779) ) ;
    buf_clk new_AGEMA_reg_buffer_11827 ( .C (clk), .D (new_AGEMA_signal_32782), .Q (new_AGEMA_signal_32783) ) ;
    buf_clk new_AGEMA_reg_buffer_11831 ( .C (clk), .D (new_AGEMA_signal_32786), .Q (new_AGEMA_signal_32787) ) ;
    buf_clk new_AGEMA_reg_buffer_11835 ( .C (clk), .D (new_AGEMA_signal_32790), .Q (new_AGEMA_signal_32791) ) ;
    buf_clk new_AGEMA_reg_buffer_11839 ( .C (clk), .D (new_AGEMA_signal_32794), .Q (new_AGEMA_signal_32795) ) ;
    buf_clk new_AGEMA_reg_buffer_11843 ( .C (clk), .D (new_AGEMA_signal_32798), .Q (new_AGEMA_signal_32799) ) ;
    buf_clk new_AGEMA_reg_buffer_11847 ( .C (clk), .D (new_AGEMA_signal_32802), .Q (new_AGEMA_signal_32803) ) ;
    buf_clk new_AGEMA_reg_buffer_11851 ( .C (clk), .D (new_AGEMA_signal_32806), .Q (new_AGEMA_signal_32807) ) ;
    buf_clk new_AGEMA_reg_buffer_11855 ( .C (clk), .D (new_AGEMA_signal_32810), .Q (new_AGEMA_signal_32811) ) ;
    buf_clk new_AGEMA_reg_buffer_11859 ( .C (clk), .D (new_AGEMA_signal_32814), .Q (new_AGEMA_signal_32815) ) ;
    buf_clk new_AGEMA_reg_buffer_11863 ( .C (clk), .D (new_AGEMA_signal_32818), .Q (new_AGEMA_signal_32819) ) ;
    buf_clk new_AGEMA_reg_buffer_11867 ( .C (clk), .D (new_AGEMA_signal_32822), .Q (new_AGEMA_signal_32823) ) ;
    buf_clk new_AGEMA_reg_buffer_11871 ( .C (clk), .D (new_AGEMA_signal_32826), .Q (new_AGEMA_signal_32827) ) ;
    buf_clk new_AGEMA_reg_buffer_11875 ( .C (clk), .D (new_AGEMA_signal_32830), .Q (new_AGEMA_signal_32831) ) ;
    buf_clk new_AGEMA_reg_buffer_11879 ( .C (clk), .D (new_AGEMA_signal_32834), .Q (new_AGEMA_signal_32835) ) ;
    buf_clk new_AGEMA_reg_buffer_11883 ( .C (clk), .D (new_AGEMA_signal_32838), .Q (new_AGEMA_signal_32839) ) ;
    buf_clk new_AGEMA_reg_buffer_11887 ( .C (clk), .D (new_AGEMA_signal_32842), .Q (new_AGEMA_signal_32843) ) ;
    buf_clk new_AGEMA_reg_buffer_11891 ( .C (clk), .D (new_AGEMA_signal_32846), .Q (new_AGEMA_signal_32847) ) ;
    buf_clk new_AGEMA_reg_buffer_11895 ( .C (clk), .D (new_AGEMA_signal_32850), .Q (new_AGEMA_signal_32851) ) ;
    buf_clk new_AGEMA_reg_buffer_11899 ( .C (clk), .D (new_AGEMA_signal_32854), .Q (new_AGEMA_signal_32855) ) ;
    buf_clk new_AGEMA_reg_buffer_11903 ( .C (clk), .D (new_AGEMA_signal_32858), .Q (new_AGEMA_signal_32859) ) ;
    buf_clk new_AGEMA_reg_buffer_11907 ( .C (clk), .D (new_AGEMA_signal_32862), .Q (new_AGEMA_signal_32863) ) ;
    buf_clk new_AGEMA_reg_buffer_11911 ( .C (clk), .D (new_AGEMA_signal_32866), .Q (new_AGEMA_signal_32867) ) ;
    buf_clk new_AGEMA_reg_buffer_11915 ( .C (clk), .D (new_AGEMA_signal_32870), .Q (new_AGEMA_signal_32871) ) ;
    buf_clk new_AGEMA_reg_buffer_11919 ( .C (clk), .D (new_AGEMA_signal_32874), .Q (new_AGEMA_signal_32875) ) ;
    buf_clk new_AGEMA_reg_buffer_11923 ( .C (clk), .D (new_AGEMA_signal_32878), .Q (new_AGEMA_signal_32879) ) ;
    buf_clk new_AGEMA_reg_buffer_11927 ( .C (clk), .D (new_AGEMA_signal_32882), .Q (new_AGEMA_signal_32883) ) ;
    buf_clk new_AGEMA_reg_buffer_11931 ( .C (clk), .D (new_AGEMA_signal_32886), .Q (new_AGEMA_signal_32887) ) ;
    buf_clk new_AGEMA_reg_buffer_11935 ( .C (clk), .D (new_AGEMA_signal_32890), .Q (new_AGEMA_signal_32891) ) ;
    buf_clk new_AGEMA_reg_buffer_11939 ( .C (clk), .D (new_AGEMA_signal_32894), .Q (new_AGEMA_signal_32895) ) ;
    buf_clk new_AGEMA_reg_buffer_11943 ( .C (clk), .D (new_AGEMA_signal_32898), .Q (new_AGEMA_signal_32899) ) ;
    buf_clk new_AGEMA_reg_buffer_11947 ( .C (clk), .D (new_AGEMA_signal_32902), .Q (new_AGEMA_signal_32903) ) ;
    buf_clk new_AGEMA_reg_buffer_11951 ( .C (clk), .D (new_AGEMA_signal_32906), .Q (new_AGEMA_signal_32907) ) ;
    buf_clk new_AGEMA_reg_buffer_11955 ( .C (clk), .D (new_AGEMA_signal_32910), .Q (new_AGEMA_signal_32911) ) ;
    buf_clk new_AGEMA_reg_buffer_11959 ( .C (clk), .D (new_AGEMA_signal_32914), .Q (new_AGEMA_signal_32915) ) ;
    buf_clk new_AGEMA_reg_buffer_11963 ( .C (clk), .D (new_AGEMA_signal_32918), .Q (new_AGEMA_signal_32919) ) ;
    buf_clk new_AGEMA_reg_buffer_11967 ( .C (clk), .D (new_AGEMA_signal_32922), .Q (new_AGEMA_signal_32923) ) ;
    buf_clk new_AGEMA_reg_buffer_11971 ( .C (clk), .D (new_AGEMA_signal_32926), .Q (new_AGEMA_signal_32927) ) ;
    buf_clk new_AGEMA_reg_buffer_11975 ( .C (clk), .D (new_AGEMA_signal_32930), .Q (new_AGEMA_signal_32931) ) ;
    buf_clk new_AGEMA_reg_buffer_11979 ( .C (clk), .D (new_AGEMA_signal_32934), .Q (new_AGEMA_signal_32935) ) ;
    buf_clk new_AGEMA_reg_buffer_11983 ( .C (clk), .D (new_AGEMA_signal_32938), .Q (new_AGEMA_signal_32939) ) ;
    buf_clk new_AGEMA_reg_buffer_11987 ( .C (clk), .D (new_AGEMA_signal_32942), .Q (new_AGEMA_signal_32943) ) ;
    buf_clk new_AGEMA_reg_buffer_11991 ( .C (clk), .D (new_AGEMA_signal_32946), .Q (new_AGEMA_signal_32947) ) ;
    buf_clk new_AGEMA_reg_buffer_11995 ( .C (clk), .D (new_AGEMA_signal_32950), .Q (new_AGEMA_signal_32951) ) ;
    buf_clk new_AGEMA_reg_buffer_11999 ( .C (clk), .D (new_AGEMA_signal_32954), .Q (new_AGEMA_signal_32955) ) ;
    buf_clk new_AGEMA_reg_buffer_12003 ( .C (clk), .D (new_AGEMA_signal_32958), .Q (new_AGEMA_signal_32959) ) ;
    buf_clk new_AGEMA_reg_buffer_12007 ( .C (clk), .D (new_AGEMA_signal_32962), .Q (new_AGEMA_signal_32963) ) ;
    buf_clk new_AGEMA_reg_buffer_12011 ( .C (clk), .D (new_AGEMA_signal_32966), .Q (new_AGEMA_signal_32967) ) ;
    buf_clk new_AGEMA_reg_buffer_12015 ( .C (clk), .D (new_AGEMA_signal_32970), .Q (new_AGEMA_signal_32971) ) ;
    buf_clk new_AGEMA_reg_buffer_12019 ( .C (clk), .D (new_AGEMA_signal_32974), .Q (new_AGEMA_signal_32975) ) ;
    buf_clk new_AGEMA_reg_buffer_12023 ( .C (clk), .D (new_AGEMA_signal_32978), .Q (new_AGEMA_signal_32979) ) ;
    buf_clk new_AGEMA_reg_buffer_12027 ( .C (clk), .D (new_AGEMA_signal_32982), .Q (new_AGEMA_signal_32983) ) ;
    buf_clk new_AGEMA_reg_buffer_12031 ( .C (clk), .D (new_AGEMA_signal_32986), .Q (new_AGEMA_signal_32987) ) ;
    buf_clk new_AGEMA_reg_buffer_12035 ( .C (clk), .D (new_AGEMA_signal_32990), .Q (new_AGEMA_signal_32991) ) ;
    buf_clk new_AGEMA_reg_buffer_12039 ( .C (clk), .D (new_AGEMA_signal_32994), .Q (new_AGEMA_signal_32995) ) ;
    buf_clk new_AGEMA_reg_buffer_12043 ( .C (clk), .D (new_AGEMA_signal_32998), .Q (new_AGEMA_signal_32999) ) ;
    buf_clk new_AGEMA_reg_buffer_12047 ( .C (clk), .D (new_AGEMA_signal_33002), .Q (new_AGEMA_signal_33003) ) ;
    buf_clk new_AGEMA_reg_buffer_12051 ( .C (clk), .D (new_AGEMA_signal_33006), .Q (new_AGEMA_signal_33007) ) ;
    buf_clk new_AGEMA_reg_buffer_12055 ( .C (clk), .D (new_AGEMA_signal_33010), .Q (new_AGEMA_signal_33011) ) ;
    buf_clk new_AGEMA_reg_buffer_12059 ( .C (clk), .D (new_AGEMA_signal_33014), .Q (new_AGEMA_signal_33015) ) ;
    buf_clk new_AGEMA_reg_buffer_12063 ( .C (clk), .D (new_AGEMA_signal_33018), .Q (new_AGEMA_signal_33019) ) ;
    buf_clk new_AGEMA_reg_buffer_12067 ( .C (clk), .D (new_AGEMA_signal_33022), .Q (new_AGEMA_signal_33023) ) ;
    buf_clk new_AGEMA_reg_buffer_12071 ( .C (clk), .D (new_AGEMA_signal_33026), .Q (new_AGEMA_signal_33027) ) ;
    buf_clk new_AGEMA_reg_buffer_12075 ( .C (clk), .D (new_AGEMA_signal_33030), .Q (new_AGEMA_signal_33031) ) ;
    buf_clk new_AGEMA_reg_buffer_12079 ( .C (clk), .D (new_AGEMA_signal_33034), .Q (new_AGEMA_signal_33035) ) ;
    buf_clk new_AGEMA_reg_buffer_12083 ( .C (clk), .D (new_AGEMA_signal_33038), .Q (new_AGEMA_signal_33039) ) ;
    buf_clk new_AGEMA_reg_buffer_12087 ( .C (clk), .D (new_AGEMA_signal_33042), .Q (new_AGEMA_signal_33043) ) ;
    buf_clk new_AGEMA_reg_buffer_12091 ( .C (clk), .D (new_AGEMA_signal_33046), .Q (new_AGEMA_signal_33047) ) ;
    buf_clk new_AGEMA_reg_buffer_12095 ( .C (clk), .D (new_AGEMA_signal_33050), .Q (new_AGEMA_signal_33051) ) ;
    buf_clk new_AGEMA_reg_buffer_12099 ( .C (clk), .D (new_AGEMA_signal_33054), .Q (new_AGEMA_signal_33055) ) ;
    buf_clk new_AGEMA_reg_buffer_12103 ( .C (clk), .D (new_AGEMA_signal_33058), .Q (new_AGEMA_signal_33059) ) ;
    buf_clk new_AGEMA_reg_buffer_12107 ( .C (clk), .D (new_AGEMA_signal_33062), .Q (new_AGEMA_signal_33063) ) ;
    buf_clk new_AGEMA_reg_buffer_12111 ( .C (clk), .D (new_AGEMA_signal_33066), .Q (new_AGEMA_signal_33067) ) ;
    buf_clk new_AGEMA_reg_buffer_12115 ( .C (clk), .D (new_AGEMA_signal_33070), .Q (new_AGEMA_signal_33071) ) ;
    buf_clk new_AGEMA_reg_buffer_12119 ( .C (clk), .D (new_AGEMA_signal_33074), .Q (new_AGEMA_signal_33075) ) ;
    buf_clk new_AGEMA_reg_buffer_12123 ( .C (clk), .D (new_AGEMA_signal_33078), .Q (new_AGEMA_signal_33079) ) ;
    buf_clk new_AGEMA_reg_buffer_12127 ( .C (clk), .D (new_AGEMA_signal_33082), .Q (new_AGEMA_signal_33083) ) ;
    buf_clk new_AGEMA_reg_buffer_12131 ( .C (clk), .D (new_AGEMA_signal_33086), .Q (new_AGEMA_signal_33087) ) ;
    buf_clk new_AGEMA_reg_buffer_12135 ( .C (clk), .D (new_AGEMA_signal_33090), .Q (new_AGEMA_signal_33091) ) ;
    buf_clk new_AGEMA_reg_buffer_12139 ( .C (clk), .D (new_AGEMA_signal_33094), .Q (new_AGEMA_signal_33095) ) ;
    buf_clk new_AGEMA_reg_buffer_12143 ( .C (clk), .D (new_AGEMA_signal_33098), .Q (new_AGEMA_signal_33099) ) ;
    buf_clk new_AGEMA_reg_buffer_12147 ( .C (clk), .D (new_AGEMA_signal_33102), .Q (new_AGEMA_signal_33103) ) ;
    buf_clk new_AGEMA_reg_buffer_12151 ( .C (clk), .D (new_AGEMA_signal_33106), .Q (new_AGEMA_signal_33107) ) ;
    buf_clk new_AGEMA_reg_buffer_12155 ( .C (clk), .D (new_AGEMA_signal_33110), .Q (new_AGEMA_signal_33111) ) ;
    buf_clk new_AGEMA_reg_buffer_12159 ( .C (clk), .D (new_AGEMA_signal_33114), .Q (new_AGEMA_signal_33115) ) ;
    buf_clk new_AGEMA_reg_buffer_12163 ( .C (clk), .D (new_AGEMA_signal_33118), .Q (new_AGEMA_signal_33119) ) ;
    buf_clk new_AGEMA_reg_buffer_12167 ( .C (clk), .D (new_AGEMA_signal_33122), .Q (new_AGEMA_signal_33123) ) ;
    buf_clk new_AGEMA_reg_buffer_12171 ( .C (clk), .D (new_AGEMA_signal_33126), .Q (new_AGEMA_signal_33127) ) ;
    buf_clk new_AGEMA_reg_buffer_12175 ( .C (clk), .D (new_AGEMA_signal_33130), .Q (new_AGEMA_signal_33131) ) ;
    buf_clk new_AGEMA_reg_buffer_12179 ( .C (clk), .D (new_AGEMA_signal_33134), .Q (new_AGEMA_signal_33135) ) ;
    buf_clk new_AGEMA_reg_buffer_12183 ( .C (clk), .D (new_AGEMA_signal_33138), .Q (new_AGEMA_signal_33139) ) ;
    buf_clk new_AGEMA_reg_buffer_12187 ( .C (clk), .D (new_AGEMA_signal_33142), .Q (new_AGEMA_signal_33143) ) ;
    buf_clk new_AGEMA_reg_buffer_12191 ( .C (clk), .D (new_AGEMA_signal_33146), .Q (new_AGEMA_signal_33147) ) ;
    buf_clk new_AGEMA_reg_buffer_12195 ( .C (clk), .D (new_AGEMA_signal_33150), .Q (new_AGEMA_signal_33151) ) ;
    buf_clk new_AGEMA_reg_buffer_12199 ( .C (clk), .D (new_AGEMA_signal_33154), .Q (new_AGEMA_signal_33155) ) ;
    buf_clk new_AGEMA_reg_buffer_12203 ( .C (clk), .D (new_AGEMA_signal_33158), .Q (new_AGEMA_signal_33159) ) ;
    buf_clk new_AGEMA_reg_buffer_12207 ( .C (clk), .D (new_AGEMA_signal_33162), .Q (new_AGEMA_signal_33163) ) ;
    buf_clk new_AGEMA_reg_buffer_12211 ( .C (clk), .D (new_AGEMA_signal_33166), .Q (new_AGEMA_signal_33167) ) ;
    buf_clk new_AGEMA_reg_buffer_12215 ( .C (clk), .D (new_AGEMA_signal_33170), .Q (new_AGEMA_signal_33171) ) ;
    buf_clk new_AGEMA_reg_buffer_12219 ( .C (clk), .D (new_AGEMA_signal_33174), .Q (new_AGEMA_signal_33175) ) ;
    buf_clk new_AGEMA_reg_buffer_12223 ( .C (clk), .D (new_AGEMA_signal_33178), .Q (new_AGEMA_signal_33179) ) ;
    buf_clk new_AGEMA_reg_buffer_12227 ( .C (clk), .D (new_AGEMA_signal_33182), .Q (new_AGEMA_signal_33183) ) ;
    buf_clk new_AGEMA_reg_buffer_12231 ( .C (clk), .D (new_AGEMA_signal_33186), .Q (new_AGEMA_signal_33187) ) ;
    buf_clk new_AGEMA_reg_buffer_12235 ( .C (clk), .D (new_AGEMA_signal_33190), .Q (new_AGEMA_signal_33191) ) ;
    buf_clk new_AGEMA_reg_buffer_12239 ( .C (clk), .D (new_AGEMA_signal_33194), .Q (new_AGEMA_signal_33195) ) ;
    buf_clk new_AGEMA_reg_buffer_12243 ( .C (clk), .D (new_AGEMA_signal_33198), .Q (new_AGEMA_signal_33199) ) ;
    buf_clk new_AGEMA_reg_buffer_12247 ( .C (clk), .D (new_AGEMA_signal_33202), .Q (new_AGEMA_signal_33203) ) ;
    buf_clk new_AGEMA_reg_buffer_12251 ( .C (clk), .D (new_AGEMA_signal_33206), .Q (new_AGEMA_signal_33207) ) ;
    buf_clk new_AGEMA_reg_buffer_12255 ( .C (clk), .D (new_AGEMA_signal_33210), .Q (new_AGEMA_signal_33211) ) ;
    buf_clk new_AGEMA_reg_buffer_12259 ( .C (clk), .D (new_AGEMA_signal_33214), .Q (new_AGEMA_signal_33215) ) ;
    buf_clk new_AGEMA_reg_buffer_12263 ( .C (clk), .D (new_AGEMA_signal_33218), .Q (new_AGEMA_signal_33219) ) ;
    buf_clk new_AGEMA_reg_buffer_12267 ( .C (clk), .D (new_AGEMA_signal_33222), .Q (new_AGEMA_signal_33223) ) ;
    buf_clk new_AGEMA_reg_buffer_12271 ( .C (clk), .D (new_AGEMA_signal_33226), .Q (new_AGEMA_signal_33227) ) ;
    buf_clk new_AGEMA_reg_buffer_12275 ( .C (clk), .D (new_AGEMA_signal_33230), .Q (new_AGEMA_signal_33231) ) ;
    buf_clk new_AGEMA_reg_buffer_12279 ( .C (clk), .D (new_AGEMA_signal_33234), .Q (new_AGEMA_signal_33235) ) ;
    buf_clk new_AGEMA_reg_buffer_12283 ( .C (clk), .D (new_AGEMA_signal_33238), .Q (new_AGEMA_signal_33239) ) ;
    buf_clk new_AGEMA_reg_buffer_12287 ( .C (clk), .D (new_AGEMA_signal_33242), .Q (new_AGEMA_signal_33243) ) ;
    buf_clk new_AGEMA_reg_buffer_12291 ( .C (clk), .D (new_AGEMA_signal_33246), .Q (new_AGEMA_signal_33247) ) ;
    buf_clk new_AGEMA_reg_buffer_12295 ( .C (clk), .D (new_AGEMA_signal_33250), .Q (new_AGEMA_signal_33251) ) ;
    buf_clk new_AGEMA_reg_buffer_12299 ( .C (clk), .D (new_AGEMA_signal_33254), .Q (new_AGEMA_signal_33255) ) ;
    buf_clk new_AGEMA_reg_buffer_12303 ( .C (clk), .D (new_AGEMA_signal_33258), .Q (new_AGEMA_signal_33259) ) ;
    buf_clk new_AGEMA_reg_buffer_12307 ( .C (clk), .D (new_AGEMA_signal_33262), .Q (new_AGEMA_signal_33263) ) ;
    buf_clk new_AGEMA_reg_buffer_12311 ( .C (clk), .D (new_AGEMA_signal_33266), .Q (new_AGEMA_signal_33267) ) ;
    buf_clk new_AGEMA_reg_buffer_12315 ( .C (clk), .D (new_AGEMA_signal_33270), .Q (new_AGEMA_signal_33271) ) ;
    buf_clk new_AGEMA_reg_buffer_12319 ( .C (clk), .D (new_AGEMA_signal_33274), .Q (new_AGEMA_signal_33275) ) ;
    buf_clk new_AGEMA_reg_buffer_12323 ( .C (clk), .D (new_AGEMA_signal_33278), .Q (new_AGEMA_signal_33279) ) ;
    buf_clk new_AGEMA_reg_buffer_12327 ( .C (clk), .D (new_AGEMA_signal_33282), .Q (new_AGEMA_signal_33283) ) ;
    buf_clk new_AGEMA_reg_buffer_12331 ( .C (clk), .D (new_AGEMA_signal_33286), .Q (new_AGEMA_signal_33287) ) ;
    buf_clk new_AGEMA_reg_buffer_12335 ( .C (clk), .D (new_AGEMA_signal_33290), .Q (new_AGEMA_signal_33291) ) ;
    buf_clk new_AGEMA_reg_buffer_12339 ( .C (clk), .D (new_AGEMA_signal_33294), .Q (new_AGEMA_signal_33295) ) ;
    buf_clk new_AGEMA_reg_buffer_12343 ( .C (clk), .D (new_AGEMA_signal_33298), .Q (new_AGEMA_signal_33299) ) ;
    buf_clk new_AGEMA_reg_buffer_12347 ( .C (clk), .D (new_AGEMA_signal_33302), .Q (new_AGEMA_signal_33303) ) ;
    buf_clk new_AGEMA_reg_buffer_12351 ( .C (clk), .D (new_AGEMA_signal_33306), .Q (new_AGEMA_signal_33307) ) ;
    buf_clk new_AGEMA_reg_buffer_12355 ( .C (clk), .D (new_AGEMA_signal_33310), .Q (new_AGEMA_signal_33311) ) ;
    buf_clk new_AGEMA_reg_buffer_12359 ( .C (clk), .D (new_AGEMA_signal_33314), .Q (new_AGEMA_signal_33315) ) ;
    buf_clk new_AGEMA_reg_buffer_12363 ( .C (clk), .D (new_AGEMA_signal_33318), .Q (new_AGEMA_signal_33319) ) ;
    buf_clk new_AGEMA_reg_buffer_12367 ( .C (clk), .D (new_AGEMA_signal_33322), .Q (new_AGEMA_signal_33323) ) ;
    buf_clk new_AGEMA_reg_buffer_12371 ( .C (clk), .D (new_AGEMA_signal_33326), .Q (new_AGEMA_signal_33327) ) ;
    buf_clk new_AGEMA_reg_buffer_12375 ( .C (clk), .D (new_AGEMA_signal_33330), .Q (new_AGEMA_signal_33331) ) ;
    buf_clk new_AGEMA_reg_buffer_12379 ( .C (clk), .D (new_AGEMA_signal_33334), .Q (new_AGEMA_signal_33335) ) ;
    buf_clk new_AGEMA_reg_buffer_12383 ( .C (clk), .D (new_AGEMA_signal_33338), .Q (new_AGEMA_signal_33339) ) ;
    buf_clk new_AGEMA_reg_buffer_12387 ( .C (clk), .D (new_AGEMA_signal_33342), .Q (new_AGEMA_signal_33343) ) ;
    buf_clk new_AGEMA_reg_buffer_12391 ( .C (clk), .D (new_AGEMA_signal_33346), .Q (new_AGEMA_signal_33347) ) ;
    buf_clk new_AGEMA_reg_buffer_12395 ( .C (clk), .D (new_AGEMA_signal_33350), .Q (new_AGEMA_signal_33351) ) ;
    buf_clk new_AGEMA_reg_buffer_12399 ( .C (clk), .D (new_AGEMA_signal_33354), .Q (new_AGEMA_signal_33355) ) ;
    buf_clk new_AGEMA_reg_buffer_12403 ( .C (clk), .D (new_AGEMA_signal_33358), .Q (new_AGEMA_signal_33359) ) ;
    buf_clk new_AGEMA_reg_buffer_12407 ( .C (clk), .D (new_AGEMA_signal_33362), .Q (new_AGEMA_signal_33363) ) ;
    buf_clk new_AGEMA_reg_buffer_12411 ( .C (clk), .D (new_AGEMA_signal_33366), .Q (new_AGEMA_signal_33367) ) ;
    buf_clk new_AGEMA_reg_buffer_12415 ( .C (clk), .D (new_AGEMA_signal_33370), .Q (new_AGEMA_signal_33371) ) ;
    buf_clk new_AGEMA_reg_buffer_12419 ( .C (clk), .D (new_AGEMA_signal_33374), .Q (new_AGEMA_signal_33375) ) ;
    buf_clk new_AGEMA_reg_buffer_12423 ( .C (clk), .D (new_AGEMA_signal_33378), .Q (new_AGEMA_signal_33379) ) ;
    buf_clk new_AGEMA_reg_buffer_12427 ( .C (clk), .D (new_AGEMA_signal_33382), .Q (new_AGEMA_signal_33383) ) ;
    buf_clk new_AGEMA_reg_buffer_12431 ( .C (clk), .D (new_AGEMA_signal_33386), .Q (new_AGEMA_signal_33387) ) ;
    buf_clk new_AGEMA_reg_buffer_12435 ( .C (clk), .D (new_AGEMA_signal_33390), .Q (new_AGEMA_signal_33391) ) ;
    buf_clk new_AGEMA_reg_buffer_12439 ( .C (clk), .D (new_AGEMA_signal_33394), .Q (new_AGEMA_signal_33395) ) ;
    buf_clk new_AGEMA_reg_buffer_12443 ( .C (clk), .D (new_AGEMA_signal_33398), .Q (new_AGEMA_signal_33399) ) ;
    buf_clk new_AGEMA_reg_buffer_12447 ( .C (clk), .D (new_AGEMA_signal_33402), .Q (new_AGEMA_signal_33403) ) ;
    buf_clk new_AGEMA_reg_buffer_12451 ( .C (clk), .D (new_AGEMA_signal_33406), .Q (new_AGEMA_signal_33407) ) ;
    buf_clk new_AGEMA_reg_buffer_12455 ( .C (clk), .D (new_AGEMA_signal_33410), .Q (new_AGEMA_signal_33411) ) ;
    buf_clk new_AGEMA_reg_buffer_12459 ( .C (clk), .D (new_AGEMA_signal_33414), .Q (new_AGEMA_signal_33415) ) ;
    buf_clk new_AGEMA_reg_buffer_12463 ( .C (clk), .D (new_AGEMA_signal_33418), .Q (new_AGEMA_signal_33419) ) ;
    buf_clk new_AGEMA_reg_buffer_12467 ( .C (clk), .D (new_AGEMA_signal_33422), .Q (new_AGEMA_signal_33423) ) ;
    buf_clk new_AGEMA_reg_buffer_12471 ( .C (clk), .D (new_AGEMA_signal_33426), .Q (new_AGEMA_signal_33427) ) ;
    buf_clk new_AGEMA_reg_buffer_12475 ( .C (clk), .D (new_AGEMA_signal_33430), .Q (new_AGEMA_signal_33431) ) ;
    buf_clk new_AGEMA_reg_buffer_12479 ( .C (clk), .D (new_AGEMA_signal_33434), .Q (new_AGEMA_signal_33435) ) ;
    buf_clk new_AGEMA_reg_buffer_12483 ( .C (clk), .D (new_AGEMA_signal_33438), .Q (new_AGEMA_signal_33439) ) ;
    buf_clk new_AGEMA_reg_buffer_12487 ( .C (clk), .D (new_AGEMA_signal_33442), .Q (new_AGEMA_signal_33443) ) ;
    buf_clk new_AGEMA_reg_buffer_12491 ( .C (clk), .D (new_AGEMA_signal_33446), .Q (new_AGEMA_signal_33447) ) ;
    buf_clk new_AGEMA_reg_buffer_12495 ( .C (clk), .D (new_AGEMA_signal_33450), .Q (new_AGEMA_signal_33451) ) ;
    buf_clk new_AGEMA_reg_buffer_12499 ( .C (clk), .D (new_AGEMA_signal_33454), .Q (new_AGEMA_signal_33455) ) ;
    buf_clk new_AGEMA_reg_buffer_12503 ( .C (clk), .D (new_AGEMA_signal_33458), .Q (new_AGEMA_signal_33459) ) ;
    buf_clk new_AGEMA_reg_buffer_12507 ( .C (clk), .D (new_AGEMA_signal_33462), .Q (new_AGEMA_signal_33463) ) ;
    buf_clk new_AGEMA_reg_buffer_12511 ( .C (clk), .D (new_AGEMA_signal_33466), .Q (new_AGEMA_signal_33467) ) ;
    buf_clk new_AGEMA_reg_buffer_12515 ( .C (clk), .D (new_AGEMA_signal_33470), .Q (new_AGEMA_signal_33471) ) ;
    buf_clk new_AGEMA_reg_buffer_12519 ( .C (clk), .D (new_AGEMA_signal_33474), .Q (new_AGEMA_signal_33475) ) ;
    buf_clk new_AGEMA_reg_buffer_12523 ( .C (clk), .D (new_AGEMA_signal_33478), .Q (new_AGEMA_signal_33479) ) ;
    buf_clk new_AGEMA_reg_buffer_12527 ( .C (clk), .D (new_AGEMA_signal_33482), .Q (new_AGEMA_signal_33483) ) ;
    buf_clk new_AGEMA_reg_buffer_12531 ( .C (clk), .D (new_AGEMA_signal_33486), .Q (new_AGEMA_signal_33487) ) ;
    buf_clk new_AGEMA_reg_buffer_12535 ( .C (clk), .D (new_AGEMA_signal_33490), .Q (new_AGEMA_signal_33491) ) ;
    buf_clk new_AGEMA_reg_buffer_12539 ( .C (clk), .D (new_AGEMA_signal_33494), .Q (new_AGEMA_signal_33495) ) ;
    buf_clk new_AGEMA_reg_buffer_12543 ( .C (clk), .D (new_AGEMA_signal_33498), .Q (new_AGEMA_signal_33499) ) ;
    buf_clk new_AGEMA_reg_buffer_12547 ( .C (clk), .D (new_AGEMA_signal_33502), .Q (new_AGEMA_signal_33503) ) ;
    buf_clk new_AGEMA_reg_buffer_12551 ( .C (clk), .D (new_AGEMA_signal_33506), .Q (new_AGEMA_signal_33507) ) ;
    buf_clk new_AGEMA_reg_buffer_12555 ( .C (clk), .D (new_AGEMA_signal_33510), .Q (new_AGEMA_signal_33511) ) ;
    buf_clk new_AGEMA_reg_buffer_12559 ( .C (clk), .D (new_AGEMA_signal_33514), .Q (new_AGEMA_signal_33515) ) ;
    buf_clk new_AGEMA_reg_buffer_12563 ( .C (clk), .D (new_AGEMA_signal_33518), .Q (new_AGEMA_signal_33519) ) ;
    buf_clk new_AGEMA_reg_buffer_12567 ( .C (clk), .D (new_AGEMA_signal_33522), .Q (new_AGEMA_signal_33523) ) ;
    buf_clk new_AGEMA_reg_buffer_12571 ( .C (clk), .D (new_AGEMA_signal_33526), .Q (new_AGEMA_signal_33527) ) ;
    buf_clk new_AGEMA_reg_buffer_12575 ( .C (clk), .D (new_AGEMA_signal_33530), .Q (new_AGEMA_signal_33531) ) ;
    buf_clk new_AGEMA_reg_buffer_12579 ( .C (clk), .D (new_AGEMA_signal_33534), .Q (new_AGEMA_signal_33535) ) ;
    buf_clk new_AGEMA_reg_buffer_12583 ( .C (clk), .D (new_AGEMA_signal_33538), .Q (new_AGEMA_signal_33539) ) ;
    buf_clk new_AGEMA_reg_buffer_12587 ( .C (clk), .D (new_AGEMA_signal_33542), .Q (new_AGEMA_signal_33543) ) ;
    buf_clk new_AGEMA_reg_buffer_12591 ( .C (clk), .D (new_AGEMA_signal_33546), .Q (new_AGEMA_signal_33547) ) ;
    buf_clk new_AGEMA_reg_buffer_12595 ( .C (clk), .D (new_AGEMA_signal_33550), .Q (new_AGEMA_signal_33551) ) ;
    buf_clk new_AGEMA_reg_buffer_12599 ( .C (clk), .D (new_AGEMA_signal_33554), .Q (new_AGEMA_signal_33555) ) ;
    buf_clk new_AGEMA_reg_buffer_12603 ( .C (clk), .D (new_AGEMA_signal_33558), .Q (new_AGEMA_signal_33559) ) ;
    buf_clk new_AGEMA_reg_buffer_12607 ( .C (clk), .D (new_AGEMA_signal_33562), .Q (new_AGEMA_signal_33563) ) ;
    buf_clk new_AGEMA_reg_buffer_12611 ( .C (clk), .D (new_AGEMA_signal_33566), .Q (new_AGEMA_signal_33567) ) ;
    buf_clk new_AGEMA_reg_buffer_12615 ( .C (clk), .D (new_AGEMA_signal_33570), .Q (new_AGEMA_signal_33571) ) ;
    buf_clk new_AGEMA_reg_buffer_12619 ( .C (clk), .D (new_AGEMA_signal_33574), .Q (new_AGEMA_signal_33575) ) ;
    buf_clk new_AGEMA_reg_buffer_12623 ( .C (clk), .D (new_AGEMA_signal_33578), .Q (new_AGEMA_signal_33579) ) ;
    buf_clk new_AGEMA_reg_buffer_12627 ( .C (clk), .D (new_AGEMA_signal_33582), .Q (new_AGEMA_signal_33583) ) ;
    buf_clk new_AGEMA_reg_buffer_12631 ( .C (clk), .D (new_AGEMA_signal_33586), .Q (new_AGEMA_signal_33587) ) ;
    buf_clk new_AGEMA_reg_buffer_12635 ( .C (clk), .D (new_AGEMA_signal_33590), .Q (new_AGEMA_signal_33591) ) ;
    buf_clk new_AGEMA_reg_buffer_12639 ( .C (clk), .D (new_AGEMA_signal_33594), .Q (new_AGEMA_signal_33595) ) ;
    buf_clk new_AGEMA_reg_buffer_12643 ( .C (clk), .D (new_AGEMA_signal_33598), .Q (new_AGEMA_signal_33599) ) ;
    buf_clk new_AGEMA_reg_buffer_12647 ( .C (clk), .D (new_AGEMA_signal_33602), .Q (new_AGEMA_signal_33603) ) ;
    buf_clk new_AGEMA_reg_buffer_12651 ( .C (clk), .D (new_AGEMA_signal_33606), .Q (new_AGEMA_signal_33607) ) ;
    buf_clk new_AGEMA_reg_buffer_12655 ( .C (clk), .D (new_AGEMA_signal_33610), .Q (new_AGEMA_signal_33611) ) ;
    buf_clk new_AGEMA_reg_buffer_12659 ( .C (clk), .D (new_AGEMA_signal_33614), .Q (new_AGEMA_signal_33615) ) ;
    buf_clk new_AGEMA_reg_buffer_12663 ( .C (clk), .D (new_AGEMA_signal_33618), .Q (new_AGEMA_signal_33619) ) ;
    buf_clk new_AGEMA_reg_buffer_12667 ( .C (clk), .D (new_AGEMA_signal_33622), .Q (new_AGEMA_signal_33623) ) ;
    buf_clk new_AGEMA_reg_buffer_12671 ( .C (clk), .D (new_AGEMA_signal_33626), .Q (new_AGEMA_signal_33627) ) ;
    buf_clk new_AGEMA_reg_buffer_12675 ( .C (clk), .D (new_AGEMA_signal_33630), .Q (new_AGEMA_signal_33631) ) ;
    buf_clk new_AGEMA_reg_buffer_12679 ( .C (clk), .D (new_AGEMA_signal_33634), .Q (new_AGEMA_signal_33635) ) ;
    buf_clk new_AGEMA_reg_buffer_12683 ( .C (clk), .D (new_AGEMA_signal_33638), .Q (new_AGEMA_signal_33639) ) ;
    buf_clk new_AGEMA_reg_buffer_12687 ( .C (clk), .D (new_AGEMA_signal_33642), .Q (new_AGEMA_signal_33643) ) ;
    buf_clk new_AGEMA_reg_buffer_12691 ( .C (clk), .D (new_AGEMA_signal_33646), .Q (new_AGEMA_signal_33647) ) ;
    buf_clk new_AGEMA_reg_buffer_12695 ( .C (clk), .D (new_AGEMA_signal_33650), .Q (new_AGEMA_signal_33651) ) ;
    buf_clk new_AGEMA_reg_buffer_12699 ( .C (clk), .D (new_AGEMA_signal_33654), .Q (new_AGEMA_signal_33655) ) ;
    buf_clk new_AGEMA_reg_buffer_12703 ( .C (clk), .D (new_AGEMA_signal_33658), .Q (new_AGEMA_signal_33659) ) ;
    buf_clk new_AGEMA_reg_buffer_12707 ( .C (clk), .D (new_AGEMA_signal_33662), .Q (new_AGEMA_signal_33663) ) ;
    buf_clk new_AGEMA_reg_buffer_12711 ( .C (clk), .D (new_AGEMA_signal_33666), .Q (new_AGEMA_signal_33667) ) ;
    buf_clk new_AGEMA_reg_buffer_12715 ( .C (clk), .D (new_AGEMA_signal_33670), .Q (new_AGEMA_signal_33671) ) ;
    buf_clk new_AGEMA_reg_buffer_12719 ( .C (clk), .D (new_AGEMA_signal_33674), .Q (new_AGEMA_signal_33675) ) ;
    buf_clk new_AGEMA_reg_buffer_12723 ( .C (clk), .D (new_AGEMA_signal_33678), .Q (new_AGEMA_signal_33679) ) ;
    buf_clk new_AGEMA_reg_buffer_12727 ( .C (clk), .D (new_AGEMA_signal_33682), .Q (new_AGEMA_signal_33683) ) ;
    buf_clk new_AGEMA_reg_buffer_12731 ( .C (clk), .D (new_AGEMA_signal_33686), .Q (new_AGEMA_signal_33687) ) ;
    buf_clk new_AGEMA_reg_buffer_12735 ( .C (clk), .D (new_AGEMA_signal_33690), .Q (new_AGEMA_signal_33691) ) ;
    buf_clk new_AGEMA_reg_buffer_12739 ( .C (clk), .D (new_AGEMA_signal_33694), .Q (new_AGEMA_signal_33695) ) ;
    buf_clk new_AGEMA_reg_buffer_12743 ( .C (clk), .D (new_AGEMA_signal_33698), .Q (new_AGEMA_signal_33699) ) ;
    buf_clk new_AGEMA_reg_buffer_12747 ( .C (clk), .D (new_AGEMA_signal_33702), .Q (new_AGEMA_signal_33703) ) ;
    buf_clk new_AGEMA_reg_buffer_12751 ( .C (clk), .D (new_AGEMA_signal_33706), .Q (new_AGEMA_signal_33707) ) ;
    buf_clk new_AGEMA_reg_buffer_12755 ( .C (clk), .D (new_AGEMA_signal_33710), .Q (new_AGEMA_signal_33711) ) ;
    buf_clk new_AGEMA_reg_buffer_12759 ( .C (clk), .D (new_AGEMA_signal_33714), .Q (new_AGEMA_signal_33715) ) ;
    buf_clk new_AGEMA_reg_buffer_12763 ( .C (clk), .D (new_AGEMA_signal_33718), .Q (new_AGEMA_signal_33719) ) ;
    buf_clk new_AGEMA_reg_buffer_12767 ( .C (clk), .D (new_AGEMA_signal_33722), .Q (new_AGEMA_signal_33723) ) ;
    buf_clk new_AGEMA_reg_buffer_12771 ( .C (clk), .D (new_AGEMA_signal_33726), .Q (new_AGEMA_signal_33727) ) ;
    buf_clk new_AGEMA_reg_buffer_12775 ( .C (clk), .D (new_AGEMA_signal_33730), .Q (new_AGEMA_signal_33731) ) ;
    buf_clk new_AGEMA_reg_buffer_12779 ( .C (clk), .D (new_AGEMA_signal_33734), .Q (new_AGEMA_signal_33735) ) ;
    buf_clk new_AGEMA_reg_buffer_12783 ( .C (clk), .D (new_AGEMA_signal_33738), .Q (new_AGEMA_signal_33739) ) ;
    buf_clk new_AGEMA_reg_buffer_12787 ( .C (clk), .D (new_AGEMA_signal_33742), .Q (new_AGEMA_signal_33743) ) ;
    buf_clk new_AGEMA_reg_buffer_12791 ( .C (clk), .D (new_AGEMA_signal_33746), .Q (new_AGEMA_signal_33747) ) ;
    buf_clk new_AGEMA_reg_buffer_12795 ( .C (clk), .D (new_AGEMA_signal_33750), .Q (new_AGEMA_signal_33751) ) ;
    buf_clk new_AGEMA_reg_buffer_12799 ( .C (clk), .D (new_AGEMA_signal_33754), .Q (new_AGEMA_signal_33755) ) ;
    buf_clk new_AGEMA_reg_buffer_12803 ( .C (clk), .D (new_AGEMA_signal_33758), .Q (new_AGEMA_signal_33759) ) ;
    buf_clk new_AGEMA_reg_buffer_12807 ( .C (clk), .D (new_AGEMA_signal_33762), .Q (new_AGEMA_signal_33763) ) ;
    buf_clk new_AGEMA_reg_buffer_12811 ( .C (clk), .D (new_AGEMA_signal_33766), .Q (new_AGEMA_signal_33767) ) ;
    buf_clk new_AGEMA_reg_buffer_12815 ( .C (clk), .D (new_AGEMA_signal_33770), .Q (new_AGEMA_signal_33771) ) ;
    buf_clk new_AGEMA_reg_buffer_12819 ( .C (clk), .D (new_AGEMA_signal_33774), .Q (new_AGEMA_signal_33775) ) ;
    buf_clk new_AGEMA_reg_buffer_12823 ( .C (clk), .D (new_AGEMA_signal_33778), .Q (new_AGEMA_signal_33779) ) ;
    buf_clk new_AGEMA_reg_buffer_12827 ( .C (clk), .D (new_AGEMA_signal_33782), .Q (new_AGEMA_signal_33783) ) ;
    buf_clk new_AGEMA_reg_buffer_12831 ( .C (clk), .D (new_AGEMA_signal_33786), .Q (new_AGEMA_signal_33787) ) ;
    buf_clk new_AGEMA_reg_buffer_12835 ( .C (clk), .D (new_AGEMA_signal_33790), .Q (new_AGEMA_signal_33791) ) ;
    buf_clk new_AGEMA_reg_buffer_12839 ( .C (clk), .D (new_AGEMA_signal_33794), .Q (new_AGEMA_signal_33795) ) ;
    buf_clk new_AGEMA_reg_buffer_12843 ( .C (clk), .D (new_AGEMA_signal_33798), .Q (new_AGEMA_signal_33799) ) ;
    buf_clk new_AGEMA_reg_buffer_12847 ( .C (clk), .D (new_AGEMA_signal_33802), .Q (new_AGEMA_signal_33803) ) ;
    buf_clk new_AGEMA_reg_buffer_12851 ( .C (clk), .D (new_AGEMA_signal_33806), .Q (new_AGEMA_signal_33807) ) ;
    buf_clk new_AGEMA_reg_buffer_12855 ( .C (clk), .D (new_AGEMA_signal_33810), .Q (new_AGEMA_signal_33811) ) ;
    buf_clk new_AGEMA_reg_buffer_12859 ( .C (clk), .D (new_AGEMA_signal_33814), .Q (new_AGEMA_signal_33815) ) ;
    buf_clk new_AGEMA_reg_buffer_12863 ( .C (clk), .D (new_AGEMA_signal_33818), .Q (new_AGEMA_signal_33819) ) ;
    buf_clk new_AGEMA_reg_buffer_12867 ( .C (clk), .D (new_AGEMA_signal_33822), .Q (new_AGEMA_signal_33823) ) ;
    buf_clk new_AGEMA_reg_buffer_12871 ( .C (clk), .D (new_AGEMA_signal_33826), .Q (new_AGEMA_signal_33827) ) ;
    buf_clk new_AGEMA_reg_buffer_12875 ( .C (clk), .D (new_AGEMA_signal_33830), .Q (new_AGEMA_signal_33831) ) ;
    buf_clk new_AGEMA_reg_buffer_12879 ( .C (clk), .D (new_AGEMA_signal_33834), .Q (new_AGEMA_signal_33835) ) ;
    buf_clk new_AGEMA_reg_buffer_12883 ( .C (clk), .D (new_AGEMA_signal_33838), .Q (new_AGEMA_signal_33839) ) ;
    buf_clk new_AGEMA_reg_buffer_12887 ( .C (clk), .D (new_AGEMA_signal_33842), .Q (new_AGEMA_signal_33843) ) ;
    buf_clk new_AGEMA_reg_buffer_12891 ( .C (clk), .D (new_AGEMA_signal_33846), .Q (new_AGEMA_signal_33847) ) ;
    buf_clk new_AGEMA_reg_buffer_12895 ( .C (clk), .D (new_AGEMA_signal_33850), .Q (new_AGEMA_signal_33851) ) ;
    buf_clk new_AGEMA_reg_buffer_12899 ( .C (clk), .D (new_AGEMA_signal_33854), .Q (new_AGEMA_signal_33855) ) ;
    buf_clk new_AGEMA_reg_buffer_12903 ( .C (clk), .D (new_AGEMA_signal_33858), .Q (new_AGEMA_signal_33859) ) ;
    buf_clk new_AGEMA_reg_buffer_12907 ( .C (clk), .D (new_AGEMA_signal_33862), .Q (new_AGEMA_signal_33863) ) ;
    buf_clk new_AGEMA_reg_buffer_12911 ( .C (clk), .D (new_AGEMA_signal_33866), .Q (new_AGEMA_signal_33867) ) ;
    buf_clk new_AGEMA_reg_buffer_12915 ( .C (clk), .D (new_AGEMA_signal_33870), .Q (new_AGEMA_signal_33871) ) ;
    buf_clk new_AGEMA_reg_buffer_12919 ( .C (clk), .D (new_AGEMA_signal_33874), .Q (new_AGEMA_signal_33875) ) ;
    buf_clk new_AGEMA_reg_buffer_12923 ( .C (clk), .D (new_AGEMA_signal_33878), .Q (new_AGEMA_signal_33879) ) ;
    buf_clk new_AGEMA_reg_buffer_12927 ( .C (clk), .D (new_AGEMA_signal_33882), .Q (new_AGEMA_signal_33883) ) ;
    buf_clk new_AGEMA_reg_buffer_12931 ( .C (clk), .D (new_AGEMA_signal_33886), .Q (new_AGEMA_signal_33887) ) ;
    buf_clk new_AGEMA_reg_buffer_12935 ( .C (clk), .D (new_AGEMA_signal_33890), .Q (new_AGEMA_signal_33891) ) ;
    buf_clk new_AGEMA_reg_buffer_12939 ( .C (clk), .D (new_AGEMA_signal_33894), .Q (new_AGEMA_signal_33895) ) ;
    buf_clk new_AGEMA_reg_buffer_12943 ( .C (clk), .D (new_AGEMA_signal_33898), .Q (new_AGEMA_signal_33899) ) ;
    buf_clk new_AGEMA_reg_buffer_12947 ( .C (clk), .D (new_AGEMA_signal_33902), .Q (new_AGEMA_signal_33903) ) ;
    buf_clk new_AGEMA_reg_buffer_12951 ( .C (clk), .D (new_AGEMA_signal_33906), .Q (new_AGEMA_signal_33907) ) ;
    buf_clk new_AGEMA_reg_buffer_12955 ( .C (clk), .D (new_AGEMA_signal_33910), .Q (new_AGEMA_signal_33911) ) ;
    buf_clk new_AGEMA_reg_buffer_12959 ( .C (clk), .D (new_AGEMA_signal_33914), .Q (new_AGEMA_signal_33915) ) ;
    buf_clk new_AGEMA_reg_buffer_12963 ( .C (clk), .D (new_AGEMA_signal_33918), .Q (new_AGEMA_signal_33919) ) ;
    buf_clk new_AGEMA_reg_buffer_12967 ( .C (clk), .D (new_AGEMA_signal_33922), .Q (new_AGEMA_signal_33923) ) ;
    buf_clk new_AGEMA_reg_buffer_12971 ( .C (clk), .D (new_AGEMA_signal_33926), .Q (new_AGEMA_signal_33927) ) ;
    buf_clk new_AGEMA_reg_buffer_12975 ( .C (clk), .D (new_AGEMA_signal_33930), .Q (new_AGEMA_signal_33931) ) ;
    buf_clk new_AGEMA_reg_buffer_12979 ( .C (clk), .D (new_AGEMA_signal_33934), .Q (new_AGEMA_signal_33935) ) ;
    buf_clk new_AGEMA_reg_buffer_12983 ( .C (clk), .D (new_AGEMA_signal_33938), .Q (new_AGEMA_signal_33939) ) ;
    buf_clk new_AGEMA_reg_buffer_12987 ( .C (clk), .D (new_AGEMA_signal_33942), .Q (new_AGEMA_signal_33943) ) ;
    buf_clk new_AGEMA_reg_buffer_12991 ( .C (clk), .D (new_AGEMA_signal_33946), .Q (new_AGEMA_signal_33947) ) ;
    buf_clk new_AGEMA_reg_buffer_12995 ( .C (clk), .D (new_AGEMA_signal_33950), .Q (new_AGEMA_signal_33951) ) ;
    buf_clk new_AGEMA_reg_buffer_12999 ( .C (clk), .D (new_AGEMA_signal_33954), .Q (new_AGEMA_signal_33955) ) ;
    buf_clk new_AGEMA_reg_buffer_13003 ( .C (clk), .D (new_AGEMA_signal_33958), .Q (new_AGEMA_signal_33959) ) ;
    buf_clk new_AGEMA_reg_buffer_13007 ( .C (clk), .D (new_AGEMA_signal_33962), .Q (new_AGEMA_signal_33963) ) ;
    buf_clk new_AGEMA_reg_buffer_13011 ( .C (clk), .D (new_AGEMA_signal_33966), .Q (new_AGEMA_signal_33967) ) ;
    buf_clk new_AGEMA_reg_buffer_13015 ( .C (clk), .D (new_AGEMA_signal_33970), .Q (new_AGEMA_signal_33971) ) ;
    buf_clk new_AGEMA_reg_buffer_13019 ( .C (clk), .D (new_AGEMA_signal_33974), .Q (new_AGEMA_signal_33975) ) ;
    buf_clk new_AGEMA_reg_buffer_13023 ( .C (clk), .D (new_AGEMA_signal_33978), .Q (new_AGEMA_signal_33979) ) ;
    buf_clk new_AGEMA_reg_buffer_13027 ( .C (clk), .D (new_AGEMA_signal_33982), .Q (new_AGEMA_signal_33983) ) ;
    buf_clk new_AGEMA_reg_buffer_13031 ( .C (clk), .D (new_AGEMA_signal_33986), .Q (new_AGEMA_signal_33987) ) ;
    buf_clk new_AGEMA_reg_buffer_13035 ( .C (clk), .D (new_AGEMA_signal_33990), .Q (new_AGEMA_signal_33991) ) ;
    buf_clk new_AGEMA_reg_buffer_13039 ( .C (clk), .D (new_AGEMA_signal_33994), .Q (new_AGEMA_signal_33995) ) ;
    buf_clk new_AGEMA_reg_buffer_13043 ( .C (clk), .D (new_AGEMA_signal_33998), .Q (new_AGEMA_signal_33999) ) ;
    buf_clk new_AGEMA_reg_buffer_13047 ( .C (clk), .D (new_AGEMA_signal_34002), .Q (new_AGEMA_signal_34003) ) ;
    buf_clk new_AGEMA_reg_buffer_13051 ( .C (clk), .D (new_AGEMA_signal_34006), .Q (new_AGEMA_signal_34007) ) ;
    buf_clk new_AGEMA_reg_buffer_13055 ( .C (clk), .D (new_AGEMA_signal_34010), .Q (new_AGEMA_signal_34011) ) ;
    buf_clk new_AGEMA_reg_buffer_13059 ( .C (clk), .D (new_AGEMA_signal_34014), .Q (new_AGEMA_signal_34015) ) ;
    buf_clk new_AGEMA_reg_buffer_13063 ( .C (clk), .D (new_AGEMA_signal_34018), .Q (new_AGEMA_signal_34019) ) ;
    buf_clk new_AGEMA_reg_buffer_13067 ( .C (clk), .D (new_AGEMA_signal_34022), .Q (new_AGEMA_signal_34023) ) ;
    buf_clk new_AGEMA_reg_buffer_13071 ( .C (clk), .D (new_AGEMA_signal_34026), .Q (new_AGEMA_signal_34027) ) ;
    buf_clk new_AGEMA_reg_buffer_13075 ( .C (clk), .D (new_AGEMA_signal_34030), .Q (new_AGEMA_signal_34031) ) ;
    buf_clk new_AGEMA_reg_buffer_13079 ( .C (clk), .D (new_AGEMA_signal_34034), .Q (new_AGEMA_signal_34035) ) ;
    buf_clk new_AGEMA_reg_buffer_13083 ( .C (clk), .D (new_AGEMA_signal_34038), .Q (new_AGEMA_signal_34039) ) ;
    buf_clk new_AGEMA_reg_buffer_13087 ( .C (clk), .D (new_AGEMA_signal_34042), .Q (new_AGEMA_signal_34043) ) ;
    buf_clk new_AGEMA_reg_buffer_13091 ( .C (clk), .D (new_AGEMA_signal_34046), .Q (new_AGEMA_signal_34047) ) ;
    buf_clk new_AGEMA_reg_buffer_13095 ( .C (clk), .D (new_AGEMA_signal_34050), .Q (new_AGEMA_signal_34051) ) ;
    buf_clk new_AGEMA_reg_buffer_13099 ( .C (clk), .D (new_AGEMA_signal_34054), .Q (new_AGEMA_signal_34055) ) ;
    buf_clk new_AGEMA_reg_buffer_13103 ( .C (clk), .D (new_AGEMA_signal_34058), .Q (new_AGEMA_signal_34059) ) ;
    buf_clk new_AGEMA_reg_buffer_13107 ( .C (clk), .D (new_AGEMA_signal_34062), .Q (new_AGEMA_signal_34063) ) ;
    buf_clk new_AGEMA_reg_buffer_13111 ( .C (clk), .D (new_AGEMA_signal_34066), .Q (new_AGEMA_signal_34067) ) ;
    buf_clk new_AGEMA_reg_buffer_13115 ( .C (clk), .D (new_AGEMA_signal_34070), .Q (new_AGEMA_signal_34071) ) ;
    buf_clk new_AGEMA_reg_buffer_13119 ( .C (clk), .D (new_AGEMA_signal_34074), .Q (new_AGEMA_signal_34075) ) ;
    buf_clk new_AGEMA_reg_buffer_13123 ( .C (clk), .D (new_AGEMA_signal_34078), .Q (new_AGEMA_signal_34079) ) ;
    buf_clk new_AGEMA_reg_buffer_13127 ( .C (clk), .D (new_AGEMA_signal_34082), .Q (new_AGEMA_signal_34083) ) ;
    buf_clk new_AGEMA_reg_buffer_13131 ( .C (clk), .D (new_AGEMA_signal_34086), .Q (new_AGEMA_signal_34087) ) ;
    buf_clk new_AGEMA_reg_buffer_13135 ( .C (clk), .D (new_AGEMA_signal_34090), .Q (new_AGEMA_signal_34091) ) ;
    buf_clk new_AGEMA_reg_buffer_13139 ( .C (clk), .D (new_AGEMA_signal_34094), .Q (new_AGEMA_signal_34095) ) ;
    buf_clk new_AGEMA_reg_buffer_13143 ( .C (clk), .D (new_AGEMA_signal_34098), .Q (new_AGEMA_signal_34099) ) ;
    buf_clk new_AGEMA_reg_buffer_13147 ( .C (clk), .D (new_AGEMA_signal_34102), .Q (new_AGEMA_signal_34103) ) ;
    buf_clk new_AGEMA_reg_buffer_13151 ( .C (clk), .D (new_AGEMA_signal_34106), .Q (new_AGEMA_signal_34107) ) ;
    buf_clk new_AGEMA_reg_buffer_13155 ( .C (clk), .D (new_AGEMA_signal_34110), .Q (new_AGEMA_signal_34111) ) ;
    buf_clk new_AGEMA_reg_buffer_13159 ( .C (clk), .D (new_AGEMA_signal_34114), .Q (new_AGEMA_signal_34115) ) ;
    buf_clk new_AGEMA_reg_buffer_13163 ( .C (clk), .D (new_AGEMA_signal_34118), .Q (new_AGEMA_signal_34119) ) ;
    buf_clk new_AGEMA_reg_buffer_13167 ( .C (clk), .D (new_AGEMA_signal_34122), .Q (new_AGEMA_signal_34123) ) ;
    buf_clk new_AGEMA_reg_buffer_13171 ( .C (clk), .D (new_AGEMA_signal_34126), .Q (new_AGEMA_signal_34127) ) ;
    buf_clk new_AGEMA_reg_buffer_13175 ( .C (clk), .D (new_AGEMA_signal_34130), .Q (new_AGEMA_signal_34131) ) ;
    buf_clk new_AGEMA_reg_buffer_13179 ( .C (clk), .D (new_AGEMA_signal_34134), .Q (new_AGEMA_signal_34135) ) ;
    buf_clk new_AGEMA_reg_buffer_13183 ( .C (clk), .D (new_AGEMA_signal_34138), .Q (new_AGEMA_signal_34139) ) ;
    buf_clk new_AGEMA_reg_buffer_13187 ( .C (clk), .D (new_AGEMA_signal_34142), .Q (new_AGEMA_signal_34143) ) ;
    buf_clk new_AGEMA_reg_buffer_13191 ( .C (clk), .D (new_AGEMA_signal_34146), .Q (new_AGEMA_signal_34147) ) ;
    buf_clk new_AGEMA_reg_buffer_13195 ( .C (clk), .D (new_AGEMA_signal_34150), .Q (new_AGEMA_signal_34151) ) ;
    buf_clk new_AGEMA_reg_buffer_13199 ( .C (clk), .D (new_AGEMA_signal_34154), .Q (new_AGEMA_signal_34155) ) ;
    buf_clk new_AGEMA_reg_buffer_13203 ( .C (clk), .D (new_AGEMA_signal_34158), .Q (new_AGEMA_signal_34159) ) ;
    buf_clk new_AGEMA_reg_buffer_13207 ( .C (clk), .D (new_AGEMA_signal_34162), .Q (new_AGEMA_signal_34163) ) ;
    buf_clk new_AGEMA_reg_buffer_13211 ( .C (clk), .D (new_AGEMA_signal_34166), .Q (new_AGEMA_signal_34167) ) ;
    buf_clk new_AGEMA_reg_buffer_13215 ( .C (clk), .D (new_AGEMA_signal_34170), .Q (new_AGEMA_signal_34171) ) ;
    buf_clk new_AGEMA_reg_buffer_13219 ( .C (clk), .D (new_AGEMA_signal_34174), .Q (new_AGEMA_signal_34175) ) ;
    buf_clk new_AGEMA_reg_buffer_13223 ( .C (clk), .D (new_AGEMA_signal_34178), .Q (new_AGEMA_signal_34179) ) ;
    buf_clk new_AGEMA_reg_buffer_13227 ( .C (clk), .D (new_AGEMA_signal_34182), .Q (new_AGEMA_signal_34183) ) ;
    buf_clk new_AGEMA_reg_buffer_13231 ( .C (clk), .D (new_AGEMA_signal_34186), .Q (new_AGEMA_signal_34187) ) ;
    buf_clk new_AGEMA_reg_buffer_13235 ( .C (clk), .D (new_AGEMA_signal_34190), .Q (new_AGEMA_signal_34191) ) ;
    buf_clk new_AGEMA_reg_buffer_13239 ( .C (clk), .D (new_AGEMA_signal_34194), .Q (new_AGEMA_signal_34195) ) ;
    buf_clk new_AGEMA_reg_buffer_13243 ( .C (clk), .D (new_AGEMA_signal_34198), .Q (new_AGEMA_signal_34199) ) ;
    buf_clk new_AGEMA_reg_buffer_13247 ( .C (clk), .D (new_AGEMA_signal_34202), .Q (new_AGEMA_signal_34203) ) ;
    buf_clk new_AGEMA_reg_buffer_13251 ( .C (clk), .D (new_AGEMA_signal_34206), .Q (new_AGEMA_signal_34207) ) ;
    buf_clk new_AGEMA_reg_buffer_13255 ( .C (clk), .D (new_AGEMA_signal_34210), .Q (new_AGEMA_signal_34211) ) ;
    buf_clk new_AGEMA_reg_buffer_13259 ( .C (clk), .D (new_AGEMA_signal_34214), .Q (new_AGEMA_signal_34215) ) ;
    buf_clk new_AGEMA_reg_buffer_13263 ( .C (clk), .D (new_AGEMA_signal_34218), .Q (new_AGEMA_signal_34219) ) ;
    buf_clk new_AGEMA_reg_buffer_13267 ( .C (clk), .D (new_AGEMA_signal_34222), .Q (new_AGEMA_signal_34223) ) ;
    buf_clk new_AGEMA_reg_buffer_13271 ( .C (clk), .D (new_AGEMA_signal_34226), .Q (new_AGEMA_signal_34227) ) ;
    buf_clk new_AGEMA_reg_buffer_13275 ( .C (clk), .D (new_AGEMA_signal_34230), .Q (new_AGEMA_signal_34231) ) ;
    buf_clk new_AGEMA_reg_buffer_13279 ( .C (clk), .D (new_AGEMA_signal_34234), .Q (new_AGEMA_signal_34235) ) ;
    buf_clk new_AGEMA_reg_buffer_13283 ( .C (clk), .D (new_AGEMA_signal_34238), .Q (new_AGEMA_signal_34239) ) ;
    buf_clk new_AGEMA_reg_buffer_13287 ( .C (clk), .D (new_AGEMA_signal_34242), .Q (new_AGEMA_signal_34243) ) ;
    buf_clk new_AGEMA_reg_buffer_13291 ( .C (clk), .D (new_AGEMA_signal_34246), .Q (new_AGEMA_signal_34247) ) ;
    buf_clk new_AGEMA_reg_buffer_13295 ( .C (clk), .D (new_AGEMA_signal_34250), .Q (new_AGEMA_signal_34251) ) ;
    buf_clk new_AGEMA_reg_buffer_13299 ( .C (clk), .D (new_AGEMA_signal_34254), .Q (new_AGEMA_signal_34255) ) ;
    buf_clk new_AGEMA_reg_buffer_13303 ( .C (clk), .D (new_AGEMA_signal_34258), .Q (new_AGEMA_signal_34259) ) ;
    buf_clk new_AGEMA_reg_buffer_13307 ( .C (clk), .D (new_AGEMA_signal_34262), .Q (new_AGEMA_signal_34263) ) ;
    buf_clk new_AGEMA_reg_buffer_13311 ( .C (clk), .D (new_AGEMA_signal_34266), .Q (new_AGEMA_signal_34267) ) ;
    buf_clk new_AGEMA_reg_buffer_13315 ( .C (clk), .D (new_AGEMA_signal_34270), .Q (new_AGEMA_signal_34271) ) ;
    buf_clk new_AGEMA_reg_buffer_13319 ( .C (clk), .D (new_AGEMA_signal_34274), .Q (new_AGEMA_signal_34275) ) ;
    buf_clk new_AGEMA_reg_buffer_13323 ( .C (clk), .D (new_AGEMA_signal_34278), .Q (new_AGEMA_signal_34279) ) ;
    buf_clk new_AGEMA_reg_buffer_13327 ( .C (clk), .D (new_AGEMA_signal_34282), .Q (new_AGEMA_signal_34283) ) ;
    buf_clk new_AGEMA_reg_buffer_13331 ( .C (clk), .D (new_AGEMA_signal_34286), .Q (new_AGEMA_signal_34287) ) ;
    buf_clk new_AGEMA_reg_buffer_13335 ( .C (clk), .D (new_AGEMA_signal_34290), .Q (new_AGEMA_signal_34291) ) ;
    buf_clk new_AGEMA_reg_buffer_13339 ( .C (clk), .D (new_AGEMA_signal_34294), .Q (new_AGEMA_signal_34295) ) ;
    buf_clk new_AGEMA_reg_buffer_13343 ( .C (clk), .D (new_AGEMA_signal_34298), .Q (new_AGEMA_signal_34299) ) ;
    buf_clk new_AGEMA_reg_buffer_13347 ( .C (clk), .D (new_AGEMA_signal_34302), .Q (new_AGEMA_signal_34303) ) ;
    buf_clk new_AGEMA_reg_buffer_13351 ( .C (clk), .D (new_AGEMA_signal_34306), .Q (new_AGEMA_signal_34307) ) ;
    buf_clk new_AGEMA_reg_buffer_13355 ( .C (clk), .D (new_AGEMA_signal_34310), .Q (new_AGEMA_signal_34311) ) ;
    buf_clk new_AGEMA_reg_buffer_13359 ( .C (clk), .D (new_AGEMA_signal_34314), .Q (new_AGEMA_signal_34315) ) ;
    buf_clk new_AGEMA_reg_buffer_13363 ( .C (clk), .D (new_AGEMA_signal_34318), .Q (new_AGEMA_signal_34319) ) ;
    buf_clk new_AGEMA_reg_buffer_13367 ( .C (clk), .D (new_AGEMA_signal_34322), .Q (new_AGEMA_signal_34323) ) ;
    buf_clk new_AGEMA_reg_buffer_13371 ( .C (clk), .D (new_AGEMA_signal_34326), .Q (new_AGEMA_signal_34327) ) ;
    buf_clk new_AGEMA_reg_buffer_13375 ( .C (clk), .D (new_AGEMA_signal_34330), .Q (new_AGEMA_signal_34331) ) ;
    buf_clk new_AGEMA_reg_buffer_13379 ( .C (clk), .D (new_AGEMA_signal_34334), .Q (new_AGEMA_signal_34335) ) ;
    buf_clk new_AGEMA_reg_buffer_13383 ( .C (clk), .D (new_AGEMA_signal_34338), .Q (new_AGEMA_signal_34339) ) ;
    buf_clk new_AGEMA_reg_buffer_13387 ( .C (clk), .D (new_AGEMA_signal_34342), .Q (new_AGEMA_signal_34343) ) ;
    buf_clk new_AGEMA_reg_buffer_13391 ( .C (clk), .D (new_AGEMA_signal_34346), .Q (new_AGEMA_signal_34347) ) ;
    buf_clk new_AGEMA_reg_buffer_13395 ( .C (clk), .D (new_AGEMA_signal_34350), .Q (new_AGEMA_signal_34351) ) ;
    buf_clk new_AGEMA_reg_buffer_13399 ( .C (clk), .D (new_AGEMA_signal_34354), .Q (new_AGEMA_signal_34355) ) ;
    buf_clk new_AGEMA_reg_buffer_13403 ( .C (clk), .D (new_AGEMA_signal_34358), .Q (new_AGEMA_signal_34359) ) ;
    buf_clk new_AGEMA_reg_buffer_13407 ( .C (clk), .D (new_AGEMA_signal_34362), .Q (new_AGEMA_signal_34363) ) ;
    buf_clk new_AGEMA_reg_buffer_13411 ( .C (clk), .D (new_AGEMA_signal_34366), .Q (new_AGEMA_signal_34367) ) ;
    buf_clk new_AGEMA_reg_buffer_13415 ( .C (clk), .D (new_AGEMA_signal_34370), .Q (new_AGEMA_signal_34371) ) ;
    buf_clk new_AGEMA_reg_buffer_13419 ( .C (clk), .D (new_AGEMA_signal_34374), .Q (new_AGEMA_signal_34375) ) ;
    buf_clk new_AGEMA_reg_buffer_13423 ( .C (clk), .D (new_AGEMA_signal_34378), .Q (new_AGEMA_signal_34379) ) ;
    buf_clk new_AGEMA_reg_buffer_13427 ( .C (clk), .D (new_AGEMA_signal_34382), .Q (new_AGEMA_signal_34383) ) ;
    buf_clk new_AGEMA_reg_buffer_13431 ( .C (clk), .D (new_AGEMA_signal_34386), .Q (new_AGEMA_signal_34387) ) ;
    buf_clk new_AGEMA_reg_buffer_13435 ( .C (clk), .D (new_AGEMA_signal_34390), .Q (new_AGEMA_signal_34391) ) ;
    buf_clk new_AGEMA_reg_buffer_13439 ( .C (clk), .D (new_AGEMA_signal_34394), .Q (new_AGEMA_signal_34395) ) ;
    buf_clk new_AGEMA_reg_buffer_13443 ( .C (clk), .D (new_AGEMA_signal_34398), .Q (new_AGEMA_signal_34399) ) ;
    buf_clk new_AGEMA_reg_buffer_13447 ( .C (clk), .D (new_AGEMA_signal_34402), .Q (new_AGEMA_signal_34403) ) ;
    buf_clk new_AGEMA_reg_buffer_13451 ( .C (clk), .D (new_AGEMA_signal_34406), .Q (new_AGEMA_signal_34407) ) ;
    buf_clk new_AGEMA_reg_buffer_13455 ( .C (clk), .D (new_AGEMA_signal_34410), .Q (new_AGEMA_signal_34411) ) ;
    buf_clk new_AGEMA_reg_buffer_13459 ( .C (clk), .D (new_AGEMA_signal_34414), .Q (new_AGEMA_signal_34415) ) ;
    buf_clk new_AGEMA_reg_buffer_13463 ( .C (clk), .D (new_AGEMA_signal_34418), .Q (new_AGEMA_signal_34419) ) ;
    buf_clk new_AGEMA_reg_buffer_13467 ( .C (clk), .D (new_AGEMA_signal_34422), .Q (new_AGEMA_signal_34423) ) ;
    buf_clk new_AGEMA_reg_buffer_13471 ( .C (clk), .D (new_AGEMA_signal_34426), .Q (new_AGEMA_signal_34427) ) ;
    buf_clk new_AGEMA_reg_buffer_13475 ( .C (clk), .D (new_AGEMA_signal_34430), .Q (new_AGEMA_signal_34431) ) ;
    buf_clk new_AGEMA_reg_buffer_13479 ( .C (clk), .D (new_AGEMA_signal_34434), .Q (new_AGEMA_signal_34435) ) ;
    buf_clk new_AGEMA_reg_buffer_13483 ( .C (clk), .D (new_AGEMA_signal_34438), .Q (new_AGEMA_signal_34439) ) ;
    buf_clk new_AGEMA_reg_buffer_13487 ( .C (clk), .D (new_AGEMA_signal_34442), .Q (new_AGEMA_signal_34443) ) ;
    buf_clk new_AGEMA_reg_buffer_13491 ( .C (clk), .D (new_AGEMA_signal_34446), .Q (new_AGEMA_signal_34447) ) ;
    buf_clk new_AGEMA_reg_buffer_13495 ( .C (clk), .D (new_AGEMA_signal_34450), .Q (new_AGEMA_signal_34451) ) ;
    buf_clk new_AGEMA_reg_buffer_13499 ( .C (clk), .D (new_AGEMA_signal_34454), .Q (new_AGEMA_signal_34455) ) ;
    buf_clk new_AGEMA_reg_buffer_13503 ( .C (clk), .D (new_AGEMA_signal_34458), .Q (new_AGEMA_signal_34459) ) ;
    buf_clk new_AGEMA_reg_buffer_13507 ( .C (clk), .D (new_AGEMA_signal_34462), .Q (new_AGEMA_signal_34463) ) ;
    buf_clk new_AGEMA_reg_buffer_13511 ( .C (clk), .D (new_AGEMA_signal_34466), .Q (new_AGEMA_signal_34467) ) ;
    buf_clk new_AGEMA_reg_buffer_13515 ( .C (clk), .D (new_AGEMA_signal_34470), .Q (new_AGEMA_signal_34471) ) ;
    buf_clk new_AGEMA_reg_buffer_13519 ( .C (clk), .D (new_AGEMA_signal_34474), .Q (new_AGEMA_signal_34475) ) ;
    buf_clk new_AGEMA_reg_buffer_13523 ( .C (clk), .D (new_AGEMA_signal_34478), .Q (new_AGEMA_signal_34479) ) ;
    buf_clk new_AGEMA_reg_buffer_13527 ( .C (clk), .D (new_AGEMA_signal_34482), .Q (new_AGEMA_signal_34483) ) ;
    buf_clk new_AGEMA_reg_buffer_13531 ( .C (clk), .D (new_AGEMA_signal_34486), .Q (new_AGEMA_signal_34487) ) ;
    buf_clk new_AGEMA_reg_buffer_13535 ( .C (clk), .D (new_AGEMA_signal_34490), .Q (new_AGEMA_signal_34491) ) ;
    buf_clk new_AGEMA_reg_buffer_13539 ( .C (clk), .D (new_AGEMA_signal_34494), .Q (new_AGEMA_signal_34495) ) ;
    buf_clk new_AGEMA_reg_buffer_13543 ( .C (clk), .D (new_AGEMA_signal_34498), .Q (new_AGEMA_signal_34499) ) ;
    buf_clk new_AGEMA_reg_buffer_13547 ( .C (clk), .D (new_AGEMA_signal_34502), .Q (new_AGEMA_signal_34503) ) ;
    buf_clk new_AGEMA_reg_buffer_13551 ( .C (clk), .D (new_AGEMA_signal_34506), .Q (new_AGEMA_signal_34507) ) ;
    buf_clk new_AGEMA_reg_buffer_13555 ( .C (clk), .D (new_AGEMA_signal_34510), .Q (new_AGEMA_signal_34511) ) ;
    buf_clk new_AGEMA_reg_buffer_13559 ( .C (clk), .D (new_AGEMA_signal_34514), .Q (new_AGEMA_signal_34515) ) ;
    buf_clk new_AGEMA_reg_buffer_13563 ( .C (clk), .D (new_AGEMA_signal_34518), .Q (new_AGEMA_signal_34519) ) ;
    buf_clk new_AGEMA_reg_buffer_13567 ( .C (clk), .D (new_AGEMA_signal_34522), .Q (new_AGEMA_signal_34523) ) ;
    buf_clk new_AGEMA_reg_buffer_13571 ( .C (clk), .D (new_AGEMA_signal_34526), .Q (new_AGEMA_signal_34527) ) ;
    buf_clk new_AGEMA_reg_buffer_13575 ( .C (clk), .D (new_AGEMA_signal_34530), .Q (new_AGEMA_signal_34531) ) ;
    buf_clk new_AGEMA_reg_buffer_13579 ( .C (clk), .D (new_AGEMA_signal_34534), .Q (new_AGEMA_signal_34535) ) ;
    buf_clk new_AGEMA_reg_buffer_13583 ( .C (clk), .D (new_AGEMA_signal_34538), .Q (new_AGEMA_signal_34539) ) ;
    buf_clk new_AGEMA_reg_buffer_13587 ( .C (clk), .D (new_AGEMA_signal_34542), .Q (new_AGEMA_signal_34543) ) ;
    buf_clk new_AGEMA_reg_buffer_13591 ( .C (clk), .D (new_AGEMA_signal_34546), .Q (new_AGEMA_signal_34547) ) ;
    buf_clk new_AGEMA_reg_buffer_13595 ( .C (clk), .D (new_AGEMA_signal_34550), .Q (new_AGEMA_signal_34551) ) ;
    buf_clk new_AGEMA_reg_buffer_13599 ( .C (clk), .D (new_AGEMA_signal_34554), .Q (new_AGEMA_signal_34555) ) ;
    buf_clk new_AGEMA_reg_buffer_13603 ( .C (clk), .D (new_AGEMA_signal_34558), .Q (new_AGEMA_signal_34559) ) ;
    buf_clk new_AGEMA_reg_buffer_13607 ( .C (clk), .D (new_AGEMA_signal_34562), .Q (new_AGEMA_signal_34563) ) ;
    buf_clk new_AGEMA_reg_buffer_13611 ( .C (clk), .D (new_AGEMA_signal_34566), .Q (new_AGEMA_signal_34567) ) ;
    buf_clk new_AGEMA_reg_buffer_13615 ( .C (clk), .D (new_AGEMA_signal_34570), .Q (new_AGEMA_signal_34571) ) ;
    buf_clk new_AGEMA_reg_buffer_13619 ( .C (clk), .D (new_AGEMA_signal_34574), .Q (new_AGEMA_signal_34575) ) ;
    buf_clk new_AGEMA_reg_buffer_13623 ( .C (clk), .D (new_AGEMA_signal_34578), .Q (new_AGEMA_signal_34579) ) ;
    buf_clk new_AGEMA_reg_buffer_13627 ( .C (clk), .D (new_AGEMA_signal_34582), .Q (new_AGEMA_signal_34583) ) ;
    buf_clk new_AGEMA_reg_buffer_13631 ( .C (clk), .D (new_AGEMA_signal_34586), .Q (new_AGEMA_signal_34587) ) ;
    buf_clk new_AGEMA_reg_buffer_13635 ( .C (clk), .D (new_AGEMA_signal_34590), .Q (new_AGEMA_signal_34591) ) ;
    buf_clk new_AGEMA_reg_buffer_13639 ( .C (clk), .D (new_AGEMA_signal_34594), .Q (new_AGEMA_signal_34595) ) ;
    buf_clk new_AGEMA_reg_buffer_13643 ( .C (clk), .D (new_AGEMA_signal_34598), .Q (new_AGEMA_signal_34599) ) ;
    buf_clk new_AGEMA_reg_buffer_13647 ( .C (clk), .D (new_AGEMA_signal_34602), .Q (new_AGEMA_signal_34603) ) ;
    buf_clk new_AGEMA_reg_buffer_13651 ( .C (clk), .D (new_AGEMA_signal_34606), .Q (new_AGEMA_signal_34607) ) ;
    buf_clk new_AGEMA_reg_buffer_13655 ( .C (clk), .D (new_AGEMA_signal_34610), .Q (new_AGEMA_signal_34611) ) ;
    buf_clk new_AGEMA_reg_buffer_13659 ( .C (clk), .D (new_AGEMA_signal_34614), .Q (new_AGEMA_signal_34615) ) ;
    buf_clk new_AGEMA_reg_buffer_13663 ( .C (clk), .D (new_AGEMA_signal_34618), .Q (new_AGEMA_signal_34619) ) ;
    buf_clk new_AGEMA_reg_buffer_13667 ( .C (clk), .D (new_AGEMA_signal_34622), .Q (new_AGEMA_signal_34623) ) ;
    buf_clk new_AGEMA_reg_buffer_13671 ( .C (clk), .D (new_AGEMA_signal_34626), .Q (new_AGEMA_signal_34627) ) ;
    buf_clk new_AGEMA_reg_buffer_13675 ( .C (clk), .D (new_AGEMA_signal_34630), .Q (new_AGEMA_signal_34631) ) ;
    buf_clk new_AGEMA_reg_buffer_13679 ( .C (clk), .D (new_AGEMA_signal_34634), .Q (new_AGEMA_signal_34635) ) ;
    buf_clk new_AGEMA_reg_buffer_13683 ( .C (clk), .D (new_AGEMA_signal_34638), .Q (new_AGEMA_signal_34639) ) ;
    buf_clk new_AGEMA_reg_buffer_13687 ( .C (clk), .D (new_AGEMA_signal_34642), .Q (new_AGEMA_signal_34643) ) ;
    buf_clk new_AGEMA_reg_buffer_13691 ( .C (clk), .D (new_AGEMA_signal_34646), .Q (new_AGEMA_signal_34647) ) ;
    buf_clk new_AGEMA_reg_buffer_13695 ( .C (clk), .D (new_AGEMA_signal_34650), .Q (new_AGEMA_signal_34651) ) ;
    buf_clk new_AGEMA_reg_buffer_13699 ( .C (clk), .D (new_AGEMA_signal_34654), .Q (new_AGEMA_signal_34655) ) ;
    buf_clk new_AGEMA_reg_buffer_13703 ( .C (clk), .D (new_AGEMA_signal_34658), .Q (new_AGEMA_signal_34659) ) ;
    buf_clk new_AGEMA_reg_buffer_13707 ( .C (clk), .D (new_AGEMA_signal_34662), .Q (new_AGEMA_signal_34663) ) ;
    buf_clk new_AGEMA_reg_buffer_13711 ( .C (clk), .D (new_AGEMA_signal_34666), .Q (new_AGEMA_signal_34667) ) ;
    buf_clk new_AGEMA_reg_buffer_13715 ( .C (clk), .D (new_AGEMA_signal_34670), .Q (new_AGEMA_signal_34671) ) ;
    buf_clk new_AGEMA_reg_buffer_13719 ( .C (clk), .D (new_AGEMA_signal_34674), .Q (new_AGEMA_signal_34675) ) ;
    buf_clk new_AGEMA_reg_buffer_13723 ( .C (clk), .D (new_AGEMA_signal_34678), .Q (new_AGEMA_signal_34679) ) ;
    buf_clk new_AGEMA_reg_buffer_13727 ( .C (clk), .D (new_AGEMA_signal_34682), .Q (new_AGEMA_signal_34683) ) ;
    buf_clk new_AGEMA_reg_buffer_13731 ( .C (clk), .D (new_AGEMA_signal_34686), .Q (new_AGEMA_signal_34687) ) ;
    buf_clk new_AGEMA_reg_buffer_13735 ( .C (clk), .D (new_AGEMA_signal_34690), .Q (new_AGEMA_signal_34691) ) ;
    buf_clk new_AGEMA_reg_buffer_13739 ( .C (clk), .D (new_AGEMA_signal_34694), .Q (new_AGEMA_signal_34695) ) ;
    buf_clk new_AGEMA_reg_buffer_13743 ( .C (clk), .D (new_AGEMA_signal_34698), .Q (new_AGEMA_signal_34699) ) ;
    buf_clk new_AGEMA_reg_buffer_13747 ( .C (clk), .D (new_AGEMA_signal_34702), .Q (new_AGEMA_signal_34703) ) ;
    buf_clk new_AGEMA_reg_buffer_13751 ( .C (clk), .D (new_AGEMA_signal_34706), .Q (new_AGEMA_signal_34707) ) ;
    buf_clk new_AGEMA_reg_buffer_13755 ( .C (clk), .D (new_AGEMA_signal_34710), .Q (new_AGEMA_signal_34711) ) ;
    buf_clk new_AGEMA_reg_buffer_13759 ( .C (clk), .D (new_AGEMA_signal_34714), .Q (new_AGEMA_signal_34715) ) ;
    buf_clk new_AGEMA_reg_buffer_13763 ( .C (clk), .D (new_AGEMA_signal_34718), .Q (new_AGEMA_signal_34719) ) ;
    buf_clk new_AGEMA_reg_buffer_13767 ( .C (clk), .D (new_AGEMA_signal_34722), .Q (new_AGEMA_signal_34723) ) ;
    buf_clk new_AGEMA_reg_buffer_13771 ( .C (clk), .D (new_AGEMA_signal_34726), .Q (new_AGEMA_signal_34727) ) ;
    buf_clk new_AGEMA_reg_buffer_13775 ( .C (clk), .D (new_AGEMA_signal_34730), .Q (new_AGEMA_signal_34731) ) ;
    buf_clk new_AGEMA_reg_buffer_13779 ( .C (clk), .D (new_AGEMA_signal_34734), .Q (new_AGEMA_signal_34735) ) ;
    buf_clk new_AGEMA_reg_buffer_13783 ( .C (clk), .D (new_AGEMA_signal_34738), .Q (new_AGEMA_signal_34739) ) ;
    buf_clk new_AGEMA_reg_buffer_13787 ( .C (clk), .D (new_AGEMA_signal_34742), .Q (new_AGEMA_signal_34743) ) ;
    buf_clk new_AGEMA_reg_buffer_13791 ( .C (clk), .D (new_AGEMA_signal_34746), .Q (new_AGEMA_signal_34747) ) ;
    buf_clk new_AGEMA_reg_buffer_13795 ( .C (clk), .D (new_AGEMA_signal_34750), .Q (new_AGEMA_signal_34751) ) ;
    buf_clk new_AGEMA_reg_buffer_13799 ( .C (clk), .D (new_AGEMA_signal_34754), .Q (new_AGEMA_signal_34755) ) ;
    buf_clk new_AGEMA_reg_buffer_13803 ( .C (clk), .D (new_AGEMA_signal_34758), .Q (new_AGEMA_signal_34759) ) ;
    buf_clk new_AGEMA_reg_buffer_13807 ( .C (clk), .D (new_AGEMA_signal_34762), .Q (new_AGEMA_signal_34763) ) ;
    buf_clk new_AGEMA_reg_buffer_13811 ( .C (clk), .D (new_AGEMA_signal_34766), .Q (new_AGEMA_signal_34767) ) ;
    buf_clk new_AGEMA_reg_buffer_13815 ( .C (clk), .D (new_AGEMA_signal_34770), .Q (new_AGEMA_signal_34771) ) ;
    buf_clk new_AGEMA_reg_buffer_13819 ( .C (clk), .D (new_AGEMA_signal_34774), .Q (new_AGEMA_signal_34775) ) ;
    buf_clk new_AGEMA_reg_buffer_13823 ( .C (clk), .D (new_AGEMA_signal_34778), .Q (new_AGEMA_signal_34779) ) ;
    buf_clk new_AGEMA_reg_buffer_13827 ( .C (clk), .D (new_AGEMA_signal_34782), .Q (new_AGEMA_signal_34783) ) ;
    buf_clk new_AGEMA_reg_buffer_13831 ( .C (clk), .D (new_AGEMA_signal_34786), .Q (new_AGEMA_signal_34787) ) ;
    buf_clk new_AGEMA_reg_buffer_13835 ( .C (clk), .D (new_AGEMA_signal_34790), .Q (new_AGEMA_signal_34791) ) ;
    buf_clk new_AGEMA_reg_buffer_13839 ( .C (clk), .D (new_AGEMA_signal_34794), .Q (new_AGEMA_signal_34795) ) ;
    buf_clk new_AGEMA_reg_buffer_13843 ( .C (clk), .D (new_AGEMA_signal_34798), .Q (new_AGEMA_signal_34799) ) ;
    buf_clk new_AGEMA_reg_buffer_13847 ( .C (clk), .D (new_AGEMA_signal_34802), .Q (new_AGEMA_signal_34803) ) ;
    buf_clk new_AGEMA_reg_buffer_13851 ( .C (clk), .D (new_AGEMA_signal_34806), .Q (new_AGEMA_signal_34807) ) ;
    buf_clk new_AGEMA_reg_buffer_13855 ( .C (clk), .D (new_AGEMA_signal_34810), .Q (new_AGEMA_signal_34811) ) ;
    buf_clk new_AGEMA_reg_buffer_13859 ( .C (clk), .D (new_AGEMA_signal_34814), .Q (new_AGEMA_signal_34815) ) ;
    buf_clk new_AGEMA_reg_buffer_13863 ( .C (clk), .D (new_AGEMA_signal_34818), .Q (new_AGEMA_signal_34819) ) ;
    buf_clk new_AGEMA_reg_buffer_13867 ( .C (clk), .D (new_AGEMA_signal_34822), .Q (new_AGEMA_signal_34823) ) ;
    buf_clk new_AGEMA_reg_buffer_13871 ( .C (clk), .D (new_AGEMA_signal_34826), .Q (new_AGEMA_signal_34827) ) ;
    buf_clk new_AGEMA_reg_buffer_13875 ( .C (clk), .D (new_AGEMA_signal_34830), .Q (new_AGEMA_signal_34831) ) ;
    buf_clk new_AGEMA_reg_buffer_13879 ( .C (clk), .D (new_AGEMA_signal_34834), .Q (new_AGEMA_signal_34835) ) ;
    buf_clk new_AGEMA_reg_buffer_13883 ( .C (clk), .D (new_AGEMA_signal_34838), .Q (new_AGEMA_signal_34839) ) ;
    buf_clk new_AGEMA_reg_buffer_13887 ( .C (clk), .D (new_AGEMA_signal_34842), .Q (new_AGEMA_signal_34843) ) ;
    buf_clk new_AGEMA_reg_buffer_13891 ( .C (clk), .D (new_AGEMA_signal_34846), .Q (new_AGEMA_signal_34847) ) ;
    buf_clk new_AGEMA_reg_buffer_13895 ( .C (clk), .D (new_AGEMA_signal_34850), .Q (new_AGEMA_signal_34851) ) ;
    buf_clk new_AGEMA_reg_buffer_13899 ( .C (clk), .D (new_AGEMA_signal_34854), .Q (new_AGEMA_signal_34855) ) ;
    buf_clk new_AGEMA_reg_buffer_13903 ( .C (clk), .D (new_AGEMA_signal_34858), .Q (new_AGEMA_signal_34859) ) ;
    buf_clk new_AGEMA_reg_buffer_13907 ( .C (clk), .D (new_AGEMA_signal_34862), .Q (new_AGEMA_signal_34863) ) ;
    buf_clk new_AGEMA_reg_buffer_13911 ( .C (clk), .D (new_AGEMA_signal_34866), .Q (new_AGEMA_signal_34867) ) ;
    buf_clk new_AGEMA_reg_buffer_13915 ( .C (clk), .D (new_AGEMA_signal_34870), .Q (new_AGEMA_signal_34871) ) ;
    buf_clk new_AGEMA_reg_buffer_13919 ( .C (clk), .D (new_AGEMA_signal_34874), .Q (new_AGEMA_signal_34875) ) ;
    buf_clk new_AGEMA_reg_buffer_13923 ( .C (clk), .D (new_AGEMA_signal_34878), .Q (new_AGEMA_signal_34879) ) ;
    buf_clk new_AGEMA_reg_buffer_13927 ( .C (clk), .D (new_AGEMA_signal_34882), .Q (new_AGEMA_signal_34883) ) ;
    buf_clk new_AGEMA_reg_buffer_13931 ( .C (clk), .D (new_AGEMA_signal_34886), .Q (new_AGEMA_signal_34887) ) ;
    buf_clk new_AGEMA_reg_buffer_13935 ( .C (clk), .D (new_AGEMA_signal_34890), .Q (new_AGEMA_signal_34891) ) ;
    buf_clk new_AGEMA_reg_buffer_13939 ( .C (clk), .D (new_AGEMA_signal_34894), .Q (new_AGEMA_signal_34895) ) ;
    buf_clk new_AGEMA_reg_buffer_13943 ( .C (clk), .D (new_AGEMA_signal_34898), .Q (new_AGEMA_signal_34899) ) ;
    buf_clk new_AGEMA_reg_buffer_13947 ( .C (clk), .D (new_AGEMA_signal_34902), .Q (new_AGEMA_signal_34903) ) ;
    buf_clk new_AGEMA_reg_buffer_13951 ( .C (clk), .D (new_AGEMA_signal_34906), .Q (new_AGEMA_signal_34907) ) ;
    buf_clk new_AGEMA_reg_buffer_13955 ( .C (clk), .D (new_AGEMA_signal_34910), .Q (new_AGEMA_signal_34911) ) ;
    buf_clk new_AGEMA_reg_buffer_13959 ( .C (clk), .D (new_AGEMA_signal_34914), .Q (new_AGEMA_signal_34915) ) ;
    buf_clk new_AGEMA_reg_buffer_13963 ( .C (clk), .D (new_AGEMA_signal_34918), .Q (new_AGEMA_signal_34919) ) ;
    buf_clk new_AGEMA_reg_buffer_13967 ( .C (clk), .D (new_AGEMA_signal_34922), .Q (new_AGEMA_signal_34923) ) ;
    buf_clk new_AGEMA_reg_buffer_13971 ( .C (clk), .D (new_AGEMA_signal_34926), .Q (new_AGEMA_signal_34927) ) ;
    buf_clk new_AGEMA_reg_buffer_13975 ( .C (clk), .D (new_AGEMA_signal_34930), .Q (new_AGEMA_signal_34931) ) ;
    buf_clk new_AGEMA_reg_buffer_13979 ( .C (clk), .D (new_AGEMA_signal_34934), .Q (new_AGEMA_signal_34935) ) ;
    buf_clk new_AGEMA_reg_buffer_13983 ( .C (clk), .D (new_AGEMA_signal_34938), .Q (new_AGEMA_signal_34939) ) ;
    buf_clk new_AGEMA_reg_buffer_13987 ( .C (clk), .D (new_AGEMA_signal_34942), .Q (new_AGEMA_signal_34943) ) ;
    buf_clk new_AGEMA_reg_buffer_13991 ( .C (clk), .D (new_AGEMA_signal_34946), .Q (new_AGEMA_signal_34947) ) ;
    buf_clk new_AGEMA_reg_buffer_13995 ( .C (clk), .D (new_AGEMA_signal_34950), .Q (new_AGEMA_signal_34951) ) ;
    buf_clk new_AGEMA_reg_buffer_13999 ( .C (clk), .D (new_AGEMA_signal_34954), .Q (new_AGEMA_signal_34955) ) ;
    buf_clk new_AGEMA_reg_buffer_14003 ( .C (clk), .D (new_AGEMA_signal_34958), .Q (new_AGEMA_signal_34959) ) ;
    buf_clk new_AGEMA_reg_buffer_14007 ( .C (clk), .D (new_AGEMA_signal_34962), .Q (new_AGEMA_signal_34963) ) ;
    buf_clk new_AGEMA_reg_buffer_14011 ( .C (clk), .D (new_AGEMA_signal_34966), .Q (new_AGEMA_signal_34967) ) ;
    buf_clk new_AGEMA_reg_buffer_14015 ( .C (clk), .D (new_AGEMA_signal_34970), .Q (new_AGEMA_signal_34971) ) ;
    buf_clk new_AGEMA_reg_buffer_14019 ( .C (clk), .D (new_AGEMA_signal_34974), .Q (new_AGEMA_signal_34975) ) ;
    buf_clk new_AGEMA_reg_buffer_14023 ( .C (clk), .D (new_AGEMA_signal_34978), .Q (new_AGEMA_signal_34979) ) ;
    buf_clk new_AGEMA_reg_buffer_14027 ( .C (clk), .D (new_AGEMA_signal_34982), .Q (new_AGEMA_signal_34983) ) ;
    buf_clk new_AGEMA_reg_buffer_14031 ( .C (clk), .D (new_AGEMA_signal_34986), .Q (new_AGEMA_signal_34987) ) ;
    buf_clk new_AGEMA_reg_buffer_14035 ( .C (clk), .D (new_AGEMA_signal_34990), .Q (new_AGEMA_signal_34991) ) ;
    buf_clk new_AGEMA_reg_buffer_14039 ( .C (clk), .D (new_AGEMA_signal_34994), .Q (new_AGEMA_signal_34995) ) ;
    buf_clk new_AGEMA_reg_buffer_14043 ( .C (clk), .D (new_AGEMA_signal_34998), .Q (new_AGEMA_signal_34999) ) ;
    buf_clk new_AGEMA_reg_buffer_14047 ( .C (clk), .D (new_AGEMA_signal_35002), .Q (new_AGEMA_signal_35003) ) ;
    buf_clk new_AGEMA_reg_buffer_14051 ( .C (clk), .D (new_AGEMA_signal_35006), .Q (new_AGEMA_signal_35007) ) ;
    buf_clk new_AGEMA_reg_buffer_14055 ( .C (clk), .D (new_AGEMA_signal_35010), .Q (new_AGEMA_signal_35011) ) ;
    buf_clk new_AGEMA_reg_buffer_14059 ( .C (clk), .D (new_AGEMA_signal_35014), .Q (new_AGEMA_signal_35015) ) ;
    buf_clk new_AGEMA_reg_buffer_14063 ( .C (clk), .D (new_AGEMA_signal_35018), .Q (new_AGEMA_signal_35019) ) ;
    buf_clk new_AGEMA_reg_buffer_14067 ( .C (clk), .D (new_AGEMA_signal_35022), .Q (new_AGEMA_signal_35023) ) ;
    buf_clk new_AGEMA_reg_buffer_14071 ( .C (clk), .D (new_AGEMA_signal_35026), .Q (new_AGEMA_signal_35027) ) ;
    buf_clk new_AGEMA_reg_buffer_14075 ( .C (clk), .D (new_AGEMA_signal_35030), .Q (new_AGEMA_signal_35031) ) ;
    buf_clk new_AGEMA_reg_buffer_14079 ( .C (clk), .D (new_AGEMA_signal_35034), .Q (new_AGEMA_signal_35035) ) ;
    buf_clk new_AGEMA_reg_buffer_14083 ( .C (clk), .D (new_AGEMA_signal_35038), .Q (new_AGEMA_signal_35039) ) ;
    buf_clk new_AGEMA_reg_buffer_14087 ( .C (clk), .D (new_AGEMA_signal_35042), .Q (new_AGEMA_signal_35043) ) ;
    buf_clk new_AGEMA_reg_buffer_14091 ( .C (clk), .D (new_AGEMA_signal_35046), .Q (new_AGEMA_signal_35047) ) ;
    buf_clk new_AGEMA_reg_buffer_14095 ( .C (clk), .D (new_AGEMA_signal_35050), .Q (new_AGEMA_signal_35051) ) ;
    buf_clk new_AGEMA_reg_buffer_14099 ( .C (clk), .D (new_AGEMA_signal_35054), .Q (new_AGEMA_signal_35055) ) ;
    buf_clk new_AGEMA_reg_buffer_14103 ( .C (clk), .D (new_AGEMA_signal_35058), .Q (new_AGEMA_signal_35059) ) ;
    buf_clk new_AGEMA_reg_buffer_14107 ( .C (clk), .D (new_AGEMA_signal_35062), .Q (new_AGEMA_signal_35063) ) ;
    buf_clk new_AGEMA_reg_buffer_14111 ( .C (clk), .D (new_AGEMA_signal_35066), .Q (new_AGEMA_signal_35067) ) ;
    buf_clk new_AGEMA_reg_buffer_14115 ( .C (clk), .D (new_AGEMA_signal_35070), .Q (new_AGEMA_signal_35071) ) ;
    buf_clk new_AGEMA_reg_buffer_14119 ( .C (clk), .D (new_AGEMA_signal_35074), .Q (new_AGEMA_signal_35075) ) ;
    buf_clk new_AGEMA_reg_buffer_14123 ( .C (clk), .D (new_AGEMA_signal_35078), .Q (new_AGEMA_signal_35079) ) ;
    buf_clk new_AGEMA_reg_buffer_14127 ( .C (clk), .D (new_AGEMA_signal_35082), .Q (new_AGEMA_signal_35083) ) ;
    buf_clk new_AGEMA_reg_buffer_14131 ( .C (clk), .D (new_AGEMA_signal_35086), .Q (new_AGEMA_signal_35087) ) ;
    buf_clk new_AGEMA_reg_buffer_14135 ( .C (clk), .D (new_AGEMA_signal_35090), .Q (new_AGEMA_signal_35091) ) ;
    buf_clk new_AGEMA_reg_buffer_14139 ( .C (clk), .D (new_AGEMA_signal_35094), .Q (new_AGEMA_signal_35095) ) ;
    buf_clk new_AGEMA_reg_buffer_14143 ( .C (clk), .D (new_AGEMA_signal_35098), .Q (new_AGEMA_signal_35099) ) ;
    buf_clk new_AGEMA_reg_buffer_14147 ( .C (clk), .D (new_AGEMA_signal_35102), .Q (new_AGEMA_signal_35103) ) ;
    buf_clk new_AGEMA_reg_buffer_14151 ( .C (clk), .D (new_AGEMA_signal_35106), .Q (new_AGEMA_signal_35107) ) ;
    buf_clk new_AGEMA_reg_buffer_14155 ( .C (clk), .D (new_AGEMA_signal_35110), .Q (new_AGEMA_signal_35111) ) ;
    buf_clk new_AGEMA_reg_buffer_14159 ( .C (clk), .D (new_AGEMA_signal_35114), .Q (new_AGEMA_signal_35115) ) ;
    buf_clk new_AGEMA_reg_buffer_14163 ( .C (clk), .D (new_AGEMA_signal_35118), .Q (new_AGEMA_signal_35119) ) ;
    buf_clk new_AGEMA_reg_buffer_14167 ( .C (clk), .D (new_AGEMA_signal_35122), .Q (new_AGEMA_signal_35123) ) ;
    buf_clk new_AGEMA_reg_buffer_14171 ( .C (clk), .D (new_AGEMA_signal_35126), .Q (new_AGEMA_signal_35127) ) ;
    buf_clk new_AGEMA_reg_buffer_14175 ( .C (clk), .D (new_AGEMA_signal_35130), .Q (new_AGEMA_signal_35131) ) ;
    buf_clk new_AGEMA_reg_buffer_14179 ( .C (clk), .D (new_AGEMA_signal_35134), .Q (new_AGEMA_signal_35135) ) ;
    buf_clk new_AGEMA_reg_buffer_14183 ( .C (clk), .D (new_AGEMA_signal_35138), .Q (new_AGEMA_signal_35139) ) ;
    buf_clk new_AGEMA_reg_buffer_14187 ( .C (clk), .D (new_AGEMA_signal_35142), .Q (new_AGEMA_signal_35143) ) ;
    buf_clk new_AGEMA_reg_buffer_14191 ( .C (clk), .D (new_AGEMA_signal_35146), .Q (new_AGEMA_signal_35147) ) ;
    buf_clk new_AGEMA_reg_buffer_14195 ( .C (clk), .D (new_AGEMA_signal_35150), .Q (new_AGEMA_signal_35151) ) ;
    buf_clk new_AGEMA_reg_buffer_14199 ( .C (clk), .D (new_AGEMA_signal_35154), .Q (new_AGEMA_signal_35155) ) ;
    buf_clk new_AGEMA_reg_buffer_14203 ( .C (clk), .D (new_AGEMA_signal_35158), .Q (new_AGEMA_signal_35159) ) ;
    buf_clk new_AGEMA_reg_buffer_14207 ( .C (clk), .D (new_AGEMA_signal_35162), .Q (new_AGEMA_signal_35163) ) ;
    buf_clk new_AGEMA_reg_buffer_14211 ( .C (clk), .D (new_AGEMA_signal_35166), .Q (new_AGEMA_signal_35167) ) ;
    buf_clk new_AGEMA_reg_buffer_14215 ( .C (clk), .D (new_AGEMA_signal_35170), .Q (new_AGEMA_signal_35171) ) ;
    buf_clk new_AGEMA_reg_buffer_14219 ( .C (clk), .D (new_AGEMA_signal_35174), .Q (new_AGEMA_signal_35175) ) ;
    buf_clk new_AGEMA_reg_buffer_14223 ( .C (clk), .D (new_AGEMA_signal_35178), .Q (new_AGEMA_signal_35179) ) ;
    buf_clk new_AGEMA_reg_buffer_14227 ( .C (clk), .D (new_AGEMA_signal_35182), .Q (new_AGEMA_signal_35183) ) ;
    buf_clk new_AGEMA_reg_buffer_14231 ( .C (clk), .D (new_AGEMA_signal_35186), .Q (new_AGEMA_signal_35187) ) ;
    buf_clk new_AGEMA_reg_buffer_14235 ( .C (clk), .D (new_AGEMA_signal_35190), .Q (new_AGEMA_signal_35191) ) ;
    buf_clk new_AGEMA_reg_buffer_14239 ( .C (clk), .D (new_AGEMA_signal_35194), .Q (new_AGEMA_signal_35195) ) ;
    buf_clk new_AGEMA_reg_buffer_14243 ( .C (clk), .D (new_AGEMA_signal_35198), .Q (new_AGEMA_signal_35199) ) ;
    buf_clk new_AGEMA_reg_buffer_14247 ( .C (clk), .D (new_AGEMA_signal_35202), .Q (new_AGEMA_signal_35203) ) ;
    buf_clk new_AGEMA_reg_buffer_14251 ( .C (clk), .D (new_AGEMA_signal_35206), .Q (new_AGEMA_signal_35207) ) ;
    buf_clk new_AGEMA_reg_buffer_14255 ( .C (clk), .D (new_AGEMA_signal_35210), .Q (new_AGEMA_signal_35211) ) ;
    buf_clk new_AGEMA_reg_buffer_14259 ( .C (clk), .D (new_AGEMA_signal_35214), .Q (new_AGEMA_signal_35215) ) ;
    buf_clk new_AGEMA_reg_buffer_14263 ( .C (clk), .D (new_AGEMA_signal_35218), .Q (new_AGEMA_signal_35219) ) ;
    buf_clk new_AGEMA_reg_buffer_14267 ( .C (clk), .D (new_AGEMA_signal_35222), .Q (new_AGEMA_signal_35223) ) ;
    buf_clk new_AGEMA_reg_buffer_14271 ( .C (clk), .D (new_AGEMA_signal_35226), .Q (new_AGEMA_signal_35227) ) ;
    buf_clk new_AGEMA_reg_buffer_14275 ( .C (clk), .D (new_AGEMA_signal_35230), .Q (new_AGEMA_signal_35231) ) ;
    buf_clk new_AGEMA_reg_buffer_14279 ( .C (clk), .D (new_AGEMA_signal_35234), .Q (new_AGEMA_signal_35235) ) ;
    buf_clk new_AGEMA_reg_buffer_14283 ( .C (clk), .D (new_AGEMA_signal_35238), .Q (new_AGEMA_signal_35239) ) ;
    buf_clk new_AGEMA_reg_buffer_14287 ( .C (clk), .D (new_AGEMA_signal_35242), .Q (new_AGEMA_signal_35243) ) ;
    buf_clk new_AGEMA_reg_buffer_14291 ( .C (clk), .D (new_AGEMA_signal_35246), .Q (new_AGEMA_signal_35247) ) ;
    buf_clk new_AGEMA_reg_buffer_14295 ( .C (clk), .D (new_AGEMA_signal_35250), .Q (new_AGEMA_signal_35251) ) ;
    buf_clk new_AGEMA_reg_buffer_14299 ( .C (clk), .D (new_AGEMA_signal_35254), .Q (new_AGEMA_signal_35255) ) ;
    buf_clk new_AGEMA_reg_buffer_14303 ( .C (clk), .D (new_AGEMA_signal_35258), .Q (new_AGEMA_signal_35259) ) ;
    buf_clk new_AGEMA_reg_buffer_14307 ( .C (clk), .D (new_AGEMA_signal_35262), .Q (new_AGEMA_signal_35263) ) ;
    buf_clk new_AGEMA_reg_buffer_14311 ( .C (clk), .D (new_AGEMA_signal_35266), .Q (new_AGEMA_signal_35267) ) ;
    buf_clk new_AGEMA_reg_buffer_14315 ( .C (clk), .D (new_AGEMA_signal_35270), .Q (new_AGEMA_signal_35271) ) ;
    buf_clk new_AGEMA_reg_buffer_14319 ( .C (clk), .D (new_AGEMA_signal_35274), .Q (new_AGEMA_signal_35275) ) ;
    buf_clk new_AGEMA_reg_buffer_14323 ( .C (clk), .D (new_AGEMA_signal_35278), .Q (new_AGEMA_signal_35279) ) ;
    buf_clk new_AGEMA_reg_buffer_14327 ( .C (clk), .D (new_AGEMA_signal_35282), .Q (new_AGEMA_signal_35283) ) ;
    buf_clk new_AGEMA_reg_buffer_14331 ( .C (clk), .D (new_AGEMA_signal_35286), .Q (new_AGEMA_signal_35287) ) ;
    buf_clk new_AGEMA_reg_buffer_14335 ( .C (clk), .D (new_AGEMA_signal_35290), .Q (new_AGEMA_signal_35291) ) ;
    buf_clk new_AGEMA_reg_buffer_14339 ( .C (clk), .D (new_AGEMA_signal_35294), .Q (new_AGEMA_signal_35295) ) ;
    buf_clk new_AGEMA_reg_buffer_14343 ( .C (clk), .D (new_AGEMA_signal_35298), .Q (new_AGEMA_signal_35299) ) ;
    buf_clk new_AGEMA_reg_buffer_14347 ( .C (clk), .D (new_AGEMA_signal_35302), .Q (new_AGEMA_signal_35303) ) ;
    buf_clk new_AGEMA_reg_buffer_14351 ( .C (clk), .D (new_AGEMA_signal_35306), .Q (new_AGEMA_signal_35307) ) ;
    buf_clk new_AGEMA_reg_buffer_14355 ( .C (clk), .D (new_AGEMA_signal_35310), .Q (new_AGEMA_signal_35311) ) ;
    buf_clk new_AGEMA_reg_buffer_14359 ( .C (clk), .D (new_AGEMA_signal_35314), .Q (new_AGEMA_signal_35315) ) ;
    buf_clk new_AGEMA_reg_buffer_14363 ( .C (clk), .D (new_AGEMA_signal_35318), .Q (new_AGEMA_signal_35319) ) ;
    buf_clk new_AGEMA_reg_buffer_14367 ( .C (clk), .D (new_AGEMA_signal_35322), .Q (new_AGEMA_signal_35323) ) ;
    buf_clk new_AGEMA_reg_buffer_14371 ( .C (clk), .D (new_AGEMA_signal_35326), .Q (new_AGEMA_signal_35327) ) ;
    buf_clk new_AGEMA_reg_buffer_14375 ( .C (clk), .D (new_AGEMA_signal_35330), .Q (new_AGEMA_signal_35331) ) ;
    buf_clk new_AGEMA_reg_buffer_14379 ( .C (clk), .D (new_AGEMA_signal_35334), .Q (new_AGEMA_signal_35335) ) ;
    buf_clk new_AGEMA_reg_buffer_14383 ( .C (clk), .D (new_AGEMA_signal_35338), .Q (new_AGEMA_signal_35339) ) ;
    buf_clk new_AGEMA_reg_buffer_14387 ( .C (clk), .D (new_AGEMA_signal_35342), .Q (new_AGEMA_signal_35343) ) ;
    buf_clk new_AGEMA_reg_buffer_14391 ( .C (clk), .D (new_AGEMA_signal_35346), .Q (new_AGEMA_signal_35347) ) ;
    buf_clk new_AGEMA_reg_buffer_14395 ( .C (clk), .D (new_AGEMA_signal_35350), .Q (new_AGEMA_signal_35351) ) ;
    buf_clk new_AGEMA_reg_buffer_14399 ( .C (clk), .D (new_AGEMA_signal_35354), .Q (new_AGEMA_signal_35355) ) ;
    buf_clk new_AGEMA_reg_buffer_14403 ( .C (clk), .D (new_AGEMA_signal_35358), .Q (new_AGEMA_signal_35359) ) ;
    buf_clk new_AGEMA_reg_buffer_14407 ( .C (clk), .D (new_AGEMA_signal_35362), .Q (new_AGEMA_signal_35363) ) ;
    buf_clk new_AGEMA_reg_buffer_14411 ( .C (clk), .D (new_AGEMA_signal_35366), .Q (new_AGEMA_signal_35367) ) ;
    buf_clk new_AGEMA_reg_buffer_14415 ( .C (clk), .D (new_AGEMA_signal_35370), .Q (new_AGEMA_signal_35371) ) ;
    buf_clk new_AGEMA_reg_buffer_14419 ( .C (clk), .D (new_AGEMA_signal_35374), .Q (new_AGEMA_signal_35375) ) ;
    buf_clk new_AGEMA_reg_buffer_14423 ( .C (clk), .D (new_AGEMA_signal_35378), .Q (new_AGEMA_signal_35379) ) ;
    buf_clk new_AGEMA_reg_buffer_14427 ( .C (clk), .D (new_AGEMA_signal_35382), .Q (new_AGEMA_signal_35383) ) ;
    buf_clk new_AGEMA_reg_buffer_14431 ( .C (clk), .D (new_AGEMA_signal_35386), .Q (new_AGEMA_signal_35387) ) ;
    buf_clk new_AGEMA_reg_buffer_14435 ( .C (clk), .D (new_AGEMA_signal_35390), .Q (new_AGEMA_signal_35391) ) ;
    buf_clk new_AGEMA_reg_buffer_14439 ( .C (clk), .D (new_AGEMA_signal_35394), .Q (new_AGEMA_signal_35395) ) ;
    buf_clk new_AGEMA_reg_buffer_14443 ( .C (clk), .D (new_AGEMA_signal_35398), .Q (new_AGEMA_signal_35399) ) ;
    buf_clk new_AGEMA_reg_buffer_14447 ( .C (clk), .D (new_AGEMA_signal_35402), .Q (new_AGEMA_signal_35403) ) ;
    buf_clk new_AGEMA_reg_buffer_14451 ( .C (clk), .D (new_AGEMA_signal_35406), .Q (new_AGEMA_signal_35407) ) ;
    buf_clk new_AGEMA_reg_buffer_14455 ( .C (clk), .D (new_AGEMA_signal_35410), .Q (new_AGEMA_signal_35411) ) ;
    buf_clk new_AGEMA_reg_buffer_14459 ( .C (clk), .D (new_AGEMA_signal_35414), .Q (new_AGEMA_signal_35415) ) ;
    buf_clk new_AGEMA_reg_buffer_14463 ( .C (clk), .D (new_AGEMA_signal_35418), .Q (new_AGEMA_signal_35419) ) ;
    buf_clk new_AGEMA_reg_buffer_14467 ( .C (clk), .D (new_AGEMA_signal_35422), .Q (new_AGEMA_signal_35423) ) ;
    buf_clk new_AGEMA_reg_buffer_14471 ( .C (clk), .D (new_AGEMA_signal_35426), .Q (new_AGEMA_signal_35427) ) ;
    buf_clk new_AGEMA_reg_buffer_14475 ( .C (clk), .D (new_AGEMA_signal_35430), .Q (new_AGEMA_signal_35431) ) ;
    buf_clk new_AGEMA_reg_buffer_14479 ( .C (clk), .D (new_AGEMA_signal_35434), .Q (new_AGEMA_signal_35435) ) ;
    buf_clk new_AGEMA_reg_buffer_14483 ( .C (clk), .D (new_AGEMA_signal_35438), .Q (new_AGEMA_signal_35439) ) ;
    buf_clk new_AGEMA_reg_buffer_14487 ( .C (clk), .D (new_AGEMA_signal_35442), .Q (new_AGEMA_signal_35443) ) ;
    buf_clk new_AGEMA_reg_buffer_14491 ( .C (clk), .D (new_AGEMA_signal_35446), .Q (new_AGEMA_signal_35447) ) ;
    buf_clk new_AGEMA_reg_buffer_14495 ( .C (clk), .D (new_AGEMA_signal_35450), .Q (new_AGEMA_signal_35451) ) ;
    buf_clk new_AGEMA_reg_buffer_14499 ( .C (clk), .D (new_AGEMA_signal_35454), .Q (new_AGEMA_signal_35455) ) ;
    buf_clk new_AGEMA_reg_buffer_14503 ( .C (clk), .D (new_AGEMA_signal_35458), .Q (new_AGEMA_signal_35459) ) ;
    buf_clk new_AGEMA_reg_buffer_14507 ( .C (clk), .D (new_AGEMA_signal_35462), .Q (new_AGEMA_signal_35463) ) ;
    buf_clk new_AGEMA_reg_buffer_14511 ( .C (clk), .D (new_AGEMA_signal_35466), .Q (new_AGEMA_signal_35467) ) ;
    buf_clk new_AGEMA_reg_buffer_14515 ( .C (clk), .D (new_AGEMA_signal_35470), .Q (new_AGEMA_signal_35471) ) ;
    buf_clk new_AGEMA_reg_buffer_14519 ( .C (clk), .D (new_AGEMA_signal_35474), .Q (new_AGEMA_signal_35475) ) ;
    buf_clk new_AGEMA_reg_buffer_14523 ( .C (clk), .D (new_AGEMA_signal_35478), .Q (new_AGEMA_signal_35479) ) ;
    buf_clk new_AGEMA_reg_buffer_14527 ( .C (clk), .D (new_AGEMA_signal_35482), .Q (new_AGEMA_signal_35483) ) ;
    buf_clk new_AGEMA_reg_buffer_14531 ( .C (clk), .D (new_AGEMA_signal_35486), .Q (new_AGEMA_signal_35487) ) ;
    buf_clk new_AGEMA_reg_buffer_14535 ( .C (clk), .D (new_AGEMA_signal_35490), .Q (new_AGEMA_signal_35491) ) ;
    buf_clk new_AGEMA_reg_buffer_14539 ( .C (clk), .D (new_AGEMA_signal_35494), .Q (new_AGEMA_signal_35495) ) ;
    buf_clk new_AGEMA_reg_buffer_14543 ( .C (clk), .D (new_AGEMA_signal_35498), .Q (new_AGEMA_signal_35499) ) ;
    buf_clk new_AGEMA_reg_buffer_14547 ( .C (clk), .D (new_AGEMA_signal_35502), .Q (new_AGEMA_signal_35503) ) ;
    buf_clk new_AGEMA_reg_buffer_14551 ( .C (clk), .D (new_AGEMA_signal_35506), .Q (new_AGEMA_signal_35507) ) ;
    buf_clk new_AGEMA_reg_buffer_14555 ( .C (clk), .D (new_AGEMA_signal_35510), .Q (new_AGEMA_signal_35511) ) ;
    buf_clk new_AGEMA_reg_buffer_14559 ( .C (clk), .D (new_AGEMA_signal_35514), .Q (new_AGEMA_signal_35515) ) ;
    buf_clk new_AGEMA_reg_buffer_14563 ( .C (clk), .D (new_AGEMA_signal_35518), .Q (new_AGEMA_signal_35519) ) ;
    buf_clk new_AGEMA_reg_buffer_14567 ( .C (clk), .D (new_AGEMA_signal_35522), .Q (new_AGEMA_signal_35523) ) ;
    buf_clk new_AGEMA_reg_buffer_14571 ( .C (clk), .D (new_AGEMA_signal_35526), .Q (new_AGEMA_signal_35527) ) ;
    buf_clk new_AGEMA_reg_buffer_14575 ( .C (clk), .D (new_AGEMA_signal_35530), .Q (new_AGEMA_signal_35531) ) ;
    buf_clk new_AGEMA_reg_buffer_14579 ( .C (clk), .D (new_AGEMA_signal_35534), .Q (new_AGEMA_signal_35535) ) ;
    buf_clk new_AGEMA_reg_buffer_14583 ( .C (clk), .D (new_AGEMA_signal_35538), .Q (new_AGEMA_signal_35539) ) ;
    buf_clk new_AGEMA_reg_buffer_14587 ( .C (clk), .D (new_AGEMA_signal_35542), .Q (new_AGEMA_signal_35543) ) ;
    buf_clk new_AGEMA_reg_buffer_14591 ( .C (clk), .D (new_AGEMA_signal_35546), .Q (new_AGEMA_signal_35547) ) ;
    buf_clk new_AGEMA_reg_buffer_14595 ( .C (clk), .D (new_AGEMA_signal_35550), .Q (new_AGEMA_signal_35551) ) ;
    buf_clk new_AGEMA_reg_buffer_14599 ( .C (clk), .D (new_AGEMA_signal_35554), .Q (new_AGEMA_signal_35555) ) ;
    buf_clk new_AGEMA_reg_buffer_14603 ( .C (clk), .D (new_AGEMA_signal_35558), .Q (new_AGEMA_signal_35559) ) ;
    buf_clk new_AGEMA_reg_buffer_14607 ( .C (clk), .D (new_AGEMA_signal_35562), .Q (new_AGEMA_signal_35563) ) ;
    buf_clk new_AGEMA_reg_buffer_14611 ( .C (clk), .D (new_AGEMA_signal_35566), .Q (new_AGEMA_signal_35567) ) ;
    buf_clk new_AGEMA_reg_buffer_14615 ( .C (clk), .D (new_AGEMA_signal_35570), .Q (new_AGEMA_signal_35571) ) ;
    buf_clk new_AGEMA_reg_buffer_14619 ( .C (clk), .D (new_AGEMA_signal_35574), .Q (new_AGEMA_signal_35575) ) ;
    buf_clk new_AGEMA_reg_buffer_14623 ( .C (clk), .D (new_AGEMA_signal_35578), .Q (new_AGEMA_signal_35579) ) ;
    buf_clk new_AGEMA_reg_buffer_14627 ( .C (clk), .D (new_AGEMA_signal_35582), .Q (new_AGEMA_signal_35583) ) ;
    buf_clk new_AGEMA_reg_buffer_14631 ( .C (clk), .D (new_AGEMA_signal_35586), .Q (new_AGEMA_signal_35587) ) ;
    buf_clk new_AGEMA_reg_buffer_14635 ( .C (clk), .D (new_AGEMA_signal_35590), .Q (new_AGEMA_signal_35591) ) ;
    buf_clk new_AGEMA_reg_buffer_14639 ( .C (clk), .D (new_AGEMA_signal_35594), .Q (new_AGEMA_signal_35595) ) ;
    buf_clk new_AGEMA_reg_buffer_14643 ( .C (clk), .D (new_AGEMA_signal_35598), .Q (new_AGEMA_signal_35599) ) ;
    buf_clk new_AGEMA_reg_buffer_14647 ( .C (clk), .D (new_AGEMA_signal_35602), .Q (new_AGEMA_signal_35603) ) ;
    buf_clk new_AGEMA_reg_buffer_14651 ( .C (clk), .D (new_AGEMA_signal_35606), .Q (new_AGEMA_signal_35607) ) ;
    buf_clk new_AGEMA_reg_buffer_14655 ( .C (clk), .D (new_AGEMA_signal_35610), .Q (new_AGEMA_signal_35611) ) ;
    buf_clk new_AGEMA_reg_buffer_14659 ( .C (clk), .D (new_AGEMA_signal_35614), .Q (new_AGEMA_signal_35615) ) ;
    buf_clk new_AGEMA_reg_buffer_14663 ( .C (clk), .D (new_AGEMA_signal_35618), .Q (new_AGEMA_signal_35619) ) ;
    buf_clk new_AGEMA_reg_buffer_14667 ( .C (clk), .D (new_AGEMA_signal_35622), .Q (new_AGEMA_signal_35623) ) ;
    buf_clk new_AGEMA_reg_buffer_14671 ( .C (clk), .D (new_AGEMA_signal_35626), .Q (new_AGEMA_signal_35627) ) ;
    buf_clk new_AGEMA_reg_buffer_14675 ( .C (clk), .D (new_AGEMA_signal_35630), .Q (new_AGEMA_signal_35631) ) ;
    buf_clk new_AGEMA_reg_buffer_14679 ( .C (clk), .D (new_AGEMA_signal_35634), .Q (new_AGEMA_signal_35635) ) ;
    buf_clk new_AGEMA_reg_buffer_14683 ( .C (clk), .D (new_AGEMA_signal_35638), .Q (new_AGEMA_signal_35639) ) ;
    buf_clk new_AGEMA_reg_buffer_14687 ( .C (clk), .D (new_AGEMA_signal_35642), .Q (new_AGEMA_signal_35643) ) ;
    buf_clk new_AGEMA_reg_buffer_14691 ( .C (clk), .D (new_AGEMA_signal_35646), .Q (new_AGEMA_signal_35647) ) ;
    buf_clk new_AGEMA_reg_buffer_14695 ( .C (clk), .D (new_AGEMA_signal_35650), .Q (new_AGEMA_signal_35651) ) ;
    buf_clk new_AGEMA_reg_buffer_14699 ( .C (clk), .D (new_AGEMA_signal_35654), .Q (new_AGEMA_signal_35655) ) ;
    buf_clk new_AGEMA_reg_buffer_14703 ( .C (clk), .D (new_AGEMA_signal_35658), .Q (new_AGEMA_signal_35659) ) ;
    buf_clk new_AGEMA_reg_buffer_14707 ( .C (clk), .D (new_AGEMA_signal_35662), .Q (new_AGEMA_signal_35663) ) ;
    buf_clk new_AGEMA_reg_buffer_14711 ( .C (clk), .D (new_AGEMA_signal_35666), .Q (new_AGEMA_signal_35667) ) ;
    buf_clk new_AGEMA_reg_buffer_14715 ( .C (clk), .D (new_AGEMA_signal_35670), .Q (new_AGEMA_signal_35671) ) ;
    buf_clk new_AGEMA_reg_buffer_14719 ( .C (clk), .D (new_AGEMA_signal_35674), .Q (new_AGEMA_signal_35675) ) ;
    buf_clk new_AGEMA_reg_buffer_14723 ( .C (clk), .D (new_AGEMA_signal_35678), .Q (new_AGEMA_signal_35679) ) ;
    buf_clk new_AGEMA_reg_buffer_14727 ( .C (clk), .D (new_AGEMA_signal_35682), .Q (new_AGEMA_signal_35683) ) ;
    buf_clk new_AGEMA_reg_buffer_14731 ( .C (clk), .D (new_AGEMA_signal_35686), .Q (new_AGEMA_signal_35687) ) ;
    buf_clk new_AGEMA_reg_buffer_14735 ( .C (clk), .D (new_AGEMA_signal_35690), .Q (new_AGEMA_signal_35691) ) ;
    buf_clk new_AGEMA_reg_buffer_14739 ( .C (clk), .D (new_AGEMA_signal_35694), .Q (new_AGEMA_signal_35695) ) ;
    buf_clk new_AGEMA_reg_buffer_14743 ( .C (clk), .D (new_AGEMA_signal_35698), .Q (new_AGEMA_signal_35699) ) ;
    buf_clk new_AGEMA_reg_buffer_14747 ( .C (clk), .D (new_AGEMA_signal_35702), .Q (new_AGEMA_signal_35703) ) ;
    buf_clk new_AGEMA_reg_buffer_14751 ( .C (clk), .D (new_AGEMA_signal_35706), .Q (new_AGEMA_signal_35707) ) ;
    buf_clk new_AGEMA_reg_buffer_14755 ( .C (clk), .D (new_AGEMA_signal_35710), .Q (new_AGEMA_signal_35711) ) ;
    buf_clk new_AGEMA_reg_buffer_14759 ( .C (clk), .D (new_AGEMA_signal_35714), .Q (new_AGEMA_signal_35715) ) ;
    buf_clk new_AGEMA_reg_buffer_14763 ( .C (clk), .D (new_AGEMA_signal_35718), .Q (new_AGEMA_signal_35719) ) ;
    buf_clk new_AGEMA_reg_buffer_14767 ( .C (clk), .D (new_AGEMA_signal_35722), .Q (new_AGEMA_signal_35723) ) ;
    buf_clk new_AGEMA_reg_buffer_14771 ( .C (clk), .D (new_AGEMA_signal_35726), .Q (new_AGEMA_signal_35727) ) ;
    buf_clk new_AGEMA_reg_buffer_14775 ( .C (clk), .D (new_AGEMA_signal_35730), .Q (new_AGEMA_signal_35731) ) ;
    buf_clk new_AGEMA_reg_buffer_14779 ( .C (clk), .D (new_AGEMA_signal_35734), .Q (new_AGEMA_signal_35735) ) ;
    buf_clk new_AGEMA_reg_buffer_14783 ( .C (clk), .D (new_AGEMA_signal_35738), .Q (new_AGEMA_signal_35739) ) ;
    buf_clk new_AGEMA_reg_buffer_14787 ( .C (clk), .D (new_AGEMA_signal_35742), .Q (new_AGEMA_signal_35743) ) ;
    buf_clk new_AGEMA_reg_buffer_14791 ( .C (clk), .D (new_AGEMA_signal_35746), .Q (new_AGEMA_signal_35747) ) ;
    buf_clk new_AGEMA_reg_buffer_14795 ( .C (clk), .D (new_AGEMA_signal_35750), .Q (new_AGEMA_signal_35751) ) ;
    buf_clk new_AGEMA_reg_buffer_14799 ( .C (clk), .D (new_AGEMA_signal_35754), .Q (new_AGEMA_signal_35755) ) ;
    buf_clk new_AGEMA_reg_buffer_14803 ( .C (clk), .D (new_AGEMA_signal_35758), .Q (new_AGEMA_signal_35759) ) ;
    buf_clk new_AGEMA_reg_buffer_14807 ( .C (clk), .D (new_AGEMA_signal_35762), .Q (new_AGEMA_signal_35763) ) ;
    buf_clk new_AGEMA_reg_buffer_14811 ( .C (clk), .D (new_AGEMA_signal_35766), .Q (new_AGEMA_signal_35767) ) ;
    buf_clk new_AGEMA_reg_buffer_14815 ( .C (clk), .D (new_AGEMA_signal_35770), .Q (new_AGEMA_signal_35771) ) ;
    buf_clk new_AGEMA_reg_buffer_14819 ( .C (clk), .D (new_AGEMA_signal_35774), .Q (new_AGEMA_signal_35775) ) ;
    buf_clk new_AGEMA_reg_buffer_14823 ( .C (clk), .D (new_AGEMA_signal_35778), .Q (new_AGEMA_signal_35779) ) ;
    buf_clk new_AGEMA_reg_buffer_14827 ( .C (clk), .D (new_AGEMA_signal_35782), .Q (new_AGEMA_signal_35783) ) ;
    buf_clk new_AGEMA_reg_buffer_14831 ( .C (clk), .D (new_AGEMA_signal_35786), .Q (new_AGEMA_signal_35787) ) ;
    buf_clk new_AGEMA_reg_buffer_14835 ( .C (clk), .D (new_AGEMA_signal_35790), .Q (new_AGEMA_signal_35791) ) ;
    buf_clk new_AGEMA_reg_buffer_14838 ( .C (clk), .D (new_AGEMA_signal_35793), .Q (new_AGEMA_signal_35794) ) ;
    buf_clk new_AGEMA_reg_buffer_14841 ( .C (clk), .D (new_AGEMA_signal_35796), .Q (new_AGEMA_signal_35797) ) ;
    buf_clk new_AGEMA_reg_buffer_14844 ( .C (clk), .D (new_AGEMA_signal_35799), .Q (new_AGEMA_signal_35800) ) ;
    buf_clk new_AGEMA_reg_buffer_14847 ( .C (clk), .D (new_AGEMA_signal_35802), .Q (new_AGEMA_signal_35803) ) ;
    buf_clk new_AGEMA_reg_buffer_14850 ( .C (clk), .D (new_AGEMA_signal_35805), .Q (new_AGEMA_signal_35806) ) ;
    buf_clk new_AGEMA_reg_buffer_14853 ( .C (clk), .D (new_AGEMA_signal_35808), .Q (new_AGEMA_signal_35809) ) ;
    buf_clk new_AGEMA_reg_buffer_14856 ( .C (clk), .D (new_AGEMA_signal_35811), .Q (new_AGEMA_signal_35812) ) ;
    buf_clk new_AGEMA_reg_buffer_14859 ( .C (clk), .D (new_AGEMA_signal_35814), .Q (new_AGEMA_signal_35815) ) ;
    buf_clk new_AGEMA_reg_buffer_14862 ( .C (clk), .D (new_AGEMA_signal_35817), .Q (new_AGEMA_signal_35818) ) ;
    buf_clk new_AGEMA_reg_buffer_14865 ( .C (clk), .D (new_AGEMA_signal_35820), .Q (new_AGEMA_signal_35821) ) ;
    buf_clk new_AGEMA_reg_buffer_14868 ( .C (clk), .D (new_AGEMA_signal_35823), .Q (new_AGEMA_signal_35824) ) ;
    buf_clk new_AGEMA_reg_buffer_14871 ( .C (clk), .D (new_AGEMA_signal_35826), .Q (new_AGEMA_signal_35827) ) ;
    buf_clk new_AGEMA_reg_buffer_14874 ( .C (clk), .D (new_AGEMA_signal_35829), .Q (new_AGEMA_signal_35830) ) ;
    buf_clk new_AGEMA_reg_buffer_14877 ( .C (clk), .D (new_AGEMA_signal_35832), .Q (new_AGEMA_signal_35833) ) ;
    buf_clk new_AGEMA_reg_buffer_14880 ( .C (clk), .D (new_AGEMA_signal_35835), .Q (new_AGEMA_signal_35836) ) ;
    buf_clk new_AGEMA_reg_buffer_14883 ( .C (clk), .D (new_AGEMA_signal_35838), .Q (new_AGEMA_signal_35839) ) ;
    buf_clk new_AGEMA_reg_buffer_14886 ( .C (clk), .D (new_AGEMA_signal_35841), .Q (new_AGEMA_signal_35842) ) ;
    buf_clk new_AGEMA_reg_buffer_14889 ( .C (clk), .D (new_AGEMA_signal_35844), .Q (new_AGEMA_signal_35845) ) ;
    buf_clk new_AGEMA_reg_buffer_14892 ( .C (clk), .D (new_AGEMA_signal_35847), .Q (new_AGEMA_signal_35848) ) ;
    buf_clk new_AGEMA_reg_buffer_14895 ( .C (clk), .D (new_AGEMA_signal_35850), .Q (new_AGEMA_signal_35851) ) ;
    buf_clk new_AGEMA_reg_buffer_14898 ( .C (clk), .D (new_AGEMA_signal_35853), .Q (new_AGEMA_signal_35854) ) ;
    buf_clk new_AGEMA_reg_buffer_14901 ( .C (clk), .D (new_AGEMA_signal_35856), .Q (new_AGEMA_signal_35857) ) ;
    buf_clk new_AGEMA_reg_buffer_14904 ( .C (clk), .D (new_AGEMA_signal_35859), .Q (new_AGEMA_signal_35860) ) ;
    buf_clk new_AGEMA_reg_buffer_14907 ( .C (clk), .D (new_AGEMA_signal_35862), .Q (new_AGEMA_signal_35863) ) ;
    buf_clk new_AGEMA_reg_buffer_14910 ( .C (clk), .D (new_AGEMA_signal_35865), .Q (new_AGEMA_signal_35866) ) ;
    buf_clk new_AGEMA_reg_buffer_14913 ( .C (clk), .D (new_AGEMA_signal_35868), .Q (new_AGEMA_signal_35869) ) ;
    buf_clk new_AGEMA_reg_buffer_14916 ( .C (clk), .D (new_AGEMA_signal_35871), .Q (new_AGEMA_signal_35872) ) ;
    buf_clk new_AGEMA_reg_buffer_14919 ( .C (clk), .D (new_AGEMA_signal_35874), .Q (new_AGEMA_signal_35875) ) ;
    buf_clk new_AGEMA_reg_buffer_14922 ( .C (clk), .D (new_AGEMA_signal_35877), .Q (new_AGEMA_signal_35878) ) ;
    buf_clk new_AGEMA_reg_buffer_14925 ( .C (clk), .D (new_AGEMA_signal_35880), .Q (new_AGEMA_signal_35881) ) ;
    buf_clk new_AGEMA_reg_buffer_14928 ( .C (clk), .D (new_AGEMA_signal_35883), .Q (new_AGEMA_signal_35884) ) ;
    buf_clk new_AGEMA_reg_buffer_14931 ( .C (clk), .D (new_AGEMA_signal_35886), .Q (new_AGEMA_signal_35887) ) ;
    buf_clk new_AGEMA_reg_buffer_14934 ( .C (clk), .D (new_AGEMA_signal_35889), .Q (new_AGEMA_signal_35890) ) ;
    buf_clk new_AGEMA_reg_buffer_14937 ( .C (clk), .D (new_AGEMA_signal_35892), .Q (new_AGEMA_signal_35893) ) ;
    buf_clk new_AGEMA_reg_buffer_14940 ( .C (clk), .D (new_AGEMA_signal_35895), .Q (new_AGEMA_signal_35896) ) ;
    buf_clk new_AGEMA_reg_buffer_14943 ( .C (clk), .D (new_AGEMA_signal_35898), .Q (new_AGEMA_signal_35899) ) ;
    buf_clk new_AGEMA_reg_buffer_14946 ( .C (clk), .D (new_AGEMA_signal_35901), .Q (new_AGEMA_signal_35902) ) ;
    buf_clk new_AGEMA_reg_buffer_14949 ( .C (clk), .D (new_AGEMA_signal_35904), .Q (new_AGEMA_signal_35905) ) ;
    buf_clk new_AGEMA_reg_buffer_14952 ( .C (clk), .D (new_AGEMA_signal_35907), .Q (new_AGEMA_signal_35908) ) ;
    buf_clk new_AGEMA_reg_buffer_14955 ( .C (clk), .D (new_AGEMA_signal_35910), .Q (new_AGEMA_signal_35911) ) ;
    buf_clk new_AGEMA_reg_buffer_14958 ( .C (clk), .D (new_AGEMA_signal_35913), .Q (new_AGEMA_signal_35914) ) ;
    buf_clk new_AGEMA_reg_buffer_14961 ( .C (clk), .D (new_AGEMA_signal_35916), .Q (new_AGEMA_signal_35917) ) ;
    buf_clk new_AGEMA_reg_buffer_14964 ( .C (clk), .D (new_AGEMA_signal_35919), .Q (new_AGEMA_signal_35920) ) ;
    buf_clk new_AGEMA_reg_buffer_14967 ( .C (clk), .D (new_AGEMA_signal_35922), .Q (new_AGEMA_signal_35923) ) ;
    buf_clk new_AGEMA_reg_buffer_14970 ( .C (clk), .D (new_AGEMA_signal_35925), .Q (new_AGEMA_signal_35926) ) ;
    buf_clk new_AGEMA_reg_buffer_14973 ( .C (clk), .D (new_AGEMA_signal_35928), .Q (new_AGEMA_signal_35929) ) ;
    buf_clk new_AGEMA_reg_buffer_14976 ( .C (clk), .D (new_AGEMA_signal_35931), .Q (new_AGEMA_signal_35932) ) ;
    buf_clk new_AGEMA_reg_buffer_14979 ( .C (clk), .D (new_AGEMA_signal_35934), .Q (new_AGEMA_signal_35935) ) ;
    buf_clk new_AGEMA_reg_buffer_14982 ( .C (clk), .D (new_AGEMA_signal_35937), .Q (new_AGEMA_signal_35938) ) ;
    buf_clk new_AGEMA_reg_buffer_14985 ( .C (clk), .D (new_AGEMA_signal_35940), .Q (new_AGEMA_signal_35941) ) ;
    buf_clk new_AGEMA_reg_buffer_14988 ( .C (clk), .D (new_AGEMA_signal_35943), .Q (new_AGEMA_signal_35944) ) ;
    buf_clk new_AGEMA_reg_buffer_14991 ( .C (clk), .D (new_AGEMA_signal_35946), .Q (new_AGEMA_signal_35947) ) ;
    buf_clk new_AGEMA_reg_buffer_14994 ( .C (clk), .D (new_AGEMA_signal_35949), .Q (new_AGEMA_signal_35950) ) ;
    buf_clk new_AGEMA_reg_buffer_14997 ( .C (clk), .D (new_AGEMA_signal_35952), .Q (new_AGEMA_signal_35953) ) ;
    buf_clk new_AGEMA_reg_buffer_15000 ( .C (clk), .D (new_AGEMA_signal_35955), .Q (new_AGEMA_signal_35956) ) ;
    buf_clk new_AGEMA_reg_buffer_15003 ( .C (clk), .D (new_AGEMA_signal_35958), .Q (new_AGEMA_signal_35959) ) ;
    buf_clk new_AGEMA_reg_buffer_15006 ( .C (clk), .D (new_AGEMA_signal_35961), .Q (new_AGEMA_signal_35962) ) ;
    buf_clk new_AGEMA_reg_buffer_15009 ( .C (clk), .D (new_AGEMA_signal_35964), .Q (new_AGEMA_signal_35965) ) ;
    buf_clk new_AGEMA_reg_buffer_15012 ( .C (clk), .D (new_AGEMA_signal_35967), .Q (new_AGEMA_signal_35968) ) ;
    buf_clk new_AGEMA_reg_buffer_15015 ( .C (clk), .D (new_AGEMA_signal_35970), .Q (new_AGEMA_signal_35971) ) ;
    buf_clk new_AGEMA_reg_buffer_15018 ( .C (clk), .D (new_AGEMA_signal_35973), .Q (new_AGEMA_signal_35974) ) ;
    buf_clk new_AGEMA_reg_buffer_15021 ( .C (clk), .D (new_AGEMA_signal_35976), .Q (new_AGEMA_signal_35977) ) ;
    buf_clk new_AGEMA_reg_buffer_15024 ( .C (clk), .D (new_AGEMA_signal_35979), .Q (new_AGEMA_signal_35980) ) ;
    buf_clk new_AGEMA_reg_buffer_15027 ( .C (clk), .D (new_AGEMA_signal_35982), .Q (new_AGEMA_signal_35983) ) ;
    buf_clk new_AGEMA_reg_buffer_15030 ( .C (clk), .D (new_AGEMA_signal_35985), .Q (new_AGEMA_signal_35986) ) ;
    buf_clk new_AGEMA_reg_buffer_15033 ( .C (clk), .D (new_AGEMA_signal_35988), .Q (new_AGEMA_signal_35989) ) ;
    buf_clk new_AGEMA_reg_buffer_15036 ( .C (clk), .D (new_AGEMA_signal_35991), .Q (new_AGEMA_signal_35992) ) ;
    buf_clk new_AGEMA_reg_buffer_15039 ( .C (clk), .D (new_AGEMA_signal_35994), .Q (new_AGEMA_signal_35995) ) ;
    buf_clk new_AGEMA_reg_buffer_15042 ( .C (clk), .D (new_AGEMA_signal_35997), .Q (new_AGEMA_signal_35998) ) ;
    buf_clk new_AGEMA_reg_buffer_15045 ( .C (clk), .D (new_AGEMA_signal_36000), .Q (new_AGEMA_signal_36001) ) ;
    buf_clk new_AGEMA_reg_buffer_15048 ( .C (clk), .D (new_AGEMA_signal_36003), .Q (new_AGEMA_signal_36004) ) ;
    buf_clk new_AGEMA_reg_buffer_15051 ( .C (clk), .D (new_AGEMA_signal_36006), .Q (new_AGEMA_signal_36007) ) ;
    buf_clk new_AGEMA_reg_buffer_15054 ( .C (clk), .D (new_AGEMA_signal_36009), .Q (new_AGEMA_signal_36010) ) ;
    buf_clk new_AGEMA_reg_buffer_15057 ( .C (clk), .D (new_AGEMA_signal_36012), .Q (new_AGEMA_signal_36013) ) ;
    buf_clk new_AGEMA_reg_buffer_15060 ( .C (clk), .D (new_AGEMA_signal_36015), .Q (new_AGEMA_signal_36016) ) ;
    buf_clk new_AGEMA_reg_buffer_15063 ( .C (clk), .D (new_AGEMA_signal_36018), .Q (new_AGEMA_signal_36019) ) ;
    buf_clk new_AGEMA_reg_buffer_15066 ( .C (clk), .D (new_AGEMA_signal_36021), .Q (new_AGEMA_signal_36022) ) ;
    buf_clk new_AGEMA_reg_buffer_15069 ( .C (clk), .D (new_AGEMA_signal_36024), .Q (new_AGEMA_signal_36025) ) ;
    buf_clk new_AGEMA_reg_buffer_15072 ( .C (clk), .D (new_AGEMA_signal_36027), .Q (new_AGEMA_signal_36028) ) ;
    buf_clk new_AGEMA_reg_buffer_15075 ( .C (clk), .D (new_AGEMA_signal_36030), .Q (new_AGEMA_signal_36031) ) ;
    buf_clk new_AGEMA_reg_buffer_15078 ( .C (clk), .D (new_AGEMA_signal_36033), .Q (new_AGEMA_signal_36034) ) ;
    buf_clk new_AGEMA_reg_buffer_15081 ( .C (clk), .D (new_AGEMA_signal_36036), .Q (new_AGEMA_signal_36037) ) ;
    buf_clk new_AGEMA_reg_buffer_15084 ( .C (clk), .D (new_AGEMA_signal_36039), .Q (new_AGEMA_signal_36040) ) ;
    buf_clk new_AGEMA_reg_buffer_15087 ( .C (clk), .D (new_AGEMA_signal_36042), .Q (new_AGEMA_signal_36043) ) ;
    buf_clk new_AGEMA_reg_buffer_15090 ( .C (clk), .D (new_AGEMA_signal_36045), .Q (new_AGEMA_signal_36046) ) ;
    buf_clk new_AGEMA_reg_buffer_15093 ( .C (clk), .D (new_AGEMA_signal_36048), .Q (new_AGEMA_signal_36049) ) ;
    buf_clk new_AGEMA_reg_buffer_15096 ( .C (clk), .D (new_AGEMA_signal_36051), .Q (new_AGEMA_signal_36052) ) ;
    buf_clk new_AGEMA_reg_buffer_15099 ( .C (clk), .D (new_AGEMA_signal_36054), .Q (new_AGEMA_signal_36055) ) ;
    buf_clk new_AGEMA_reg_buffer_15102 ( .C (clk), .D (new_AGEMA_signal_36057), .Q (new_AGEMA_signal_36058) ) ;
    buf_clk new_AGEMA_reg_buffer_15105 ( .C (clk), .D (new_AGEMA_signal_36060), .Q (new_AGEMA_signal_36061) ) ;
    buf_clk new_AGEMA_reg_buffer_15108 ( .C (clk), .D (new_AGEMA_signal_36063), .Q (new_AGEMA_signal_36064) ) ;
    buf_clk new_AGEMA_reg_buffer_15111 ( .C (clk), .D (new_AGEMA_signal_36066), .Q (new_AGEMA_signal_36067) ) ;
    buf_clk new_AGEMA_reg_buffer_15114 ( .C (clk), .D (new_AGEMA_signal_36069), .Q (new_AGEMA_signal_36070) ) ;
    buf_clk new_AGEMA_reg_buffer_15117 ( .C (clk), .D (new_AGEMA_signal_36072), .Q (new_AGEMA_signal_36073) ) ;
    buf_clk new_AGEMA_reg_buffer_15120 ( .C (clk), .D (new_AGEMA_signal_36075), .Q (new_AGEMA_signal_36076) ) ;
    buf_clk new_AGEMA_reg_buffer_15123 ( .C (clk), .D (new_AGEMA_signal_36078), .Q (new_AGEMA_signal_36079) ) ;
    buf_clk new_AGEMA_reg_buffer_15126 ( .C (clk), .D (new_AGEMA_signal_36081), .Q (new_AGEMA_signal_36082) ) ;
    buf_clk new_AGEMA_reg_buffer_15129 ( .C (clk), .D (new_AGEMA_signal_36084), .Q (new_AGEMA_signal_36085) ) ;
    buf_clk new_AGEMA_reg_buffer_15132 ( .C (clk), .D (new_AGEMA_signal_36087), .Q (new_AGEMA_signal_36088) ) ;
    buf_clk new_AGEMA_reg_buffer_15135 ( .C (clk), .D (new_AGEMA_signal_36090), .Q (new_AGEMA_signal_36091) ) ;
    buf_clk new_AGEMA_reg_buffer_15138 ( .C (clk), .D (new_AGEMA_signal_36093), .Q (new_AGEMA_signal_36094) ) ;
    buf_clk new_AGEMA_reg_buffer_15141 ( .C (clk), .D (new_AGEMA_signal_36096), .Q (new_AGEMA_signal_36097) ) ;
    buf_clk new_AGEMA_reg_buffer_15144 ( .C (clk), .D (new_AGEMA_signal_36099), .Q (new_AGEMA_signal_36100) ) ;
    buf_clk new_AGEMA_reg_buffer_15147 ( .C (clk), .D (new_AGEMA_signal_36102), .Q (new_AGEMA_signal_36103) ) ;
    buf_clk new_AGEMA_reg_buffer_15150 ( .C (clk), .D (new_AGEMA_signal_36105), .Q (new_AGEMA_signal_36106) ) ;
    buf_clk new_AGEMA_reg_buffer_15153 ( .C (clk), .D (new_AGEMA_signal_36108), .Q (new_AGEMA_signal_36109) ) ;
    buf_clk new_AGEMA_reg_buffer_15156 ( .C (clk), .D (new_AGEMA_signal_36111), .Q (new_AGEMA_signal_36112) ) ;
    buf_clk new_AGEMA_reg_buffer_15159 ( .C (clk), .D (new_AGEMA_signal_36114), .Q (new_AGEMA_signal_36115) ) ;
    buf_clk new_AGEMA_reg_buffer_15162 ( .C (clk), .D (new_AGEMA_signal_36117), .Q (new_AGEMA_signal_36118) ) ;
    buf_clk new_AGEMA_reg_buffer_15165 ( .C (clk), .D (new_AGEMA_signal_36120), .Q (new_AGEMA_signal_36121) ) ;
    buf_clk new_AGEMA_reg_buffer_15168 ( .C (clk), .D (new_AGEMA_signal_36123), .Q (new_AGEMA_signal_36124) ) ;
    buf_clk new_AGEMA_reg_buffer_15171 ( .C (clk), .D (new_AGEMA_signal_36126), .Q (new_AGEMA_signal_36127) ) ;
    buf_clk new_AGEMA_reg_buffer_15174 ( .C (clk), .D (new_AGEMA_signal_36129), .Q (new_AGEMA_signal_36130) ) ;
    buf_clk new_AGEMA_reg_buffer_15177 ( .C (clk), .D (new_AGEMA_signal_36132), .Q (new_AGEMA_signal_36133) ) ;
    buf_clk new_AGEMA_reg_buffer_15180 ( .C (clk), .D (new_AGEMA_signal_36135), .Q (new_AGEMA_signal_36136) ) ;
    buf_clk new_AGEMA_reg_buffer_15183 ( .C (clk), .D (new_AGEMA_signal_36138), .Q (new_AGEMA_signal_36139) ) ;
    buf_clk new_AGEMA_reg_buffer_15186 ( .C (clk), .D (new_AGEMA_signal_36141), .Q (new_AGEMA_signal_36142) ) ;
    buf_clk new_AGEMA_reg_buffer_15189 ( .C (clk), .D (new_AGEMA_signal_36144), .Q (new_AGEMA_signal_36145) ) ;
    buf_clk new_AGEMA_reg_buffer_15192 ( .C (clk), .D (new_AGEMA_signal_36147), .Q (new_AGEMA_signal_36148) ) ;
    buf_clk new_AGEMA_reg_buffer_15195 ( .C (clk), .D (new_AGEMA_signal_36150), .Q (new_AGEMA_signal_36151) ) ;
    buf_clk new_AGEMA_reg_buffer_15198 ( .C (clk), .D (new_AGEMA_signal_36153), .Q (new_AGEMA_signal_36154) ) ;
    buf_clk new_AGEMA_reg_buffer_15201 ( .C (clk), .D (new_AGEMA_signal_36156), .Q (new_AGEMA_signal_36157) ) ;
    buf_clk new_AGEMA_reg_buffer_15204 ( .C (clk), .D (new_AGEMA_signal_36159), .Q (new_AGEMA_signal_36160) ) ;
    buf_clk new_AGEMA_reg_buffer_15207 ( .C (clk), .D (new_AGEMA_signal_36162), .Q (new_AGEMA_signal_36163) ) ;
    buf_clk new_AGEMA_reg_buffer_15210 ( .C (clk), .D (new_AGEMA_signal_36165), .Q (new_AGEMA_signal_36166) ) ;
    buf_clk new_AGEMA_reg_buffer_15213 ( .C (clk), .D (new_AGEMA_signal_36168), .Q (new_AGEMA_signal_36169) ) ;
    buf_clk new_AGEMA_reg_buffer_15216 ( .C (clk), .D (new_AGEMA_signal_36171), .Q (new_AGEMA_signal_36172) ) ;
    buf_clk new_AGEMA_reg_buffer_15219 ( .C (clk), .D (new_AGEMA_signal_36174), .Q (new_AGEMA_signal_36175) ) ;
    buf_clk new_AGEMA_reg_buffer_15222 ( .C (clk), .D (new_AGEMA_signal_36177), .Q (new_AGEMA_signal_36178) ) ;
    buf_clk new_AGEMA_reg_buffer_15225 ( .C (clk), .D (new_AGEMA_signal_36180), .Q (new_AGEMA_signal_36181) ) ;
    buf_clk new_AGEMA_reg_buffer_15228 ( .C (clk), .D (new_AGEMA_signal_36183), .Q (new_AGEMA_signal_36184) ) ;
    buf_clk new_AGEMA_reg_buffer_15231 ( .C (clk), .D (new_AGEMA_signal_36186), .Q (new_AGEMA_signal_36187) ) ;
    buf_clk new_AGEMA_reg_buffer_15234 ( .C (clk), .D (new_AGEMA_signal_36189), .Q (new_AGEMA_signal_36190) ) ;
    buf_clk new_AGEMA_reg_buffer_15237 ( .C (clk), .D (new_AGEMA_signal_36192), .Q (new_AGEMA_signal_36193) ) ;
    buf_clk new_AGEMA_reg_buffer_15240 ( .C (clk), .D (new_AGEMA_signal_36195), .Q (new_AGEMA_signal_36196) ) ;
    buf_clk new_AGEMA_reg_buffer_15243 ( .C (clk), .D (new_AGEMA_signal_36198), .Q (new_AGEMA_signal_36199) ) ;
    buf_clk new_AGEMA_reg_buffer_15246 ( .C (clk), .D (new_AGEMA_signal_36201), .Q (new_AGEMA_signal_36202) ) ;
    buf_clk new_AGEMA_reg_buffer_15249 ( .C (clk), .D (new_AGEMA_signal_36204), .Q (new_AGEMA_signal_36205) ) ;
    buf_clk new_AGEMA_reg_buffer_15252 ( .C (clk), .D (new_AGEMA_signal_36207), .Q (new_AGEMA_signal_36208) ) ;
    buf_clk new_AGEMA_reg_buffer_15255 ( .C (clk), .D (new_AGEMA_signal_36210), .Q (new_AGEMA_signal_36211) ) ;
    buf_clk new_AGEMA_reg_buffer_15258 ( .C (clk), .D (new_AGEMA_signal_36213), .Q (new_AGEMA_signal_36214) ) ;
    buf_clk new_AGEMA_reg_buffer_15261 ( .C (clk), .D (new_AGEMA_signal_36216), .Q (new_AGEMA_signal_36217) ) ;
    buf_clk new_AGEMA_reg_buffer_15264 ( .C (clk), .D (new_AGEMA_signal_36219), .Q (new_AGEMA_signal_36220) ) ;
    buf_clk new_AGEMA_reg_buffer_15267 ( .C (clk), .D (new_AGEMA_signal_36222), .Q (new_AGEMA_signal_36223) ) ;
    buf_clk new_AGEMA_reg_buffer_15270 ( .C (clk), .D (new_AGEMA_signal_36225), .Q (new_AGEMA_signal_36226) ) ;
    buf_clk new_AGEMA_reg_buffer_15273 ( .C (clk), .D (new_AGEMA_signal_36228), .Q (new_AGEMA_signal_36229) ) ;
    buf_clk new_AGEMA_reg_buffer_15276 ( .C (clk), .D (new_AGEMA_signal_36231), .Q (new_AGEMA_signal_36232) ) ;
    buf_clk new_AGEMA_reg_buffer_15279 ( .C (clk), .D (new_AGEMA_signal_36234), .Q (new_AGEMA_signal_36235) ) ;
    buf_clk new_AGEMA_reg_buffer_15282 ( .C (clk), .D (new_AGEMA_signal_36237), .Q (new_AGEMA_signal_36238) ) ;
    buf_clk new_AGEMA_reg_buffer_15285 ( .C (clk), .D (new_AGEMA_signal_36240), .Q (new_AGEMA_signal_36241) ) ;
    buf_clk new_AGEMA_reg_buffer_15288 ( .C (clk), .D (new_AGEMA_signal_36243), .Q (new_AGEMA_signal_36244) ) ;
    buf_clk new_AGEMA_reg_buffer_15291 ( .C (clk), .D (new_AGEMA_signal_36246), .Q (new_AGEMA_signal_36247) ) ;
    buf_clk new_AGEMA_reg_buffer_15294 ( .C (clk), .D (new_AGEMA_signal_36249), .Q (new_AGEMA_signal_36250) ) ;
    buf_clk new_AGEMA_reg_buffer_15297 ( .C (clk), .D (new_AGEMA_signal_36252), .Q (new_AGEMA_signal_36253) ) ;
    buf_clk new_AGEMA_reg_buffer_15300 ( .C (clk), .D (new_AGEMA_signal_36255), .Q (new_AGEMA_signal_36256) ) ;
    buf_clk new_AGEMA_reg_buffer_15303 ( .C (clk), .D (new_AGEMA_signal_36258), .Q (new_AGEMA_signal_36259) ) ;
    buf_clk new_AGEMA_reg_buffer_15306 ( .C (clk), .D (new_AGEMA_signal_36261), .Q (new_AGEMA_signal_36262) ) ;
    buf_clk new_AGEMA_reg_buffer_15309 ( .C (clk), .D (new_AGEMA_signal_36264), .Q (new_AGEMA_signal_36265) ) ;
    buf_clk new_AGEMA_reg_buffer_15312 ( .C (clk), .D (new_AGEMA_signal_36267), .Q (new_AGEMA_signal_36268) ) ;
    buf_clk new_AGEMA_reg_buffer_15315 ( .C (clk), .D (new_AGEMA_signal_36270), .Q (new_AGEMA_signal_36271) ) ;
    buf_clk new_AGEMA_reg_buffer_15318 ( .C (clk), .D (new_AGEMA_signal_36273), .Q (new_AGEMA_signal_36274) ) ;
    buf_clk new_AGEMA_reg_buffer_15321 ( .C (clk), .D (new_AGEMA_signal_36276), .Q (new_AGEMA_signal_36277) ) ;
    buf_clk new_AGEMA_reg_buffer_15324 ( .C (clk), .D (new_AGEMA_signal_36279), .Q (new_AGEMA_signal_36280) ) ;
    buf_clk new_AGEMA_reg_buffer_15327 ( .C (clk), .D (new_AGEMA_signal_36282), .Q (new_AGEMA_signal_36283) ) ;
    buf_clk new_AGEMA_reg_buffer_15330 ( .C (clk), .D (new_AGEMA_signal_36285), .Q (new_AGEMA_signal_36286) ) ;
    buf_clk new_AGEMA_reg_buffer_15333 ( .C (clk), .D (new_AGEMA_signal_36288), .Q (new_AGEMA_signal_36289) ) ;
    buf_clk new_AGEMA_reg_buffer_15336 ( .C (clk), .D (new_AGEMA_signal_36291), .Q (new_AGEMA_signal_36292) ) ;
    buf_clk new_AGEMA_reg_buffer_15339 ( .C (clk), .D (new_AGEMA_signal_36294), .Q (new_AGEMA_signal_36295) ) ;
    buf_clk new_AGEMA_reg_buffer_15342 ( .C (clk), .D (new_AGEMA_signal_36297), .Q (new_AGEMA_signal_36298) ) ;
    buf_clk new_AGEMA_reg_buffer_15345 ( .C (clk), .D (new_AGEMA_signal_36300), .Q (new_AGEMA_signal_36301) ) ;
    buf_clk new_AGEMA_reg_buffer_15348 ( .C (clk), .D (new_AGEMA_signal_36303), .Q (new_AGEMA_signal_36304) ) ;
    buf_clk new_AGEMA_reg_buffer_15351 ( .C (clk), .D (new_AGEMA_signal_36306), .Q (new_AGEMA_signal_36307) ) ;
    buf_clk new_AGEMA_reg_buffer_15354 ( .C (clk), .D (new_AGEMA_signal_36309), .Q (new_AGEMA_signal_36310) ) ;
    buf_clk new_AGEMA_reg_buffer_15357 ( .C (clk), .D (new_AGEMA_signal_36312), .Q (new_AGEMA_signal_36313) ) ;
    buf_clk new_AGEMA_reg_buffer_15360 ( .C (clk), .D (new_AGEMA_signal_36315), .Q (new_AGEMA_signal_36316) ) ;
    buf_clk new_AGEMA_reg_buffer_15363 ( .C (clk), .D (new_AGEMA_signal_36318), .Q (new_AGEMA_signal_36319) ) ;
    buf_clk new_AGEMA_reg_buffer_15366 ( .C (clk), .D (new_AGEMA_signal_36321), .Q (new_AGEMA_signal_36322) ) ;
    buf_clk new_AGEMA_reg_buffer_15369 ( .C (clk), .D (new_AGEMA_signal_36324), .Q (new_AGEMA_signal_36325) ) ;
    buf_clk new_AGEMA_reg_buffer_15372 ( .C (clk), .D (new_AGEMA_signal_36327), .Q (new_AGEMA_signal_36328) ) ;
    buf_clk new_AGEMA_reg_buffer_15375 ( .C (clk), .D (new_AGEMA_signal_36330), .Q (new_AGEMA_signal_36331) ) ;
    buf_clk new_AGEMA_reg_buffer_15378 ( .C (clk), .D (new_AGEMA_signal_36333), .Q (new_AGEMA_signal_36334) ) ;
    buf_clk new_AGEMA_reg_buffer_15381 ( .C (clk), .D (new_AGEMA_signal_36336), .Q (new_AGEMA_signal_36337) ) ;
    buf_clk new_AGEMA_reg_buffer_15384 ( .C (clk), .D (new_AGEMA_signal_36339), .Q (new_AGEMA_signal_36340) ) ;
    buf_clk new_AGEMA_reg_buffer_15387 ( .C (clk), .D (new_AGEMA_signal_36342), .Q (new_AGEMA_signal_36343) ) ;
    buf_clk new_AGEMA_reg_buffer_15390 ( .C (clk), .D (new_AGEMA_signal_36345), .Q (new_AGEMA_signal_36346) ) ;
    buf_clk new_AGEMA_reg_buffer_15393 ( .C (clk), .D (new_AGEMA_signal_36348), .Q (new_AGEMA_signal_36349) ) ;
    buf_clk new_AGEMA_reg_buffer_15396 ( .C (clk), .D (new_AGEMA_signal_36351), .Q (new_AGEMA_signal_36352) ) ;
    buf_clk new_AGEMA_reg_buffer_15399 ( .C (clk), .D (new_AGEMA_signal_36354), .Q (new_AGEMA_signal_36355) ) ;
    buf_clk new_AGEMA_reg_buffer_15402 ( .C (clk), .D (new_AGEMA_signal_36357), .Q (new_AGEMA_signal_36358) ) ;
    buf_clk new_AGEMA_reg_buffer_15405 ( .C (clk), .D (new_AGEMA_signal_36360), .Q (new_AGEMA_signal_36361) ) ;
    buf_clk new_AGEMA_reg_buffer_15408 ( .C (clk), .D (new_AGEMA_signal_36363), .Q (new_AGEMA_signal_36364) ) ;
    buf_clk new_AGEMA_reg_buffer_15411 ( .C (clk), .D (new_AGEMA_signal_36366), .Q (new_AGEMA_signal_36367) ) ;
    buf_clk new_AGEMA_reg_buffer_15414 ( .C (clk), .D (new_AGEMA_signal_36369), .Q (new_AGEMA_signal_36370) ) ;
    buf_clk new_AGEMA_reg_buffer_15417 ( .C (clk), .D (new_AGEMA_signal_36372), .Q (new_AGEMA_signal_36373) ) ;
    buf_clk new_AGEMA_reg_buffer_15420 ( .C (clk), .D (new_AGEMA_signal_36375), .Q (new_AGEMA_signal_36376) ) ;
    buf_clk new_AGEMA_reg_buffer_15423 ( .C (clk), .D (new_AGEMA_signal_36378), .Q (new_AGEMA_signal_36379) ) ;
    buf_clk new_AGEMA_reg_buffer_15426 ( .C (clk), .D (new_AGEMA_signal_36381), .Q (new_AGEMA_signal_36382) ) ;
    buf_clk new_AGEMA_reg_buffer_15429 ( .C (clk), .D (new_AGEMA_signal_36384), .Q (new_AGEMA_signal_36385) ) ;
    buf_clk new_AGEMA_reg_buffer_15432 ( .C (clk), .D (new_AGEMA_signal_36387), .Q (new_AGEMA_signal_36388) ) ;
    buf_clk new_AGEMA_reg_buffer_15435 ( .C (clk), .D (new_AGEMA_signal_36390), .Q (new_AGEMA_signal_36391) ) ;
    buf_clk new_AGEMA_reg_buffer_15438 ( .C (clk), .D (new_AGEMA_signal_36393), .Q (new_AGEMA_signal_36394) ) ;
    buf_clk new_AGEMA_reg_buffer_15441 ( .C (clk), .D (new_AGEMA_signal_36396), .Q (new_AGEMA_signal_36397) ) ;
    buf_clk new_AGEMA_reg_buffer_15444 ( .C (clk), .D (new_AGEMA_signal_36399), .Q (new_AGEMA_signal_36400) ) ;
    buf_clk new_AGEMA_reg_buffer_15447 ( .C (clk), .D (new_AGEMA_signal_36402), .Q (new_AGEMA_signal_36403) ) ;
    buf_clk new_AGEMA_reg_buffer_15450 ( .C (clk), .D (new_AGEMA_signal_36405), .Q (new_AGEMA_signal_36406) ) ;
    buf_clk new_AGEMA_reg_buffer_15453 ( .C (clk), .D (new_AGEMA_signal_36408), .Q (new_AGEMA_signal_36409) ) ;
    buf_clk new_AGEMA_reg_buffer_15456 ( .C (clk), .D (new_AGEMA_signal_36411), .Q (new_AGEMA_signal_36412) ) ;
    buf_clk new_AGEMA_reg_buffer_15459 ( .C (clk), .D (new_AGEMA_signal_36414), .Q (new_AGEMA_signal_36415) ) ;
    buf_clk new_AGEMA_reg_buffer_15462 ( .C (clk), .D (new_AGEMA_signal_36417), .Q (new_AGEMA_signal_36418) ) ;
    buf_clk new_AGEMA_reg_buffer_15465 ( .C (clk), .D (new_AGEMA_signal_36420), .Q (new_AGEMA_signal_36421) ) ;
    buf_clk new_AGEMA_reg_buffer_15468 ( .C (clk), .D (new_AGEMA_signal_36423), .Q (new_AGEMA_signal_36424) ) ;
    buf_clk new_AGEMA_reg_buffer_15471 ( .C (clk), .D (new_AGEMA_signal_36426), .Q (new_AGEMA_signal_36427) ) ;
    buf_clk new_AGEMA_reg_buffer_15474 ( .C (clk), .D (new_AGEMA_signal_36429), .Q (new_AGEMA_signal_36430) ) ;
    buf_clk new_AGEMA_reg_buffer_15477 ( .C (clk), .D (new_AGEMA_signal_36432), .Q (new_AGEMA_signal_36433) ) ;
    buf_clk new_AGEMA_reg_buffer_15480 ( .C (clk), .D (new_AGEMA_signal_36435), .Q (new_AGEMA_signal_36436) ) ;
    buf_clk new_AGEMA_reg_buffer_15483 ( .C (clk), .D (new_AGEMA_signal_36438), .Q (new_AGEMA_signal_36439) ) ;
    buf_clk new_AGEMA_reg_buffer_15486 ( .C (clk), .D (new_AGEMA_signal_36441), .Q (new_AGEMA_signal_36442) ) ;
    buf_clk new_AGEMA_reg_buffer_15489 ( .C (clk), .D (new_AGEMA_signal_36444), .Q (new_AGEMA_signal_36445) ) ;
    buf_clk new_AGEMA_reg_buffer_15492 ( .C (clk), .D (new_AGEMA_signal_36447), .Q (new_AGEMA_signal_36448) ) ;
    buf_clk new_AGEMA_reg_buffer_15495 ( .C (clk), .D (new_AGEMA_signal_36450), .Q (new_AGEMA_signal_36451) ) ;
    buf_clk new_AGEMA_reg_buffer_15498 ( .C (clk), .D (new_AGEMA_signal_36453), .Q (new_AGEMA_signal_36454) ) ;
    buf_clk new_AGEMA_reg_buffer_15501 ( .C (clk), .D (new_AGEMA_signal_36456), .Q (new_AGEMA_signal_36457) ) ;
    buf_clk new_AGEMA_reg_buffer_15504 ( .C (clk), .D (new_AGEMA_signal_36459), .Q (new_AGEMA_signal_36460) ) ;
    buf_clk new_AGEMA_reg_buffer_15507 ( .C (clk), .D (new_AGEMA_signal_36462), .Q (new_AGEMA_signal_36463) ) ;
    buf_clk new_AGEMA_reg_buffer_15510 ( .C (clk), .D (new_AGEMA_signal_36465), .Q (new_AGEMA_signal_36466) ) ;
    buf_clk new_AGEMA_reg_buffer_15513 ( .C (clk), .D (new_AGEMA_signal_36468), .Q (new_AGEMA_signal_36469) ) ;
    buf_clk new_AGEMA_reg_buffer_15516 ( .C (clk), .D (new_AGEMA_signal_36471), .Q (new_AGEMA_signal_36472) ) ;
    buf_clk new_AGEMA_reg_buffer_15519 ( .C (clk), .D (new_AGEMA_signal_36474), .Q (new_AGEMA_signal_36475) ) ;
    buf_clk new_AGEMA_reg_buffer_15522 ( .C (clk), .D (new_AGEMA_signal_36477), .Q (new_AGEMA_signal_36478) ) ;
    buf_clk new_AGEMA_reg_buffer_15525 ( .C (clk), .D (new_AGEMA_signal_36480), .Q (new_AGEMA_signal_36481) ) ;
    buf_clk new_AGEMA_reg_buffer_15528 ( .C (clk), .D (new_AGEMA_signal_36483), .Q (new_AGEMA_signal_36484) ) ;
    buf_clk new_AGEMA_reg_buffer_15531 ( .C (clk), .D (new_AGEMA_signal_36486), .Q (new_AGEMA_signal_36487) ) ;
    buf_clk new_AGEMA_reg_buffer_15534 ( .C (clk), .D (new_AGEMA_signal_36489), .Q (new_AGEMA_signal_36490) ) ;
    buf_clk new_AGEMA_reg_buffer_15537 ( .C (clk), .D (new_AGEMA_signal_36492), .Q (new_AGEMA_signal_36493) ) ;
    buf_clk new_AGEMA_reg_buffer_15540 ( .C (clk), .D (new_AGEMA_signal_36495), .Q (new_AGEMA_signal_36496) ) ;
    buf_clk new_AGEMA_reg_buffer_15543 ( .C (clk), .D (new_AGEMA_signal_36498), .Q (new_AGEMA_signal_36499) ) ;
    buf_clk new_AGEMA_reg_buffer_15546 ( .C (clk), .D (new_AGEMA_signal_36501), .Q (new_AGEMA_signal_36502) ) ;
    buf_clk new_AGEMA_reg_buffer_15549 ( .C (clk), .D (new_AGEMA_signal_36504), .Q (new_AGEMA_signal_36505) ) ;
    buf_clk new_AGEMA_reg_buffer_15552 ( .C (clk), .D (new_AGEMA_signal_36507), .Q (new_AGEMA_signal_36508) ) ;
    buf_clk new_AGEMA_reg_buffer_15555 ( .C (clk), .D (new_AGEMA_signal_36510), .Q (new_AGEMA_signal_36511) ) ;
    buf_clk new_AGEMA_reg_buffer_15558 ( .C (clk), .D (new_AGEMA_signal_36513), .Q (new_AGEMA_signal_36514) ) ;
    buf_clk new_AGEMA_reg_buffer_15561 ( .C (clk), .D (new_AGEMA_signal_36516), .Q (new_AGEMA_signal_36517) ) ;
    buf_clk new_AGEMA_reg_buffer_15564 ( .C (clk), .D (new_AGEMA_signal_36519), .Q (new_AGEMA_signal_36520) ) ;
    buf_clk new_AGEMA_reg_buffer_15567 ( .C (clk), .D (new_AGEMA_signal_36522), .Q (new_AGEMA_signal_36523) ) ;
    buf_clk new_AGEMA_reg_buffer_15570 ( .C (clk), .D (new_AGEMA_signal_36525), .Q (new_AGEMA_signal_36526) ) ;
    buf_clk new_AGEMA_reg_buffer_15573 ( .C (clk), .D (new_AGEMA_signal_36528), .Q (new_AGEMA_signal_36529) ) ;
    buf_clk new_AGEMA_reg_buffer_15576 ( .C (clk), .D (new_AGEMA_signal_36531), .Q (new_AGEMA_signal_36532) ) ;
    buf_clk new_AGEMA_reg_buffer_15579 ( .C (clk), .D (new_AGEMA_signal_36534), .Q (new_AGEMA_signal_36535) ) ;
    buf_clk new_AGEMA_reg_buffer_15582 ( .C (clk), .D (new_AGEMA_signal_36537), .Q (new_AGEMA_signal_36538) ) ;
    buf_clk new_AGEMA_reg_buffer_15585 ( .C (clk), .D (new_AGEMA_signal_36540), .Q (new_AGEMA_signal_36541) ) ;
    buf_clk new_AGEMA_reg_buffer_15588 ( .C (clk), .D (new_AGEMA_signal_36543), .Q (new_AGEMA_signal_36544) ) ;
    buf_clk new_AGEMA_reg_buffer_15591 ( .C (clk), .D (new_AGEMA_signal_36546), .Q (new_AGEMA_signal_36547) ) ;
    buf_clk new_AGEMA_reg_buffer_15594 ( .C (clk), .D (new_AGEMA_signal_36549), .Q (new_AGEMA_signal_36550) ) ;
    buf_clk new_AGEMA_reg_buffer_15597 ( .C (clk), .D (new_AGEMA_signal_36552), .Q (new_AGEMA_signal_36553) ) ;
    buf_clk new_AGEMA_reg_buffer_15600 ( .C (clk), .D (new_AGEMA_signal_36555), .Q (new_AGEMA_signal_36556) ) ;
    buf_clk new_AGEMA_reg_buffer_15603 ( .C (clk), .D (new_AGEMA_signal_36558), .Q (new_AGEMA_signal_36559) ) ;
    buf_clk new_AGEMA_reg_buffer_15606 ( .C (clk), .D (new_AGEMA_signal_36561), .Q (new_AGEMA_signal_36562) ) ;
    buf_clk new_AGEMA_reg_buffer_15609 ( .C (clk), .D (new_AGEMA_signal_36564), .Q (new_AGEMA_signal_36565) ) ;
    buf_clk new_AGEMA_reg_buffer_15612 ( .C (clk), .D (new_AGEMA_signal_36567), .Q (new_AGEMA_signal_36568) ) ;
    buf_clk new_AGEMA_reg_buffer_15615 ( .C (clk), .D (new_AGEMA_signal_36570), .Q (new_AGEMA_signal_36571) ) ;
    buf_clk new_AGEMA_reg_buffer_15618 ( .C (clk), .D (new_AGEMA_signal_36573), .Q (new_AGEMA_signal_36574) ) ;
    buf_clk new_AGEMA_reg_buffer_15621 ( .C (clk), .D (new_AGEMA_signal_36576), .Q (new_AGEMA_signal_36577) ) ;
    buf_clk new_AGEMA_reg_buffer_15624 ( .C (clk), .D (new_AGEMA_signal_36579), .Q (new_AGEMA_signal_36580) ) ;
    buf_clk new_AGEMA_reg_buffer_15627 ( .C (clk), .D (new_AGEMA_signal_36582), .Q (new_AGEMA_signal_36583) ) ;
    buf_clk new_AGEMA_reg_buffer_15630 ( .C (clk), .D (new_AGEMA_signal_36585), .Q (new_AGEMA_signal_36586) ) ;
    buf_clk new_AGEMA_reg_buffer_15633 ( .C (clk), .D (new_AGEMA_signal_36588), .Q (new_AGEMA_signal_36589) ) ;
    buf_clk new_AGEMA_reg_buffer_15636 ( .C (clk), .D (new_AGEMA_signal_36591), .Q (new_AGEMA_signal_36592) ) ;
    buf_clk new_AGEMA_reg_buffer_15639 ( .C (clk), .D (new_AGEMA_signal_36594), .Q (new_AGEMA_signal_36595) ) ;
    buf_clk new_AGEMA_reg_buffer_15642 ( .C (clk), .D (new_AGEMA_signal_36597), .Q (new_AGEMA_signal_36598) ) ;
    buf_clk new_AGEMA_reg_buffer_15645 ( .C (clk), .D (new_AGEMA_signal_36600), .Q (new_AGEMA_signal_36601) ) ;
    buf_clk new_AGEMA_reg_buffer_15648 ( .C (clk), .D (new_AGEMA_signal_36603), .Q (new_AGEMA_signal_36604) ) ;
    buf_clk new_AGEMA_reg_buffer_15651 ( .C (clk), .D (new_AGEMA_signal_36606), .Q (new_AGEMA_signal_36607) ) ;
    buf_clk new_AGEMA_reg_buffer_15655 ( .C (clk), .D (new_AGEMA_signal_36610), .Q (new_AGEMA_signal_36611) ) ;
    buf_clk new_AGEMA_reg_buffer_15659 ( .C (clk), .D (new_AGEMA_signal_36614), .Q (new_AGEMA_signal_36615) ) ;
    buf_clk new_AGEMA_reg_buffer_15663 ( .C (clk), .D (new_AGEMA_signal_36618), .Q (new_AGEMA_signal_36619) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(3), .pipeline(1)) U858 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .a ({new_AGEMA_signal_15192, new_AGEMA_signal_15191, new_AGEMA_signal_15190, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_15474, new_AGEMA_signal_15473, new_AGEMA_signal_15472, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U859 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, new_AGEMA_signal_15715, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_16053, new_AGEMA_signal_16052, new_AGEMA_signal_16051, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U860 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_14823, new_AGEMA_signal_14822, new_AGEMA_signal_14821, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_15477, new_AGEMA_signal_15476, new_AGEMA_signal_15475, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U861 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_14820, new_AGEMA_signal_14819, new_AGEMA_signal_14818, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_15480, new_AGEMA_signal_15479, new_AGEMA_signal_15478, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U862 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_14817, new_AGEMA_signal_14816, new_AGEMA_signal_14815, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_15483, new_AGEMA_signal_15482, new_AGEMA_signal_15481, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U863 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .a ({new_AGEMA_signal_14814, new_AGEMA_signal_14813, new_AGEMA_signal_14812, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_15486, new_AGEMA_signal_15485, new_AGEMA_signal_15484, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U864 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_15714, new_AGEMA_signal_15713, new_AGEMA_signal_15712, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_16056, new_AGEMA_signal_16055, new_AGEMA_signal_16054, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U865 ( .s (new_AGEMA_signal_26128), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .a ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, new_AGEMA_signal_14899, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, new_AGEMA_signal_15487, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U866 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .a ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, new_AGEMA_signal_15745, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, new_AGEMA_signal_16057, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U867 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_15744, new_AGEMA_signal_15743, new_AGEMA_signal_15742, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_16062, new_AGEMA_signal_16061, new_AGEMA_signal_16060, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U868 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_14892, new_AGEMA_signal_14891, new_AGEMA_signal_14890, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_15492, new_AGEMA_signal_15491, new_AGEMA_signal_15490, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U869 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .a ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, new_AGEMA_signal_15187, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, new_AGEMA_signal_15493, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U870 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_14889, new_AGEMA_signal_14888, new_AGEMA_signal_14887, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_15498, new_AGEMA_signal_15497, new_AGEMA_signal_15496, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U871 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_14886, new_AGEMA_signal_14885, new_AGEMA_signal_14884, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, new_AGEMA_signal_15499, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U872 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .a ({new_AGEMA_signal_14883, new_AGEMA_signal_14882, new_AGEMA_signal_14881, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_15504, new_AGEMA_signal_15503, new_AGEMA_signal_15502, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U873 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, new_AGEMA_signal_15739, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, new_AGEMA_signal_16063, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U874 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .a ({new_AGEMA_signal_14877, new_AGEMA_signal_14876, new_AGEMA_signal_14875, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_15507, new_AGEMA_signal_15506, new_AGEMA_signal_15505, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U875 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .a ({new_AGEMA_signal_15738, new_AGEMA_signal_15737, new_AGEMA_signal_15736, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_16068, new_AGEMA_signal_16067, new_AGEMA_signal_16066, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U876 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_15732, new_AGEMA_signal_15731, new_AGEMA_signal_15730, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, new_AGEMA_signal_16069, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U877 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_14865, new_AGEMA_signal_14864, new_AGEMA_signal_14863, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_15510, new_AGEMA_signal_15509, new_AGEMA_signal_15508, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U878 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_14862, new_AGEMA_signal_14861, new_AGEMA_signal_14860, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_15513, new_AGEMA_signal_15512, new_AGEMA_signal_15511, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U879 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, new_AGEMA_signal_14857, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_15516, new_AGEMA_signal_15515, new_AGEMA_signal_15514, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U880 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .a ({new_AGEMA_signal_15855, new_AGEMA_signal_15854, new_AGEMA_signal_15853, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_16074, new_AGEMA_signal_16073, new_AGEMA_signal_16072, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U881 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .a ({new_AGEMA_signal_14856, new_AGEMA_signal_14855, new_AGEMA_signal_14854, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, new_AGEMA_signal_15517, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U882 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_15729, new_AGEMA_signal_15728, new_AGEMA_signal_15727, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_16077, new_AGEMA_signal_16076, new_AGEMA_signal_16075, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U883 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .a ({new_AGEMA_signal_14850, new_AGEMA_signal_14849, new_AGEMA_signal_14848, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_15522, new_AGEMA_signal_15521, new_AGEMA_signal_15520, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U884 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .a ({new_AGEMA_signal_15726, new_AGEMA_signal_15725, new_AGEMA_signal_15724, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_16080, new_AGEMA_signal_16079, new_AGEMA_signal_16078, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U885 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, new_AGEMA_signal_15721, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, new_AGEMA_signal_16081, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U886 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, new_AGEMA_signal_14839, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, new_AGEMA_signal_15523, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U887 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, new_AGEMA_signal_14833, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_15528, new_AGEMA_signal_15527, new_AGEMA_signal_15526, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U888 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_14832, new_AGEMA_signal_14831, new_AGEMA_signal_14830, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, new_AGEMA_signal_15529, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U889 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_15852, new_AGEMA_signal_15851, new_AGEMA_signal_15850, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_16086, new_AGEMA_signal_16085, new_AGEMA_signal_16084, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U890 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_15180, new_AGEMA_signal_15179, new_AGEMA_signal_15178, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_15534, new_AGEMA_signal_15533, new_AGEMA_signal_15532, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U891 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_15177, new_AGEMA_signal_15176, new_AGEMA_signal_15175, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, new_AGEMA_signal_15535, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U892 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_15174, new_AGEMA_signal_15173, new_AGEMA_signal_15172, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_15540, new_AGEMA_signal_15539, new_AGEMA_signal_15538, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U893 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .a ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, new_AGEMA_signal_15169, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_15543, new_AGEMA_signal_15542, new_AGEMA_signal_15541, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U894 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, new_AGEMA_signal_15847, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, new_AGEMA_signal_16087, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U895 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .a ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, new_AGEMA_signal_15163, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_15546, new_AGEMA_signal_15545, new_AGEMA_signal_15544, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U896 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .a ({new_AGEMA_signal_15846, new_AGEMA_signal_15845, new_AGEMA_signal_15844, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_16092, new_AGEMA_signal_16091, new_AGEMA_signal_16090, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U897 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, new_AGEMA_signal_15841, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, new_AGEMA_signal_16093, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U898 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_15840, new_AGEMA_signal_15839, new_AGEMA_signal_15838, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_16098, new_AGEMA_signal_16097, new_AGEMA_signal_16096, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U899 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, new_AGEMA_signal_15151, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, new_AGEMA_signal_15547, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U900 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_15150, new_AGEMA_signal_15149, new_AGEMA_signal_15148, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_15552, new_AGEMA_signal_15551, new_AGEMA_signal_15550, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U901 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, new_AGEMA_signal_15145, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, new_AGEMA_signal_15553, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U902 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .a ({new_AGEMA_signal_15144, new_AGEMA_signal_15143, new_AGEMA_signal_15142, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_15558, new_AGEMA_signal_15557, new_AGEMA_signal_15556, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U903 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, new_AGEMA_signal_15835, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, new_AGEMA_signal_16099, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U904 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .a ({new_AGEMA_signal_15138, new_AGEMA_signal_15137, new_AGEMA_signal_15136, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, new_AGEMA_signal_15559, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U905 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .a ({new_AGEMA_signal_15834, new_AGEMA_signal_15833, new_AGEMA_signal_15832, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_16104, new_AGEMA_signal_16103, new_AGEMA_signal_16102, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U906 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, new_AGEMA_signal_15829, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, new_AGEMA_signal_16105, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U907 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, new_AGEMA_signal_15127, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_15564, new_AGEMA_signal_15563, new_AGEMA_signal_15562, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U908 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .a ({new_AGEMA_signal_15126, new_AGEMA_signal_15125, new_AGEMA_signal_15124, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, new_AGEMA_signal_15565, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U909 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, new_AGEMA_signal_15121, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_15570, new_AGEMA_signal_15569, new_AGEMA_signal_15568, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U910 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_15120, new_AGEMA_signal_15119, new_AGEMA_signal_15118, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, new_AGEMA_signal_15571, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U911 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .a ({new_AGEMA_signal_15096, new_AGEMA_signal_15095, new_AGEMA_signal_15094, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_15576, new_AGEMA_signal_15575, new_AGEMA_signal_15574, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U912 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, new_AGEMA_signal_15805, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_16110, new_AGEMA_signal_16109, new_AGEMA_signal_16108, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U913 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .a ({new_AGEMA_signal_15030, new_AGEMA_signal_15029, new_AGEMA_signal_15028, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, new_AGEMA_signal_15577, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U914 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .a ({new_AGEMA_signal_15792, new_AGEMA_signal_15791, new_AGEMA_signal_15790, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_16113, new_AGEMA_signal_16112, new_AGEMA_signal_16111, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U915 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_15789, new_AGEMA_signal_15788, new_AGEMA_signal_15787, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_16116, new_AGEMA_signal_16115, new_AGEMA_signal_16114, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U916 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, new_AGEMA_signal_15013, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_15582, new_AGEMA_signal_15581, new_AGEMA_signal_15580, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U917 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_15012, new_AGEMA_signal_15011, new_AGEMA_signal_15010, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, new_AGEMA_signal_15583, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U918 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, new_AGEMA_signal_15007, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_15588, new_AGEMA_signal_15587, new_AGEMA_signal_15586, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U919 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .a ({new_AGEMA_signal_15828, new_AGEMA_signal_15827, new_AGEMA_signal_15826, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, new_AGEMA_signal_16117, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U920 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .a ({new_AGEMA_signal_15006, new_AGEMA_signal_15005, new_AGEMA_signal_15004, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_15591, new_AGEMA_signal_15590, new_AGEMA_signal_15589, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U921 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_15786, new_AGEMA_signal_15785, new_AGEMA_signal_15784, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_16122, new_AGEMA_signal_16121, new_AGEMA_signal_16120, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U922 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .a ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, new_AGEMA_signal_15091, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_15594, new_AGEMA_signal_15593, new_AGEMA_signal_15592, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U923 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .a ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, new_AGEMA_signal_15817, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_16125, new_AGEMA_signal_16124, new_AGEMA_signal_16123, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U924 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_15816, new_AGEMA_signal_15815, new_AGEMA_signal_15814, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_16128, new_AGEMA_signal_16127, new_AGEMA_signal_16126, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U925 ( .s (new_AGEMA_signal_26152), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_15084, new_AGEMA_signal_15083, new_AGEMA_signal_15082, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_15597, new_AGEMA_signal_15596, new_AGEMA_signal_15595, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U926 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, new_AGEMA_signal_15079, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_15600, new_AGEMA_signal_15599, new_AGEMA_signal_15598, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U927 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_15078, new_AGEMA_signal_15077, new_AGEMA_signal_15076, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, new_AGEMA_signal_15601, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U928 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .a ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, new_AGEMA_signal_15073, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_15606, new_AGEMA_signal_15605, new_AGEMA_signal_15604, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U929 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, new_AGEMA_signal_15811, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_16131, new_AGEMA_signal_16130, new_AGEMA_signal_16129, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U930 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, new_AGEMA_signal_15823, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_16134, new_AGEMA_signal_16133, new_AGEMA_signal_16132, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U931 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .a ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, new_AGEMA_signal_15067, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, new_AGEMA_signal_15607, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U932 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .a ({new_AGEMA_signal_15810, new_AGEMA_signal_15809, new_AGEMA_signal_15808, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, new_AGEMA_signal_16135, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U933 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_15804, new_AGEMA_signal_15803, new_AGEMA_signal_15802, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_16140, new_AGEMA_signal_16139, new_AGEMA_signal_16138, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U934 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, new_AGEMA_signal_15055, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_15612, new_AGEMA_signal_15611, new_AGEMA_signal_15610, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U935 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_15054, new_AGEMA_signal_15053, new_AGEMA_signal_15052, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_15615, new_AGEMA_signal_15614, new_AGEMA_signal_15613, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U936 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, new_AGEMA_signal_15049, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_15618, new_AGEMA_signal_15617, new_AGEMA_signal_15616, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U937 ( .s (new_AGEMA_signal_26148), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .a ({new_AGEMA_signal_15048, new_AGEMA_signal_15047, new_AGEMA_signal_15046, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, new_AGEMA_signal_15619, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U938 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, new_AGEMA_signal_15799, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_16143, new_AGEMA_signal_16142, new_AGEMA_signal_16141, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U939 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .a ({new_AGEMA_signal_15042, new_AGEMA_signal_15041, new_AGEMA_signal_15040, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_15624, new_AGEMA_signal_15623, new_AGEMA_signal_15622, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U940 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .a ({new_AGEMA_signal_15798, new_AGEMA_signal_15797, new_AGEMA_signal_15796, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_16146, new_AGEMA_signal_16145, new_AGEMA_signal_16144, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U941 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, new_AGEMA_signal_15109, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, new_AGEMA_signal_15625, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U942 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_15795, new_AGEMA_signal_15794, new_AGEMA_signal_15793, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_16149, new_AGEMA_signal_16148, new_AGEMA_signal_16147, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U943 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, new_AGEMA_signal_15031, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_15630, new_AGEMA_signal_15629, new_AGEMA_signal_15628, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U944 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, new_AGEMA_signal_15025, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, new_AGEMA_signal_15631, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U945 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_15024, new_AGEMA_signal_15023, new_AGEMA_signal_15022, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_15636, new_AGEMA_signal_15635, new_AGEMA_signal_15634, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U946 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .a ({new_AGEMA_signal_15000, new_AGEMA_signal_14999, new_AGEMA_signal_14998, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, new_AGEMA_signal_15637, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U947 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_15771, new_AGEMA_signal_15770, new_AGEMA_signal_15769, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_16152, new_AGEMA_signal_16151, new_AGEMA_signal_16150, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U948 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .a ({new_AGEMA_signal_14934, new_AGEMA_signal_14933, new_AGEMA_signal_14932, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_15642, new_AGEMA_signal_15641, new_AGEMA_signal_15640, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U949 ( .s (new_AGEMA_signal_26144), .b ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .a ({new_AGEMA_signal_15756, new_AGEMA_signal_15755, new_AGEMA_signal_15754, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_16155, new_AGEMA_signal_16154, new_AGEMA_signal_16153, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U950 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_15753, new_AGEMA_signal_15752, new_AGEMA_signal_15751, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_16158, new_AGEMA_signal_16157, new_AGEMA_signal_16156, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U951 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, new_AGEMA_signal_14917, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_15645, new_AGEMA_signal_15644, new_AGEMA_signal_15643, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U952 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_15108, new_AGEMA_signal_15107, new_AGEMA_signal_15106, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_15648, new_AGEMA_signal_15647, new_AGEMA_signal_15646, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U953 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_14916, new_AGEMA_signal_14915, new_AGEMA_signal_14914, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_15651, new_AGEMA_signal_15650, new_AGEMA_signal_15649, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U954 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, new_AGEMA_signal_14911, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_15654, new_AGEMA_signal_15653, new_AGEMA_signal_15652, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U955 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .a ({new_AGEMA_signal_14910, new_AGEMA_signal_14909, new_AGEMA_signal_14908, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, new_AGEMA_signal_15655, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U956 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_15750, new_AGEMA_signal_15749, new_AGEMA_signal_15748, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_16161, new_AGEMA_signal_16160, new_AGEMA_signal_16159, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U957 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .a ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, new_AGEMA_signal_14995, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_15660, new_AGEMA_signal_15659, new_AGEMA_signal_15658, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U958 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .a ({new_AGEMA_signal_15783, new_AGEMA_signal_15782, new_AGEMA_signal_15781, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_16164, new_AGEMA_signal_16163, new_AGEMA_signal_16162, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U959 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_15780, new_AGEMA_signal_15779, new_AGEMA_signal_15778, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_16167, new_AGEMA_signal_16166, new_AGEMA_signal_16165, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U960 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_14988, new_AGEMA_signal_14987, new_AGEMA_signal_14986, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, new_AGEMA_signal_15661, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U961 ( .s (new_AGEMA_signal_26140), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_14985, new_AGEMA_signal_14984, new_AGEMA_signal_14983, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_15666, new_AGEMA_signal_15665, new_AGEMA_signal_15664, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U962 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_14982, new_AGEMA_signal_14981, new_AGEMA_signal_14980, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, new_AGEMA_signal_15667, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U963 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, new_AGEMA_signal_15103, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_15672, new_AGEMA_signal_15671, new_AGEMA_signal_15670, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U964 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .a ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, new_AGEMA_signal_14977, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, new_AGEMA_signal_15673, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U965 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_15777, new_AGEMA_signal_15776, new_AGEMA_signal_15775, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_16170, new_AGEMA_signal_16169, new_AGEMA_signal_16168, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U966 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .a ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, new_AGEMA_signal_14971, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_15678, new_AGEMA_signal_15677, new_AGEMA_signal_15676, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U967 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .a ({new_AGEMA_signal_15774, new_AGEMA_signal_15773, new_AGEMA_signal_15772, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_16173, new_AGEMA_signal_16172, new_AGEMA_signal_16171, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U968 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_15768, new_AGEMA_signal_15767, new_AGEMA_signal_15766, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_16176, new_AGEMA_signal_16175, new_AGEMA_signal_16174, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U969 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, new_AGEMA_signal_14959, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_15681, new_AGEMA_signal_15680, new_AGEMA_signal_15679, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U970 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_14958, new_AGEMA_signal_14957, new_AGEMA_signal_14956, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_15684, new_AGEMA_signal_15683, new_AGEMA_signal_15682, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U971 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, new_AGEMA_signal_14953, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, new_AGEMA_signal_15685, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U972 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .a ({new_AGEMA_signal_14952, new_AGEMA_signal_14951, new_AGEMA_signal_14950, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_15690, new_AGEMA_signal_15689, new_AGEMA_signal_15688, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U973 ( .s (new_AGEMA_signal_26136), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_15765, new_AGEMA_signal_15764, new_AGEMA_signal_15763, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_16179, new_AGEMA_signal_16178, new_AGEMA_signal_16177, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U974 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .a ({new_AGEMA_signal_15102, new_AGEMA_signal_15101, new_AGEMA_signal_15100, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, new_AGEMA_signal_15691, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U975 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .a ({new_AGEMA_signal_14946, new_AGEMA_signal_14945, new_AGEMA_signal_14944, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_15696, new_AGEMA_signal_15695, new_AGEMA_signal_15694, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U976 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .a ({new_AGEMA_signal_15762, new_AGEMA_signal_15761, new_AGEMA_signal_15760, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_16182, new_AGEMA_signal_16181, new_AGEMA_signal_16180, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U977 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, new_AGEMA_signal_15757, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, new_AGEMA_signal_16183, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U978 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_14937, new_AGEMA_signal_14936, new_AGEMA_signal_14935, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, new_AGEMA_signal_15697, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U979 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, new_AGEMA_signal_14929, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_15702, new_AGEMA_signal_15701, new_AGEMA_signal_15700, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U980 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_14928, new_AGEMA_signal_14927, new_AGEMA_signal_14926, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, new_AGEMA_signal_15703, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U981 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .a ({new_AGEMA_signal_14904, new_AGEMA_signal_14903, new_AGEMA_signal_14902, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_15708, new_AGEMA_signal_15707, new_AGEMA_signal_15706, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U982 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_15735, new_AGEMA_signal_15734, new_AGEMA_signal_15733, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_16188, new_AGEMA_signal_16187, new_AGEMA_signal_16186, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U983 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .a ({new_AGEMA_signal_14838, new_AGEMA_signal_14837, new_AGEMA_signal_14836, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, new_AGEMA_signal_15709, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U984 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .a ({new_AGEMA_signal_15720, new_AGEMA_signal_15719, new_AGEMA_signal_15718, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, new_AGEMA_signal_16189, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) U985 ( .s (new_AGEMA_signal_26132), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_15822, new_AGEMA_signal_15821, new_AGEMA_signal_15820, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_16194, new_AGEMA_signal_16193, new_AGEMA_signal_16192, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15474, new_AGEMA_signal_15473, new_AGEMA_signal_15472, RoundOutput[0]}), .a ({new_AGEMA_signal_26172, new_AGEMA_signal_26168, new_AGEMA_signal_26164, new_AGEMA_signal_26160}), .c ({new_AGEMA_signal_16200, new_AGEMA_signal_16199, new_AGEMA_signal_16198, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, new_AGEMA_signal_16093, RoundOutput[1]}), .a ({new_AGEMA_signal_26188, new_AGEMA_signal_26184, new_AGEMA_signal_26180, new_AGEMA_signal_26176}), .c ({new_AGEMA_signal_16722, new_AGEMA_signal_16721, new_AGEMA_signal_16720, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, new_AGEMA_signal_15565, RoundOutput[2]}), .a ({new_AGEMA_signal_26204, new_AGEMA_signal_26200, new_AGEMA_signal_26196, new_AGEMA_signal_26192}), .c ({new_AGEMA_signal_16206, new_AGEMA_signal_16205, new_AGEMA_signal_16204, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, new_AGEMA_signal_16117, RoundOutput[3]}), .a ({new_AGEMA_signal_26220, new_AGEMA_signal_26216, new_AGEMA_signal_26212, new_AGEMA_signal_26208}), .c ({new_AGEMA_signal_16728, new_AGEMA_signal_16727, new_AGEMA_signal_16726, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16134, new_AGEMA_signal_16133, new_AGEMA_signal_16132, RoundOutput[4]}), .a ({new_AGEMA_signal_26236, new_AGEMA_signal_26232, new_AGEMA_signal_26228, new_AGEMA_signal_26224}), .c ({new_AGEMA_signal_16734, new_AGEMA_signal_16733, new_AGEMA_signal_16732, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, new_AGEMA_signal_15625, RoundOutput[5]}), .a ({new_AGEMA_signal_26252, new_AGEMA_signal_26248, new_AGEMA_signal_26244, new_AGEMA_signal_26240}), .c ({new_AGEMA_signal_16212, new_AGEMA_signal_16211, new_AGEMA_signal_16210, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15648, new_AGEMA_signal_15647, new_AGEMA_signal_15646, RoundOutput[6]}), .a ({new_AGEMA_signal_26268, new_AGEMA_signal_26264, new_AGEMA_signal_26260, new_AGEMA_signal_26256}), .c ({new_AGEMA_signal_16218, new_AGEMA_signal_16217, new_AGEMA_signal_16216, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15672, new_AGEMA_signal_15671, new_AGEMA_signal_15670, RoundOutput[7]}), .a ({new_AGEMA_signal_26284, new_AGEMA_signal_26280, new_AGEMA_signal_26276, new_AGEMA_signal_26272}), .c ({new_AGEMA_signal_16224, new_AGEMA_signal_16223, new_AGEMA_signal_16222, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, new_AGEMA_signal_15691, RoundOutput[8]}), .a ({new_AGEMA_signal_26300, new_AGEMA_signal_26296, new_AGEMA_signal_26292, new_AGEMA_signal_26288}), .c ({new_AGEMA_signal_16230, new_AGEMA_signal_16229, new_AGEMA_signal_16228, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16194, new_AGEMA_signal_16193, new_AGEMA_signal_16192, RoundOutput[9]}), .a ({new_AGEMA_signal_26316, new_AGEMA_signal_26312, new_AGEMA_signal_26308, new_AGEMA_signal_26304}), .c ({new_AGEMA_signal_16740, new_AGEMA_signal_16739, new_AGEMA_signal_16738, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, new_AGEMA_signal_15493, RoundOutput[10]}), .a ({new_AGEMA_signal_26332, new_AGEMA_signal_26328, new_AGEMA_signal_26324, new_AGEMA_signal_26320}), .c ({new_AGEMA_signal_16236, new_AGEMA_signal_16235, new_AGEMA_signal_16234, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16074, new_AGEMA_signal_16073, new_AGEMA_signal_16072, RoundOutput[11]}), .a ({new_AGEMA_signal_26348, new_AGEMA_signal_26344, new_AGEMA_signal_26340, new_AGEMA_signal_26336}), .c ({new_AGEMA_signal_16746, new_AGEMA_signal_16745, new_AGEMA_signal_16744, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16086, new_AGEMA_signal_16085, new_AGEMA_signal_16084, RoundOutput[12]}), .a ({new_AGEMA_signal_26364, new_AGEMA_signal_26360, new_AGEMA_signal_26356, new_AGEMA_signal_26352}), .c ({new_AGEMA_signal_16752, new_AGEMA_signal_16751, new_AGEMA_signal_16750, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15534, new_AGEMA_signal_15533, new_AGEMA_signal_15532, RoundOutput[13]}), .a ({new_AGEMA_signal_26380, new_AGEMA_signal_26376, new_AGEMA_signal_26372, new_AGEMA_signal_26368}), .c ({new_AGEMA_signal_16242, new_AGEMA_signal_16241, new_AGEMA_signal_16240, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, new_AGEMA_signal_15535, RoundOutput[14]}), .a ({new_AGEMA_signal_26396, new_AGEMA_signal_26392, new_AGEMA_signal_26388, new_AGEMA_signal_26384}), .c ({new_AGEMA_signal_16248, new_AGEMA_signal_16247, new_AGEMA_signal_16246, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15540, new_AGEMA_signal_15539, new_AGEMA_signal_15538, RoundOutput[15]}), .a ({new_AGEMA_signal_26412, new_AGEMA_signal_26408, new_AGEMA_signal_26404, new_AGEMA_signal_26400}), .c ({new_AGEMA_signal_16254, new_AGEMA_signal_16253, new_AGEMA_signal_16252, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15543, new_AGEMA_signal_15542, new_AGEMA_signal_15541, RoundOutput[16]}), .a ({new_AGEMA_signal_26428, new_AGEMA_signal_26424, new_AGEMA_signal_26420, new_AGEMA_signal_26416}), .c ({new_AGEMA_signal_16260, new_AGEMA_signal_16259, new_AGEMA_signal_16258, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, new_AGEMA_signal_16087, RoundOutput[17]}), .a ({new_AGEMA_signal_26444, new_AGEMA_signal_26440, new_AGEMA_signal_26436, new_AGEMA_signal_26432}), .c ({new_AGEMA_signal_16758, new_AGEMA_signal_16757, new_AGEMA_signal_16756, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15546, new_AGEMA_signal_15545, new_AGEMA_signal_15544, RoundOutput[18]}), .a ({new_AGEMA_signal_26460, new_AGEMA_signal_26456, new_AGEMA_signal_26452, new_AGEMA_signal_26448}), .c ({new_AGEMA_signal_16266, new_AGEMA_signal_16265, new_AGEMA_signal_16264, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16092, new_AGEMA_signal_16091, new_AGEMA_signal_16090, RoundOutput[19]}), .a ({new_AGEMA_signal_26476, new_AGEMA_signal_26472, new_AGEMA_signal_26468, new_AGEMA_signal_26464}), .c ({new_AGEMA_signal_16764, new_AGEMA_signal_16763, new_AGEMA_signal_16762, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16098, new_AGEMA_signal_16097, new_AGEMA_signal_16096, RoundOutput[20]}), .a ({new_AGEMA_signal_26492, new_AGEMA_signal_26488, new_AGEMA_signal_26484, new_AGEMA_signal_26480}), .c ({new_AGEMA_signal_16770, new_AGEMA_signal_16769, new_AGEMA_signal_16768, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, new_AGEMA_signal_15547, RoundOutput[21]}), .a ({new_AGEMA_signal_26508, new_AGEMA_signal_26504, new_AGEMA_signal_26500, new_AGEMA_signal_26496}), .c ({new_AGEMA_signal_16272, new_AGEMA_signal_16271, new_AGEMA_signal_16270, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15552, new_AGEMA_signal_15551, new_AGEMA_signal_15550, RoundOutput[22]}), .a ({new_AGEMA_signal_26524, new_AGEMA_signal_26520, new_AGEMA_signal_26516, new_AGEMA_signal_26512}), .c ({new_AGEMA_signal_16278, new_AGEMA_signal_16277, new_AGEMA_signal_16276, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, new_AGEMA_signal_15553, RoundOutput[23]}), .a ({new_AGEMA_signal_26540, new_AGEMA_signal_26536, new_AGEMA_signal_26532, new_AGEMA_signal_26528}), .c ({new_AGEMA_signal_16284, new_AGEMA_signal_16283, new_AGEMA_signal_16282, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15558, new_AGEMA_signal_15557, new_AGEMA_signal_15556, RoundOutput[24]}), .a ({new_AGEMA_signal_26556, new_AGEMA_signal_26552, new_AGEMA_signal_26548, new_AGEMA_signal_26544}), .c ({new_AGEMA_signal_16290, new_AGEMA_signal_16289, new_AGEMA_signal_16288, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, new_AGEMA_signal_16099, RoundOutput[25]}), .a ({new_AGEMA_signal_26572, new_AGEMA_signal_26568, new_AGEMA_signal_26564, new_AGEMA_signal_26560}), .c ({new_AGEMA_signal_16776, new_AGEMA_signal_16775, new_AGEMA_signal_16774, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, new_AGEMA_signal_15559, RoundOutput[26]}), .a ({new_AGEMA_signal_26588, new_AGEMA_signal_26584, new_AGEMA_signal_26580, new_AGEMA_signal_26576}), .c ({new_AGEMA_signal_16296, new_AGEMA_signal_16295, new_AGEMA_signal_16294, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16104, new_AGEMA_signal_16103, new_AGEMA_signal_16102, RoundOutput[27]}), .a ({new_AGEMA_signal_26604, new_AGEMA_signal_26600, new_AGEMA_signal_26596, new_AGEMA_signal_26592}), .c ({new_AGEMA_signal_16782, new_AGEMA_signal_16781, new_AGEMA_signal_16780, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, new_AGEMA_signal_16105, RoundOutput[28]}), .a ({new_AGEMA_signal_26620, new_AGEMA_signal_26616, new_AGEMA_signal_26612, new_AGEMA_signal_26608}), .c ({new_AGEMA_signal_16788, new_AGEMA_signal_16787, new_AGEMA_signal_16786, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15564, new_AGEMA_signal_15563, new_AGEMA_signal_15562, RoundOutput[29]}), .a ({new_AGEMA_signal_26636, new_AGEMA_signal_26632, new_AGEMA_signal_26628, new_AGEMA_signal_26624}), .c ({new_AGEMA_signal_16302, new_AGEMA_signal_16301, new_AGEMA_signal_16300, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15570, new_AGEMA_signal_15569, new_AGEMA_signal_15568, RoundOutput[30]}), .a ({new_AGEMA_signal_26652, new_AGEMA_signal_26648, new_AGEMA_signal_26644, new_AGEMA_signal_26640}), .c ({new_AGEMA_signal_16308, new_AGEMA_signal_16307, new_AGEMA_signal_16306, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, new_AGEMA_signal_15571, RoundOutput[31]}), .a ({new_AGEMA_signal_26668, new_AGEMA_signal_26664, new_AGEMA_signal_26660, new_AGEMA_signal_26656}), .c ({new_AGEMA_signal_16314, new_AGEMA_signal_16313, new_AGEMA_signal_16312, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15576, new_AGEMA_signal_15575, new_AGEMA_signal_15574, RoundOutput[32]}), .a ({new_AGEMA_signal_26684, new_AGEMA_signal_26680, new_AGEMA_signal_26676, new_AGEMA_signal_26672}), .c ({new_AGEMA_signal_16320, new_AGEMA_signal_16319, new_AGEMA_signal_16318, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16110, new_AGEMA_signal_16109, new_AGEMA_signal_16108, RoundOutput[33]}), .a ({new_AGEMA_signal_26700, new_AGEMA_signal_26696, new_AGEMA_signal_26692, new_AGEMA_signal_26688}), .c ({new_AGEMA_signal_16794, new_AGEMA_signal_16793, new_AGEMA_signal_16792, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, new_AGEMA_signal_15577, RoundOutput[34]}), .a ({new_AGEMA_signal_26716, new_AGEMA_signal_26712, new_AGEMA_signal_26708, new_AGEMA_signal_26704}), .c ({new_AGEMA_signal_16326, new_AGEMA_signal_16325, new_AGEMA_signal_16324, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16113, new_AGEMA_signal_16112, new_AGEMA_signal_16111, RoundOutput[35]}), .a ({new_AGEMA_signal_26732, new_AGEMA_signal_26728, new_AGEMA_signal_26724, new_AGEMA_signal_26720}), .c ({new_AGEMA_signal_16800, new_AGEMA_signal_16799, new_AGEMA_signal_16798, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16116, new_AGEMA_signal_16115, new_AGEMA_signal_16114, RoundOutput[36]}), .a ({new_AGEMA_signal_26748, new_AGEMA_signal_26744, new_AGEMA_signal_26740, new_AGEMA_signal_26736}), .c ({new_AGEMA_signal_16806, new_AGEMA_signal_16805, new_AGEMA_signal_16804, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15582, new_AGEMA_signal_15581, new_AGEMA_signal_15580, RoundOutput[37]}), .a ({new_AGEMA_signal_26764, new_AGEMA_signal_26760, new_AGEMA_signal_26756, new_AGEMA_signal_26752}), .c ({new_AGEMA_signal_16332, new_AGEMA_signal_16331, new_AGEMA_signal_16330, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, new_AGEMA_signal_15583, RoundOutput[38]}), .a ({new_AGEMA_signal_26780, new_AGEMA_signal_26776, new_AGEMA_signal_26772, new_AGEMA_signal_26768}), .c ({new_AGEMA_signal_16338, new_AGEMA_signal_16337, new_AGEMA_signal_16336, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15588, new_AGEMA_signal_15587, new_AGEMA_signal_15586, RoundOutput[39]}), .a ({new_AGEMA_signal_26796, new_AGEMA_signal_26792, new_AGEMA_signal_26788, new_AGEMA_signal_26784}), .c ({new_AGEMA_signal_16344, new_AGEMA_signal_16343, new_AGEMA_signal_16342, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15591, new_AGEMA_signal_15590, new_AGEMA_signal_15589, RoundOutput[40]}), .a ({new_AGEMA_signal_26812, new_AGEMA_signal_26808, new_AGEMA_signal_26804, new_AGEMA_signal_26800}), .c ({new_AGEMA_signal_16350, new_AGEMA_signal_16349, new_AGEMA_signal_16348, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16122, new_AGEMA_signal_16121, new_AGEMA_signal_16120, RoundOutput[41]}), .a ({new_AGEMA_signal_26828, new_AGEMA_signal_26824, new_AGEMA_signal_26820, new_AGEMA_signal_26816}), .c ({new_AGEMA_signal_16812, new_AGEMA_signal_16811, new_AGEMA_signal_16810, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15594, new_AGEMA_signal_15593, new_AGEMA_signal_15592, RoundOutput[42]}), .a ({new_AGEMA_signal_26844, new_AGEMA_signal_26840, new_AGEMA_signal_26836, new_AGEMA_signal_26832}), .c ({new_AGEMA_signal_16356, new_AGEMA_signal_16355, new_AGEMA_signal_16354, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16125, new_AGEMA_signal_16124, new_AGEMA_signal_16123, RoundOutput[43]}), .a ({new_AGEMA_signal_26860, new_AGEMA_signal_26856, new_AGEMA_signal_26852, new_AGEMA_signal_26848}), .c ({new_AGEMA_signal_16818, new_AGEMA_signal_16817, new_AGEMA_signal_16816, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16128, new_AGEMA_signal_16127, new_AGEMA_signal_16126, RoundOutput[44]}), .a ({new_AGEMA_signal_26876, new_AGEMA_signal_26872, new_AGEMA_signal_26868, new_AGEMA_signal_26864}), .c ({new_AGEMA_signal_16824, new_AGEMA_signal_16823, new_AGEMA_signal_16822, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15597, new_AGEMA_signal_15596, new_AGEMA_signal_15595, RoundOutput[45]}), .a ({new_AGEMA_signal_26892, new_AGEMA_signal_26888, new_AGEMA_signal_26884, new_AGEMA_signal_26880}), .c ({new_AGEMA_signal_16362, new_AGEMA_signal_16361, new_AGEMA_signal_16360, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15600, new_AGEMA_signal_15599, new_AGEMA_signal_15598, RoundOutput[46]}), .a ({new_AGEMA_signal_26908, new_AGEMA_signal_26904, new_AGEMA_signal_26900, new_AGEMA_signal_26896}), .c ({new_AGEMA_signal_16368, new_AGEMA_signal_16367, new_AGEMA_signal_16366, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, new_AGEMA_signal_15601, RoundOutput[47]}), .a ({new_AGEMA_signal_26924, new_AGEMA_signal_26920, new_AGEMA_signal_26916, new_AGEMA_signal_26912}), .c ({new_AGEMA_signal_16374, new_AGEMA_signal_16373, new_AGEMA_signal_16372, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15606, new_AGEMA_signal_15605, new_AGEMA_signal_15604, RoundOutput[48]}), .a ({new_AGEMA_signal_26940, new_AGEMA_signal_26936, new_AGEMA_signal_26932, new_AGEMA_signal_26928}), .c ({new_AGEMA_signal_16380, new_AGEMA_signal_16379, new_AGEMA_signal_16378, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16131, new_AGEMA_signal_16130, new_AGEMA_signal_16129, RoundOutput[49]}), .a ({new_AGEMA_signal_26956, new_AGEMA_signal_26952, new_AGEMA_signal_26948, new_AGEMA_signal_26944}), .c ({new_AGEMA_signal_16830, new_AGEMA_signal_16829, new_AGEMA_signal_16828, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, new_AGEMA_signal_15607, RoundOutput[50]}), .a ({new_AGEMA_signal_26972, new_AGEMA_signal_26968, new_AGEMA_signal_26964, new_AGEMA_signal_26960}), .c ({new_AGEMA_signal_16386, new_AGEMA_signal_16385, new_AGEMA_signal_16384, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, new_AGEMA_signal_16135, RoundOutput[51]}), .a ({new_AGEMA_signal_26988, new_AGEMA_signal_26984, new_AGEMA_signal_26980, new_AGEMA_signal_26976}), .c ({new_AGEMA_signal_16836, new_AGEMA_signal_16835, new_AGEMA_signal_16834, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16140, new_AGEMA_signal_16139, new_AGEMA_signal_16138, RoundOutput[52]}), .a ({new_AGEMA_signal_27004, new_AGEMA_signal_27000, new_AGEMA_signal_26996, new_AGEMA_signal_26992}), .c ({new_AGEMA_signal_16842, new_AGEMA_signal_16841, new_AGEMA_signal_16840, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15612, new_AGEMA_signal_15611, new_AGEMA_signal_15610, RoundOutput[53]}), .a ({new_AGEMA_signal_27020, new_AGEMA_signal_27016, new_AGEMA_signal_27012, new_AGEMA_signal_27008}), .c ({new_AGEMA_signal_16392, new_AGEMA_signal_16391, new_AGEMA_signal_16390, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15615, new_AGEMA_signal_15614, new_AGEMA_signal_15613, RoundOutput[54]}), .a ({new_AGEMA_signal_27036, new_AGEMA_signal_27032, new_AGEMA_signal_27028, new_AGEMA_signal_27024}), .c ({new_AGEMA_signal_16398, new_AGEMA_signal_16397, new_AGEMA_signal_16396, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15618, new_AGEMA_signal_15617, new_AGEMA_signal_15616, RoundOutput[55]}), .a ({new_AGEMA_signal_27052, new_AGEMA_signal_27048, new_AGEMA_signal_27044, new_AGEMA_signal_27040}), .c ({new_AGEMA_signal_16404, new_AGEMA_signal_16403, new_AGEMA_signal_16402, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, new_AGEMA_signal_15619, RoundOutput[56]}), .a ({new_AGEMA_signal_27068, new_AGEMA_signal_27064, new_AGEMA_signal_27060, new_AGEMA_signal_27056}), .c ({new_AGEMA_signal_16410, new_AGEMA_signal_16409, new_AGEMA_signal_16408, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16143, new_AGEMA_signal_16142, new_AGEMA_signal_16141, RoundOutput[57]}), .a ({new_AGEMA_signal_27084, new_AGEMA_signal_27080, new_AGEMA_signal_27076, new_AGEMA_signal_27072}), .c ({new_AGEMA_signal_16848, new_AGEMA_signal_16847, new_AGEMA_signal_16846, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15624, new_AGEMA_signal_15623, new_AGEMA_signal_15622, RoundOutput[58]}), .a ({new_AGEMA_signal_27100, new_AGEMA_signal_27096, new_AGEMA_signal_27092, new_AGEMA_signal_27088}), .c ({new_AGEMA_signal_16416, new_AGEMA_signal_16415, new_AGEMA_signal_16414, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16146, new_AGEMA_signal_16145, new_AGEMA_signal_16144, RoundOutput[59]}), .a ({new_AGEMA_signal_27116, new_AGEMA_signal_27112, new_AGEMA_signal_27108, new_AGEMA_signal_27104}), .c ({new_AGEMA_signal_16854, new_AGEMA_signal_16853, new_AGEMA_signal_16852, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16149, new_AGEMA_signal_16148, new_AGEMA_signal_16147, RoundOutput[60]}), .a ({new_AGEMA_signal_27132, new_AGEMA_signal_27128, new_AGEMA_signal_27124, new_AGEMA_signal_27120}), .c ({new_AGEMA_signal_16860, new_AGEMA_signal_16859, new_AGEMA_signal_16858, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15630, new_AGEMA_signal_15629, new_AGEMA_signal_15628, RoundOutput[61]}), .a ({new_AGEMA_signal_27148, new_AGEMA_signal_27144, new_AGEMA_signal_27140, new_AGEMA_signal_27136}), .c ({new_AGEMA_signal_16422, new_AGEMA_signal_16421, new_AGEMA_signal_16420, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, new_AGEMA_signal_15631, RoundOutput[62]}), .a ({new_AGEMA_signal_27164, new_AGEMA_signal_27160, new_AGEMA_signal_27156, new_AGEMA_signal_27152}), .c ({new_AGEMA_signal_16428, new_AGEMA_signal_16427, new_AGEMA_signal_16426, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15636, new_AGEMA_signal_15635, new_AGEMA_signal_15634, RoundOutput[63]}), .a ({new_AGEMA_signal_27180, new_AGEMA_signal_27176, new_AGEMA_signal_27172, new_AGEMA_signal_27168}), .c ({new_AGEMA_signal_16434, new_AGEMA_signal_16433, new_AGEMA_signal_16432, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, new_AGEMA_signal_15637, RoundOutput[64]}), .a ({new_AGEMA_signal_27196, new_AGEMA_signal_27192, new_AGEMA_signal_27188, new_AGEMA_signal_27184}), .c ({new_AGEMA_signal_16440, new_AGEMA_signal_16439, new_AGEMA_signal_16438, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16152, new_AGEMA_signal_16151, new_AGEMA_signal_16150, RoundOutput[65]}), .a ({new_AGEMA_signal_27212, new_AGEMA_signal_27208, new_AGEMA_signal_27204, new_AGEMA_signal_27200}), .c ({new_AGEMA_signal_16866, new_AGEMA_signal_16865, new_AGEMA_signal_16864, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15642, new_AGEMA_signal_15641, new_AGEMA_signal_15640, RoundOutput[66]}), .a ({new_AGEMA_signal_27228, new_AGEMA_signal_27224, new_AGEMA_signal_27220, new_AGEMA_signal_27216}), .c ({new_AGEMA_signal_16446, new_AGEMA_signal_16445, new_AGEMA_signal_16444, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16155, new_AGEMA_signal_16154, new_AGEMA_signal_16153, RoundOutput[67]}), .a ({new_AGEMA_signal_27244, new_AGEMA_signal_27240, new_AGEMA_signal_27236, new_AGEMA_signal_27232}), .c ({new_AGEMA_signal_16872, new_AGEMA_signal_16871, new_AGEMA_signal_16870, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16158, new_AGEMA_signal_16157, new_AGEMA_signal_16156, RoundOutput[68]}), .a ({new_AGEMA_signal_27260, new_AGEMA_signal_27256, new_AGEMA_signal_27252, new_AGEMA_signal_27248}), .c ({new_AGEMA_signal_16878, new_AGEMA_signal_16877, new_AGEMA_signal_16876, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15645, new_AGEMA_signal_15644, new_AGEMA_signal_15643, RoundOutput[69]}), .a ({new_AGEMA_signal_27276, new_AGEMA_signal_27272, new_AGEMA_signal_27268, new_AGEMA_signal_27264}), .c ({new_AGEMA_signal_16452, new_AGEMA_signal_16451, new_AGEMA_signal_16450, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15651, new_AGEMA_signal_15650, new_AGEMA_signal_15649, RoundOutput[70]}), .a ({new_AGEMA_signal_27292, new_AGEMA_signal_27288, new_AGEMA_signal_27284, new_AGEMA_signal_27280}), .c ({new_AGEMA_signal_16458, new_AGEMA_signal_16457, new_AGEMA_signal_16456, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15654, new_AGEMA_signal_15653, new_AGEMA_signal_15652, RoundOutput[71]}), .a ({new_AGEMA_signal_27308, new_AGEMA_signal_27304, new_AGEMA_signal_27300, new_AGEMA_signal_27296}), .c ({new_AGEMA_signal_16464, new_AGEMA_signal_16463, new_AGEMA_signal_16462, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, new_AGEMA_signal_15655, RoundOutput[72]}), .a ({new_AGEMA_signal_27324, new_AGEMA_signal_27320, new_AGEMA_signal_27316, new_AGEMA_signal_27312}), .c ({new_AGEMA_signal_16470, new_AGEMA_signal_16469, new_AGEMA_signal_16468, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16161, new_AGEMA_signal_16160, new_AGEMA_signal_16159, RoundOutput[73]}), .a ({new_AGEMA_signal_27340, new_AGEMA_signal_27336, new_AGEMA_signal_27332, new_AGEMA_signal_27328}), .c ({new_AGEMA_signal_16884, new_AGEMA_signal_16883, new_AGEMA_signal_16882, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15660, new_AGEMA_signal_15659, new_AGEMA_signal_15658, RoundOutput[74]}), .a ({new_AGEMA_signal_27356, new_AGEMA_signal_27352, new_AGEMA_signal_27348, new_AGEMA_signal_27344}), .c ({new_AGEMA_signal_16476, new_AGEMA_signal_16475, new_AGEMA_signal_16474, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16164, new_AGEMA_signal_16163, new_AGEMA_signal_16162, RoundOutput[75]}), .a ({new_AGEMA_signal_27372, new_AGEMA_signal_27368, new_AGEMA_signal_27364, new_AGEMA_signal_27360}), .c ({new_AGEMA_signal_16890, new_AGEMA_signal_16889, new_AGEMA_signal_16888, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16167, new_AGEMA_signal_16166, new_AGEMA_signal_16165, RoundOutput[76]}), .a ({new_AGEMA_signal_27388, new_AGEMA_signal_27384, new_AGEMA_signal_27380, new_AGEMA_signal_27376}), .c ({new_AGEMA_signal_16896, new_AGEMA_signal_16895, new_AGEMA_signal_16894, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, new_AGEMA_signal_15661, RoundOutput[77]}), .a ({new_AGEMA_signal_27404, new_AGEMA_signal_27400, new_AGEMA_signal_27396, new_AGEMA_signal_27392}), .c ({new_AGEMA_signal_16482, new_AGEMA_signal_16481, new_AGEMA_signal_16480, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15666, new_AGEMA_signal_15665, new_AGEMA_signal_15664, RoundOutput[78]}), .a ({new_AGEMA_signal_27420, new_AGEMA_signal_27416, new_AGEMA_signal_27412, new_AGEMA_signal_27408}), .c ({new_AGEMA_signal_16488, new_AGEMA_signal_16487, new_AGEMA_signal_16486, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, new_AGEMA_signal_15667, RoundOutput[79]}), .a ({new_AGEMA_signal_27436, new_AGEMA_signal_27432, new_AGEMA_signal_27428, new_AGEMA_signal_27424}), .c ({new_AGEMA_signal_16494, new_AGEMA_signal_16493, new_AGEMA_signal_16492, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, new_AGEMA_signal_15673, RoundOutput[80]}), .a ({new_AGEMA_signal_27452, new_AGEMA_signal_27448, new_AGEMA_signal_27444, new_AGEMA_signal_27440}), .c ({new_AGEMA_signal_16500, new_AGEMA_signal_16499, new_AGEMA_signal_16498, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16170, new_AGEMA_signal_16169, new_AGEMA_signal_16168, RoundOutput[81]}), .a ({new_AGEMA_signal_27468, new_AGEMA_signal_27464, new_AGEMA_signal_27460, new_AGEMA_signal_27456}), .c ({new_AGEMA_signal_16902, new_AGEMA_signal_16901, new_AGEMA_signal_16900, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15678, new_AGEMA_signal_15677, new_AGEMA_signal_15676, RoundOutput[82]}), .a ({new_AGEMA_signal_27484, new_AGEMA_signal_27480, new_AGEMA_signal_27476, new_AGEMA_signal_27472}), .c ({new_AGEMA_signal_16506, new_AGEMA_signal_16505, new_AGEMA_signal_16504, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16173, new_AGEMA_signal_16172, new_AGEMA_signal_16171, RoundOutput[83]}), .a ({new_AGEMA_signal_27500, new_AGEMA_signal_27496, new_AGEMA_signal_27492, new_AGEMA_signal_27488}), .c ({new_AGEMA_signal_16908, new_AGEMA_signal_16907, new_AGEMA_signal_16906, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16176, new_AGEMA_signal_16175, new_AGEMA_signal_16174, RoundOutput[84]}), .a ({new_AGEMA_signal_27516, new_AGEMA_signal_27512, new_AGEMA_signal_27508, new_AGEMA_signal_27504}), .c ({new_AGEMA_signal_16914, new_AGEMA_signal_16913, new_AGEMA_signal_16912, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15681, new_AGEMA_signal_15680, new_AGEMA_signal_15679, RoundOutput[85]}), .a ({new_AGEMA_signal_27532, new_AGEMA_signal_27528, new_AGEMA_signal_27524, new_AGEMA_signal_27520}), .c ({new_AGEMA_signal_16512, new_AGEMA_signal_16511, new_AGEMA_signal_16510, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15684, new_AGEMA_signal_15683, new_AGEMA_signal_15682, RoundOutput[86]}), .a ({new_AGEMA_signal_27548, new_AGEMA_signal_27544, new_AGEMA_signal_27540, new_AGEMA_signal_27536}), .c ({new_AGEMA_signal_16518, new_AGEMA_signal_16517, new_AGEMA_signal_16516, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, new_AGEMA_signal_15685, RoundOutput[87]}), .a ({new_AGEMA_signal_27564, new_AGEMA_signal_27560, new_AGEMA_signal_27556, new_AGEMA_signal_27552}), .c ({new_AGEMA_signal_16524, new_AGEMA_signal_16523, new_AGEMA_signal_16522, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15690, new_AGEMA_signal_15689, new_AGEMA_signal_15688, RoundOutput[88]}), .a ({new_AGEMA_signal_27580, new_AGEMA_signal_27576, new_AGEMA_signal_27572, new_AGEMA_signal_27568}), .c ({new_AGEMA_signal_16530, new_AGEMA_signal_16529, new_AGEMA_signal_16528, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16179, new_AGEMA_signal_16178, new_AGEMA_signal_16177, RoundOutput[89]}), .a ({new_AGEMA_signal_27596, new_AGEMA_signal_27592, new_AGEMA_signal_27588, new_AGEMA_signal_27584}), .c ({new_AGEMA_signal_16920, new_AGEMA_signal_16919, new_AGEMA_signal_16918, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15696, new_AGEMA_signal_15695, new_AGEMA_signal_15694, RoundOutput[90]}), .a ({new_AGEMA_signal_27612, new_AGEMA_signal_27608, new_AGEMA_signal_27604, new_AGEMA_signal_27600}), .c ({new_AGEMA_signal_16536, new_AGEMA_signal_16535, new_AGEMA_signal_16534, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16182, new_AGEMA_signal_16181, new_AGEMA_signal_16180, RoundOutput[91]}), .a ({new_AGEMA_signal_27628, new_AGEMA_signal_27624, new_AGEMA_signal_27620, new_AGEMA_signal_27616}), .c ({new_AGEMA_signal_16926, new_AGEMA_signal_16925, new_AGEMA_signal_16924, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, new_AGEMA_signal_16183, RoundOutput[92]}), .a ({new_AGEMA_signal_27644, new_AGEMA_signal_27640, new_AGEMA_signal_27636, new_AGEMA_signal_27632}), .c ({new_AGEMA_signal_16932, new_AGEMA_signal_16931, new_AGEMA_signal_16930, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, new_AGEMA_signal_15697, RoundOutput[93]}), .a ({new_AGEMA_signal_27660, new_AGEMA_signal_27656, new_AGEMA_signal_27652, new_AGEMA_signal_27648}), .c ({new_AGEMA_signal_16542, new_AGEMA_signal_16541, new_AGEMA_signal_16540, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15702, new_AGEMA_signal_15701, new_AGEMA_signal_15700, RoundOutput[94]}), .a ({new_AGEMA_signal_27676, new_AGEMA_signal_27672, new_AGEMA_signal_27668, new_AGEMA_signal_27664}), .c ({new_AGEMA_signal_16548, new_AGEMA_signal_16547, new_AGEMA_signal_16546, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, new_AGEMA_signal_15703, RoundOutput[95]}), .a ({new_AGEMA_signal_27692, new_AGEMA_signal_27688, new_AGEMA_signal_27684, new_AGEMA_signal_27680}), .c ({new_AGEMA_signal_16554, new_AGEMA_signal_16553, new_AGEMA_signal_16552, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15708, new_AGEMA_signal_15707, new_AGEMA_signal_15706, RoundOutput[96]}), .a ({new_AGEMA_signal_27708, new_AGEMA_signal_27704, new_AGEMA_signal_27700, new_AGEMA_signal_27696}), .c ({new_AGEMA_signal_16560, new_AGEMA_signal_16559, new_AGEMA_signal_16558, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16188, new_AGEMA_signal_16187, new_AGEMA_signal_16186, RoundOutput[97]}), .a ({new_AGEMA_signal_27724, new_AGEMA_signal_27720, new_AGEMA_signal_27716, new_AGEMA_signal_27712}), .c ({new_AGEMA_signal_16938, new_AGEMA_signal_16937, new_AGEMA_signal_16936, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, new_AGEMA_signal_15709, RoundOutput[98]}), .a ({new_AGEMA_signal_27740, new_AGEMA_signal_27736, new_AGEMA_signal_27732, new_AGEMA_signal_27728}), .c ({new_AGEMA_signal_16566, new_AGEMA_signal_16565, new_AGEMA_signal_16564, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, new_AGEMA_signal_16189, RoundOutput[99]}), .a ({new_AGEMA_signal_27756, new_AGEMA_signal_27752, new_AGEMA_signal_27748, new_AGEMA_signal_27744}), .c ({new_AGEMA_signal_16944, new_AGEMA_signal_16943, new_AGEMA_signal_16942, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16053, new_AGEMA_signal_16052, new_AGEMA_signal_16051, RoundOutput[100]}), .a ({new_AGEMA_signal_27772, new_AGEMA_signal_27768, new_AGEMA_signal_27764, new_AGEMA_signal_27760}), .c ({new_AGEMA_signal_16950, new_AGEMA_signal_16949, new_AGEMA_signal_16948, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15477, new_AGEMA_signal_15476, new_AGEMA_signal_15475, RoundOutput[101]}), .a ({new_AGEMA_signal_27788, new_AGEMA_signal_27784, new_AGEMA_signal_27780, new_AGEMA_signal_27776}), .c ({new_AGEMA_signal_16572, new_AGEMA_signal_16571, new_AGEMA_signal_16570, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15480, new_AGEMA_signal_15479, new_AGEMA_signal_15478, RoundOutput[102]}), .a ({new_AGEMA_signal_27804, new_AGEMA_signal_27800, new_AGEMA_signal_27796, new_AGEMA_signal_27792}), .c ({new_AGEMA_signal_16578, new_AGEMA_signal_16577, new_AGEMA_signal_16576, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15483, new_AGEMA_signal_15482, new_AGEMA_signal_15481, RoundOutput[103]}), .a ({new_AGEMA_signal_27820, new_AGEMA_signal_27816, new_AGEMA_signal_27812, new_AGEMA_signal_27808}), .c ({new_AGEMA_signal_16584, new_AGEMA_signal_16583, new_AGEMA_signal_16582, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15486, new_AGEMA_signal_15485, new_AGEMA_signal_15484, RoundOutput[104]}), .a ({new_AGEMA_signal_27836, new_AGEMA_signal_27832, new_AGEMA_signal_27828, new_AGEMA_signal_27824}), .c ({new_AGEMA_signal_16590, new_AGEMA_signal_16589, new_AGEMA_signal_16588, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16056, new_AGEMA_signal_16055, new_AGEMA_signal_16054, RoundOutput[105]}), .a ({new_AGEMA_signal_27852, new_AGEMA_signal_27848, new_AGEMA_signal_27844, new_AGEMA_signal_27840}), .c ({new_AGEMA_signal_16956, new_AGEMA_signal_16955, new_AGEMA_signal_16954, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, new_AGEMA_signal_15487, RoundOutput[106]}), .a ({new_AGEMA_signal_27868, new_AGEMA_signal_27864, new_AGEMA_signal_27860, new_AGEMA_signal_27856}), .c ({new_AGEMA_signal_16596, new_AGEMA_signal_16595, new_AGEMA_signal_16594, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, new_AGEMA_signal_16057, RoundOutput[107]}), .a ({new_AGEMA_signal_27884, new_AGEMA_signal_27880, new_AGEMA_signal_27876, new_AGEMA_signal_27872}), .c ({new_AGEMA_signal_16962, new_AGEMA_signal_16961, new_AGEMA_signal_16960, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16062, new_AGEMA_signal_16061, new_AGEMA_signal_16060, RoundOutput[108]}), .a ({new_AGEMA_signal_27900, new_AGEMA_signal_27896, new_AGEMA_signal_27892, new_AGEMA_signal_27888}), .c ({new_AGEMA_signal_16968, new_AGEMA_signal_16967, new_AGEMA_signal_16966, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15492, new_AGEMA_signal_15491, new_AGEMA_signal_15490, RoundOutput[109]}), .a ({new_AGEMA_signal_27916, new_AGEMA_signal_27912, new_AGEMA_signal_27908, new_AGEMA_signal_27904}), .c ({new_AGEMA_signal_16602, new_AGEMA_signal_16601, new_AGEMA_signal_16600, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15498, new_AGEMA_signal_15497, new_AGEMA_signal_15496, RoundOutput[110]}), .a ({new_AGEMA_signal_27932, new_AGEMA_signal_27928, new_AGEMA_signal_27924, new_AGEMA_signal_27920}), .c ({new_AGEMA_signal_16608, new_AGEMA_signal_16607, new_AGEMA_signal_16606, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, new_AGEMA_signal_15499, RoundOutput[111]}), .a ({new_AGEMA_signal_27948, new_AGEMA_signal_27944, new_AGEMA_signal_27940, new_AGEMA_signal_27936}), .c ({new_AGEMA_signal_16614, new_AGEMA_signal_16613, new_AGEMA_signal_16612, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15504, new_AGEMA_signal_15503, new_AGEMA_signal_15502, RoundOutput[112]}), .a ({new_AGEMA_signal_27964, new_AGEMA_signal_27960, new_AGEMA_signal_27956, new_AGEMA_signal_27952}), .c ({new_AGEMA_signal_16620, new_AGEMA_signal_16619, new_AGEMA_signal_16618, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, new_AGEMA_signal_16063, RoundOutput[113]}), .a ({new_AGEMA_signal_27980, new_AGEMA_signal_27976, new_AGEMA_signal_27972, new_AGEMA_signal_27968}), .c ({new_AGEMA_signal_16974, new_AGEMA_signal_16973, new_AGEMA_signal_16972, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15507, new_AGEMA_signal_15506, new_AGEMA_signal_15505, RoundOutput[114]}), .a ({new_AGEMA_signal_27996, new_AGEMA_signal_27992, new_AGEMA_signal_27988, new_AGEMA_signal_27984}), .c ({new_AGEMA_signal_16626, new_AGEMA_signal_16625, new_AGEMA_signal_16624, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16068, new_AGEMA_signal_16067, new_AGEMA_signal_16066, RoundOutput[115]}), .a ({new_AGEMA_signal_28012, new_AGEMA_signal_28008, new_AGEMA_signal_28004, new_AGEMA_signal_28000}), .c ({new_AGEMA_signal_16980, new_AGEMA_signal_16979, new_AGEMA_signal_16978, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, new_AGEMA_signal_16069, RoundOutput[116]}), .a ({new_AGEMA_signal_28028, new_AGEMA_signal_28024, new_AGEMA_signal_28020, new_AGEMA_signal_28016}), .c ({new_AGEMA_signal_16986, new_AGEMA_signal_16985, new_AGEMA_signal_16984, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15510, new_AGEMA_signal_15509, new_AGEMA_signal_15508, RoundOutput[117]}), .a ({new_AGEMA_signal_28044, new_AGEMA_signal_28040, new_AGEMA_signal_28036, new_AGEMA_signal_28032}), .c ({new_AGEMA_signal_16632, new_AGEMA_signal_16631, new_AGEMA_signal_16630, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15513, new_AGEMA_signal_15512, new_AGEMA_signal_15511, RoundOutput[118]}), .a ({new_AGEMA_signal_28060, new_AGEMA_signal_28056, new_AGEMA_signal_28052, new_AGEMA_signal_28048}), .c ({new_AGEMA_signal_16638, new_AGEMA_signal_16637, new_AGEMA_signal_16636, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15516, new_AGEMA_signal_15515, new_AGEMA_signal_15514, RoundOutput[119]}), .a ({new_AGEMA_signal_28076, new_AGEMA_signal_28072, new_AGEMA_signal_28068, new_AGEMA_signal_28064}), .c ({new_AGEMA_signal_16644, new_AGEMA_signal_16643, new_AGEMA_signal_16642, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, new_AGEMA_signal_15517, RoundOutput[120]}), .a ({new_AGEMA_signal_28092, new_AGEMA_signal_28088, new_AGEMA_signal_28084, new_AGEMA_signal_28080}), .c ({new_AGEMA_signal_16650, new_AGEMA_signal_16649, new_AGEMA_signal_16648, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16077, new_AGEMA_signal_16076, new_AGEMA_signal_16075, RoundOutput[121]}), .a ({new_AGEMA_signal_28108, new_AGEMA_signal_28104, new_AGEMA_signal_28100, new_AGEMA_signal_28096}), .c ({new_AGEMA_signal_16992, new_AGEMA_signal_16991, new_AGEMA_signal_16990, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15522, new_AGEMA_signal_15521, new_AGEMA_signal_15520, RoundOutput[122]}), .a ({new_AGEMA_signal_28124, new_AGEMA_signal_28120, new_AGEMA_signal_28116, new_AGEMA_signal_28112}), .c ({new_AGEMA_signal_16656, new_AGEMA_signal_16655, new_AGEMA_signal_16654, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16080, new_AGEMA_signal_16079, new_AGEMA_signal_16078, RoundOutput[123]}), .a ({new_AGEMA_signal_28140, new_AGEMA_signal_28136, new_AGEMA_signal_28132, new_AGEMA_signal_28128}), .c ({new_AGEMA_signal_16998, new_AGEMA_signal_16997, new_AGEMA_signal_16996, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, new_AGEMA_signal_16081, RoundOutput[124]}), .a ({new_AGEMA_signal_28156, new_AGEMA_signal_28152, new_AGEMA_signal_28148, new_AGEMA_signal_28144}), .c ({new_AGEMA_signal_17004, new_AGEMA_signal_17003, new_AGEMA_signal_17002, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, new_AGEMA_signal_15523, RoundOutput[125]}), .a ({new_AGEMA_signal_28172, new_AGEMA_signal_28168, new_AGEMA_signal_28164, new_AGEMA_signal_28160}), .c ({new_AGEMA_signal_16662, new_AGEMA_signal_16661, new_AGEMA_signal_16660, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15528, new_AGEMA_signal_15527, new_AGEMA_signal_15526, RoundOutput[126]}), .a ({new_AGEMA_signal_28188, new_AGEMA_signal_28184, new_AGEMA_signal_28180, new_AGEMA_signal_28176}), .c ({new_AGEMA_signal_16668, new_AGEMA_signal_16667, new_AGEMA_signal_16666, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, new_AGEMA_signal_15529, RoundOutput[127]}), .a ({new_AGEMA_signal_28204, new_AGEMA_signal_28200, new_AGEMA_signal_28196, new_AGEMA_signal_28192}), .c ({new_AGEMA_signal_16674, new_AGEMA_signal_16673, new_AGEMA_signal_16672, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_28216, new_AGEMA_signal_28213, new_AGEMA_signal_28210, new_AGEMA_signal_28207}), .clk (clk), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_28228, new_AGEMA_signal_28225, new_AGEMA_signal_28222, new_AGEMA_signal_28219}), .clk (clk), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_28240, new_AGEMA_signal_28237, new_AGEMA_signal_28234, new_AGEMA_signal_28231}), .clk (clk), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870], Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_28252, new_AGEMA_signal_28249, new_AGEMA_signal_28246, new_AGEMA_signal_28243}), .clk (clk), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, new_AGEMA_signal_10591, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_28264, new_AGEMA_signal_28261, new_AGEMA_signal_28258, new_AGEMA_signal_28255}), .clk (clk), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_28276, new_AGEMA_signal_28273, new_AGEMA_signal_28270, new_AGEMA_signal_28267}), .clk (clk), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_28288, new_AGEMA_signal_28285, new_AGEMA_signal_28282, new_AGEMA_signal_28279}), .clk (clk), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_28300, new_AGEMA_signal_28297, new_AGEMA_signal_28294, new_AGEMA_signal_28291}), .clk (clk), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930], Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_28312, new_AGEMA_signal_28309, new_AGEMA_signal_28306, new_AGEMA_signal_28303}), .clk (clk), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, new_AGEMA_signal_10597, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_28324, new_AGEMA_signal_28321, new_AGEMA_signal_28318, new_AGEMA_signal_28315}), .clk (clk), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_28336, new_AGEMA_signal_28333, new_AGEMA_signal_28330, new_AGEMA_signal_28327}), .clk (clk), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_28348, new_AGEMA_signal_28345, new_AGEMA_signal_28342, new_AGEMA_signal_28339}), .clk (clk), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, new_AGEMA_signal_9892, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_28360, new_AGEMA_signal_28357, new_AGEMA_signal_28354, new_AGEMA_signal_28351}), .clk (clk), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990], Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_28372, new_AGEMA_signal_28369, new_AGEMA_signal_28366, new_AGEMA_signal_28363}), .clk (clk), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_28384, new_AGEMA_signal_28381, new_AGEMA_signal_28378, new_AGEMA_signal_28375}), .clk (clk), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, new_AGEMA_signal_9898, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_28396, new_AGEMA_signal_28393, new_AGEMA_signal_28390, new_AGEMA_signal_28387}), .clk (clk), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_28408, new_AGEMA_signal_28405, new_AGEMA_signal_28402, new_AGEMA_signal_28399}), .clk (clk), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_28420, new_AGEMA_signal_28417, new_AGEMA_signal_28414, new_AGEMA_signal_28411}), .clk (clk), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050], Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, new_AGEMA_signal_10609, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, new_AGEMA_signal_10597, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, new_AGEMA_signal_10591, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11298, new_AGEMA_signal_11297, new_AGEMA_signal_11296, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_11298, new_AGEMA_signal_11297, new_AGEMA_signal_11296, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, new_AGEMA_signal_9898, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, new_AGEMA_signal_10618, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, new_AGEMA_signal_12433, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, new_AGEMA_signal_11299, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, new_AGEMA_signal_11302, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12438, new_AGEMA_signal_12437, new_AGEMA_signal_12436, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, new_AGEMA_signal_9892, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, new_AGEMA_signal_11305, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_11310, new_AGEMA_signal_11309, new_AGEMA_signal_11308, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, new_AGEMA_signal_10609, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, new_AGEMA_signal_11887, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, new_AGEMA_signal_12439, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, new_AGEMA_signal_12442, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, new_AGEMA_signal_10618, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, new_AGEMA_signal_11890, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_11310, new_AGEMA_signal_11309, new_AGEMA_signal_11308, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, new_AGEMA_signal_11893, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, new_AGEMA_signal_11302, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, new_AGEMA_signal_12445, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12450, new_AGEMA_signal_12449, new_AGEMA_signal_12448, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, new_AGEMA_signal_12451, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, new_AGEMA_signal_12454, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, new_AGEMA_signal_11299, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, new_AGEMA_signal_12457, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, new_AGEMA_signal_11305, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_12462, new_AGEMA_signal_12461, new_AGEMA_signal_12460, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, new_AGEMA_signal_12445, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_12438, new_AGEMA_signal_12437, new_AGEMA_signal_12436, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, new_AGEMA_signal_12451, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, new_AGEMA_signal_11887, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, new_AGEMA_signal_12457, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, new_AGEMA_signal_12442, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, new_AGEMA_signal_12439, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, new_AGEMA_signal_11890, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_12450, new_AGEMA_signal_12449, new_AGEMA_signal_12448, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_12462, new_AGEMA_signal_12461, new_AGEMA_signal_12460, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, new_AGEMA_signal_12433, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, new_AGEMA_signal_12454, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, new_AGEMA_signal_11893, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_28432, new_AGEMA_signal_28429, new_AGEMA_signal_28426, new_AGEMA_signal_28423}), .clk (clk), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_28444, new_AGEMA_signal_28441, new_AGEMA_signal_28438, new_AGEMA_signal_28435}), .clk (clk), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, new_AGEMA_signal_9913, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_28456, new_AGEMA_signal_28453, new_AGEMA_signal_28450, new_AGEMA_signal_28447}), .clk (clk), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_28468, new_AGEMA_signal_28465, new_AGEMA_signal_28462, new_AGEMA_signal_28459}), .clk (clk), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, new_AGEMA_signal_10627, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_28480, new_AGEMA_signal_28477, new_AGEMA_signal_28474, new_AGEMA_signal_28471}), .clk (clk), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110], Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_28492, new_AGEMA_signal_28489, new_AGEMA_signal_28486, new_AGEMA_signal_28483}), .clk (clk), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_28504, new_AGEMA_signal_28501, new_AGEMA_signal_28498, new_AGEMA_signal_28495}), .clk (clk), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_28516, new_AGEMA_signal_28513, new_AGEMA_signal_28510, new_AGEMA_signal_28507}), .clk (clk), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_28528, new_AGEMA_signal_28525, new_AGEMA_signal_28522, new_AGEMA_signal_28519}), .clk (clk), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, new_AGEMA_signal_10633, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_28540, new_AGEMA_signal_28537, new_AGEMA_signal_28534, new_AGEMA_signal_28531}), .clk (clk), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170], Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_28552, new_AGEMA_signal_28549, new_AGEMA_signal_28546, new_AGEMA_signal_28543}), .clk (clk), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_28564, new_AGEMA_signal_28561, new_AGEMA_signal_28558, new_AGEMA_signal_28555}), .clk (clk), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, new_AGEMA_signal_9928, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_28576, new_AGEMA_signal_28573, new_AGEMA_signal_28570, new_AGEMA_signal_28567}), .clk (clk), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_28588, new_AGEMA_signal_28585, new_AGEMA_signal_28582, new_AGEMA_signal_28579}), .clk (clk), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_28600, new_AGEMA_signal_28597, new_AGEMA_signal_28594, new_AGEMA_signal_28591}), .clk (clk), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230], Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, new_AGEMA_signal_9934, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_28612, new_AGEMA_signal_28609, new_AGEMA_signal_28606, new_AGEMA_signal_28603}), .clk (clk), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_28624, new_AGEMA_signal_28621, new_AGEMA_signal_28618, new_AGEMA_signal_28615}), .clk (clk), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_28636, new_AGEMA_signal_28633, new_AGEMA_signal_28630, new_AGEMA_signal_28627}), .clk (clk), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, new_AGEMA_signal_10645, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, new_AGEMA_signal_9913, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, new_AGEMA_signal_10633, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, new_AGEMA_signal_10627, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, new_AGEMA_signal_11326, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, new_AGEMA_signal_11326, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, new_AGEMA_signal_9934, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, new_AGEMA_signal_10654, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, new_AGEMA_signal_12466, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, new_AGEMA_signal_11329, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, new_AGEMA_signal_11332, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, new_AGEMA_signal_12469, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, new_AGEMA_signal_9928, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, new_AGEMA_signal_11335, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, new_AGEMA_signal_11338, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, new_AGEMA_signal_10645, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, new_AGEMA_signal_11914, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_12474, new_AGEMA_signal_12473, new_AGEMA_signal_12472, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, new_AGEMA_signal_12475, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, new_AGEMA_signal_10654, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, new_AGEMA_signal_11917, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, new_AGEMA_signal_11338, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, new_AGEMA_signal_11920, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, new_AGEMA_signal_11332, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, new_AGEMA_signal_12478, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, new_AGEMA_signal_12481, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12486, new_AGEMA_signal_12485, new_AGEMA_signal_12484, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, new_AGEMA_signal_12487, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, new_AGEMA_signal_11329, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, new_AGEMA_signal_12490, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, new_AGEMA_signal_11335, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, new_AGEMA_signal_12493, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, new_AGEMA_signal_12478, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, new_AGEMA_signal_12469, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_12486, new_AGEMA_signal_12485, new_AGEMA_signal_12484, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, new_AGEMA_signal_11914, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, new_AGEMA_signal_12490, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, new_AGEMA_signal_12475, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_12474, new_AGEMA_signal_12473, new_AGEMA_signal_12472, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, new_AGEMA_signal_11917, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, new_AGEMA_signal_12481, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, new_AGEMA_signal_12493, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, new_AGEMA_signal_12466, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, new_AGEMA_signal_12487, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, new_AGEMA_signal_11920, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_28648, new_AGEMA_signal_28645, new_AGEMA_signal_28642, new_AGEMA_signal_28639}), .clk (clk), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_28660, new_AGEMA_signal_28657, new_AGEMA_signal_28654, new_AGEMA_signal_28651}), .clk (clk), .r ({Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290], Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284]}), .c ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_28672, new_AGEMA_signal_28669, new_AGEMA_signal_28666, new_AGEMA_signal_28663}), .clk (clk), .r ({Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296]}), .c ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_28684, new_AGEMA_signal_28681, new_AGEMA_signal_28678, new_AGEMA_signal_28675}), .clk (clk), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308]}), .c ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, new_AGEMA_signal_10663, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_28696, new_AGEMA_signal_28693, new_AGEMA_signal_28690, new_AGEMA_signal_28687}), .clk (clk), .r ({Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_28708, new_AGEMA_signal_28705, new_AGEMA_signal_28702, new_AGEMA_signal_28699}), .clk (clk), .r ({Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332]}), .c ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_28720, new_AGEMA_signal_28717, new_AGEMA_signal_28714, new_AGEMA_signal_28711}), .clk (clk), .r ({Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350], Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344]}), .c ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_28732, new_AGEMA_signal_28729, new_AGEMA_signal_28726, new_AGEMA_signal_28723}), .clk (clk), .r ({Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356]}), .c ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_28744, new_AGEMA_signal_28741, new_AGEMA_signal_28738, new_AGEMA_signal_28735}), .clk (clk), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368]}), .c ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, new_AGEMA_signal_10669, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_28756, new_AGEMA_signal_28753, new_AGEMA_signal_28750, new_AGEMA_signal_28747}), .clk (clk), .r ({Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_28768, new_AGEMA_signal_28765, new_AGEMA_signal_28762, new_AGEMA_signal_28759}), .clk (clk), .r ({Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392]}), .c ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_28780, new_AGEMA_signal_28777, new_AGEMA_signal_28774, new_AGEMA_signal_28771}), .clk (clk), .r ({Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410], Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404]}), .c ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, new_AGEMA_signal_9964, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_28792, new_AGEMA_signal_28789, new_AGEMA_signal_28786, new_AGEMA_signal_28783}), .clk (clk), .r ({Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416]}), .c ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_28804, new_AGEMA_signal_28801, new_AGEMA_signal_28798, new_AGEMA_signal_28795}), .clk (clk), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428]}), .c ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_28816, new_AGEMA_signal_28813, new_AGEMA_signal_28810, new_AGEMA_signal_28807}), .clk (clk), .r ({Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, new_AGEMA_signal_9970, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_28828, new_AGEMA_signal_28825, new_AGEMA_signal_28822, new_AGEMA_signal_28819}), .clk (clk), .r ({Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452]}), .c ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_28840, new_AGEMA_signal_28837, new_AGEMA_signal_28834, new_AGEMA_signal_28831}), .clk (clk), .r ({Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470], Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464]}), .c ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_28852, new_AGEMA_signal_28849, new_AGEMA_signal_28846, new_AGEMA_signal_28843}), .clk (clk), .r ({Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476]}), .c ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, new_AGEMA_signal_10681, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, new_AGEMA_signal_10669, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, new_AGEMA_signal_10663, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, new_AGEMA_signal_11356, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, new_AGEMA_signal_11356, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, new_AGEMA_signal_9970, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, new_AGEMA_signal_10690, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, new_AGEMA_signal_12499, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, new_AGEMA_signal_11359, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, new_AGEMA_signal_11362, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, new_AGEMA_signal_12502, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, new_AGEMA_signal_9964, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, new_AGEMA_signal_11365, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, new_AGEMA_signal_11368, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, new_AGEMA_signal_10681, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, new_AGEMA_signal_11941, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, new_AGEMA_signal_12505, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_12510, new_AGEMA_signal_12509, new_AGEMA_signal_12508, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, new_AGEMA_signal_10690, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, new_AGEMA_signal_11944, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, new_AGEMA_signal_11368, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, new_AGEMA_signal_11947, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, new_AGEMA_signal_11362, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, new_AGEMA_signal_12511, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, new_AGEMA_signal_12514, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, new_AGEMA_signal_12517, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12522, new_AGEMA_signal_12521, new_AGEMA_signal_12520, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, new_AGEMA_signal_11359, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, new_AGEMA_signal_12523, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, new_AGEMA_signal_11365, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, new_AGEMA_signal_12526, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, new_AGEMA_signal_12511, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, new_AGEMA_signal_12502, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, new_AGEMA_signal_12517, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, new_AGEMA_signal_11941, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, new_AGEMA_signal_12523, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12510, new_AGEMA_signal_12509, new_AGEMA_signal_12508, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, new_AGEMA_signal_12505, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, new_AGEMA_signal_11944, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, new_AGEMA_signal_12514, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, new_AGEMA_signal_12526, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, new_AGEMA_signal_12499, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_12522, new_AGEMA_signal_12521, new_AGEMA_signal_12520, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, new_AGEMA_signal_11947, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_28864, new_AGEMA_signal_28861, new_AGEMA_signal_28858, new_AGEMA_signal_28855}), .clk (clk), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488]}), .c ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_28876, new_AGEMA_signal_28873, new_AGEMA_signal_28870, new_AGEMA_signal_28867}), .clk (clk), .r ({Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_28888, new_AGEMA_signal_28885, new_AGEMA_signal_28882, new_AGEMA_signal_28879}), .clk (clk), .r ({Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512]}), .c ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_28900, new_AGEMA_signal_28897, new_AGEMA_signal_28894, new_AGEMA_signal_28891}), .clk (clk), .r ({Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530], Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524]}), .c ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, new_AGEMA_signal_10699, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_28912, new_AGEMA_signal_28909, new_AGEMA_signal_28906, new_AGEMA_signal_28903}), .clk (clk), .r ({Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536]}), .c ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_28924, new_AGEMA_signal_28921, new_AGEMA_signal_28918, new_AGEMA_signal_28915}), .clk (clk), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548]}), .c ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_28936, new_AGEMA_signal_28933, new_AGEMA_signal_28930, new_AGEMA_signal_28927}), .clk (clk), .r ({Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_28948, new_AGEMA_signal_28945, new_AGEMA_signal_28942, new_AGEMA_signal_28939}), .clk (clk), .r ({Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572]}), .c ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_28960, new_AGEMA_signal_28957, new_AGEMA_signal_28954, new_AGEMA_signal_28951}), .clk (clk), .r ({Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590], Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584]}), .c ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, new_AGEMA_signal_10705, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_28972, new_AGEMA_signal_28969, new_AGEMA_signal_28966, new_AGEMA_signal_28963}), .clk (clk), .r ({Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596]}), .c ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_28984, new_AGEMA_signal_28981, new_AGEMA_signal_28978, new_AGEMA_signal_28975}), .clk (clk), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608]}), .c ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_28996, new_AGEMA_signal_28993, new_AGEMA_signal_28990, new_AGEMA_signal_28987}), .clk (clk), .r ({Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, new_AGEMA_signal_10000, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_29008, new_AGEMA_signal_29005, new_AGEMA_signal_29002, new_AGEMA_signal_28999}), .clk (clk), .r ({Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632]}), .c ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_29020, new_AGEMA_signal_29017, new_AGEMA_signal_29014, new_AGEMA_signal_29011}), .clk (clk), .r ({Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650], Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644]}), .c ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_29032, new_AGEMA_signal_29029, new_AGEMA_signal_29026, new_AGEMA_signal_29023}), .clk (clk), .r ({Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656]}), .c ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_29044, new_AGEMA_signal_29041, new_AGEMA_signal_29038, new_AGEMA_signal_29035}), .clk (clk), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668]}), .c ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_29056, new_AGEMA_signal_29053, new_AGEMA_signal_29050, new_AGEMA_signal_29047}), .clk (clk), .r ({Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_29068, new_AGEMA_signal_29065, new_AGEMA_signal_29062, new_AGEMA_signal_29059}), .clk (clk), .r ({Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692]}), .c ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, new_AGEMA_signal_10717, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, new_AGEMA_signal_10705, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, new_AGEMA_signal_10699, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, new_AGEMA_signal_11386, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, new_AGEMA_signal_11386, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, new_AGEMA_signal_10726, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12534, new_AGEMA_signal_12533, new_AGEMA_signal_12532, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, new_AGEMA_signal_11389, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, new_AGEMA_signal_11392, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, new_AGEMA_signal_12535, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, new_AGEMA_signal_10000, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, new_AGEMA_signal_11395, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, new_AGEMA_signal_11398, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, new_AGEMA_signal_10717, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, new_AGEMA_signal_11968, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, new_AGEMA_signal_12538, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, new_AGEMA_signal_12541, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, new_AGEMA_signal_10726, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, new_AGEMA_signal_11971, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, new_AGEMA_signal_11398, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, new_AGEMA_signal_11974, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, new_AGEMA_signal_11392, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12546, new_AGEMA_signal_12545, new_AGEMA_signal_12544, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, new_AGEMA_signal_12547, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, new_AGEMA_signal_12550, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, new_AGEMA_signal_12553, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, new_AGEMA_signal_11389, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_12558, new_AGEMA_signal_12557, new_AGEMA_signal_12556, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, new_AGEMA_signal_11395, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, new_AGEMA_signal_12559, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12546, new_AGEMA_signal_12545, new_AGEMA_signal_12544, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, new_AGEMA_signal_12535, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, new_AGEMA_signal_12550, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, new_AGEMA_signal_11968, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_12558, new_AGEMA_signal_12557, new_AGEMA_signal_12556, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, new_AGEMA_signal_12541, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, new_AGEMA_signal_12538, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, new_AGEMA_signal_11971, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, new_AGEMA_signal_12547, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, new_AGEMA_signal_12559, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_12534, new_AGEMA_signal_12533, new_AGEMA_signal_12532, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, new_AGEMA_signal_12553, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, new_AGEMA_signal_11974, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_29080, new_AGEMA_signal_29077, new_AGEMA_signal_29074, new_AGEMA_signal_29071}), .clk (clk), .r ({Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710], Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704]}), .c ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_29092, new_AGEMA_signal_29089, new_AGEMA_signal_29086, new_AGEMA_signal_29083}), .clk (clk), .r ({Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716]}), .c ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_29104, new_AGEMA_signal_29101, new_AGEMA_signal_29098, new_AGEMA_signal_29095}), .clk (clk), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728]}), .c ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_29116, new_AGEMA_signal_29113, new_AGEMA_signal_29110, new_AGEMA_signal_29107}), .clk (clk), .r ({Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, new_AGEMA_signal_10735, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_29128, new_AGEMA_signal_29125, new_AGEMA_signal_29122, new_AGEMA_signal_29119}), .clk (clk), .r ({Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752]}), .c ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_29140, new_AGEMA_signal_29137, new_AGEMA_signal_29134, new_AGEMA_signal_29131}), .clk (clk), .r ({Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770], Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764]}), .c ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_29152, new_AGEMA_signal_29149, new_AGEMA_signal_29146, new_AGEMA_signal_29143}), .clk (clk), .r ({Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776]}), .c ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_29164, new_AGEMA_signal_29161, new_AGEMA_signal_29158, new_AGEMA_signal_29155}), .clk (clk), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788]}), .c ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_29176, new_AGEMA_signal_29173, new_AGEMA_signal_29170, new_AGEMA_signal_29167}), .clk (clk), .r ({Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, new_AGEMA_signal_10741, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_29188, new_AGEMA_signal_29185, new_AGEMA_signal_29182, new_AGEMA_signal_29179}), .clk (clk), .r ({Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812]}), .c ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_29200, new_AGEMA_signal_29197, new_AGEMA_signal_29194, new_AGEMA_signal_29191}), .clk (clk), .r ({Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830], Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824]}), .c ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_29212, new_AGEMA_signal_29209, new_AGEMA_signal_29206, new_AGEMA_signal_29203}), .clk (clk), .r ({Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836]}), .c ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, new_AGEMA_signal_10036, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_29224, new_AGEMA_signal_29221, new_AGEMA_signal_29218, new_AGEMA_signal_29215}), .clk (clk), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848]}), .c ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_29236, new_AGEMA_signal_29233, new_AGEMA_signal_29230, new_AGEMA_signal_29227}), .clk (clk), .r ({Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_29248, new_AGEMA_signal_29245, new_AGEMA_signal_29242, new_AGEMA_signal_29239}), .clk (clk), .r ({Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872]}), .c ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, new_AGEMA_signal_10042, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_29260, new_AGEMA_signal_29257, new_AGEMA_signal_29254, new_AGEMA_signal_29251}), .clk (clk), .r ({Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890], Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884]}), .c ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_29272, new_AGEMA_signal_29269, new_AGEMA_signal_29266, new_AGEMA_signal_29263}), .clk (clk), .r ({Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896]}), .c ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_29284, new_AGEMA_signal_29281, new_AGEMA_signal_29278, new_AGEMA_signal_29275}), .clk (clk), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908]}), .c ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, new_AGEMA_signal_10753, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, new_AGEMA_signal_10741, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, new_AGEMA_signal_10735, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, new_AGEMA_signal_11416, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, new_AGEMA_signal_11416, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, new_AGEMA_signal_10042, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, new_AGEMA_signal_10762, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, new_AGEMA_signal_12565, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, new_AGEMA_signal_11419, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, new_AGEMA_signal_11422, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_12570, new_AGEMA_signal_12569, new_AGEMA_signal_12568, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, new_AGEMA_signal_10036, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, new_AGEMA_signal_11425, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, new_AGEMA_signal_11428, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, new_AGEMA_signal_10753, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, new_AGEMA_signal_11995, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, new_AGEMA_signal_12571, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, new_AGEMA_signal_12574, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, new_AGEMA_signal_10762, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, new_AGEMA_signal_11998, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, new_AGEMA_signal_11428, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, new_AGEMA_signal_12001, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, new_AGEMA_signal_11422, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, new_AGEMA_signal_12577, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_12582, new_AGEMA_signal_12581, new_AGEMA_signal_12580, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, new_AGEMA_signal_12583, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, new_AGEMA_signal_12586, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, new_AGEMA_signal_11419, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, new_AGEMA_signal_12589, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, new_AGEMA_signal_11425, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_12594, new_AGEMA_signal_12593, new_AGEMA_signal_12592, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, new_AGEMA_signal_12577, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_12570, new_AGEMA_signal_12569, new_AGEMA_signal_12568, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, new_AGEMA_signal_12583, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, new_AGEMA_signal_11995, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, new_AGEMA_signal_12589, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, new_AGEMA_signal_12574, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, new_AGEMA_signal_12571, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, new_AGEMA_signal_11998, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_12582, new_AGEMA_signal_12581, new_AGEMA_signal_12580, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_12594, new_AGEMA_signal_12593, new_AGEMA_signal_12592, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, new_AGEMA_signal_12565, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, new_AGEMA_signal_12586, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, new_AGEMA_signal_12001, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_29296, new_AGEMA_signal_29293, new_AGEMA_signal_29290, new_AGEMA_signal_29287}), .clk (clk), .r ({Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_29308, new_AGEMA_signal_29305, new_AGEMA_signal_29302, new_AGEMA_signal_29299}), .clk (clk), .r ({Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932]}), .c ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_29320, new_AGEMA_signal_29317, new_AGEMA_signal_29314, new_AGEMA_signal_29311}), .clk (clk), .r ({Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950], Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944]}), .c ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_29332, new_AGEMA_signal_29329, new_AGEMA_signal_29326, new_AGEMA_signal_29323}), .clk (clk), .r ({Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956]}), .c ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, new_AGEMA_signal_10771, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_29344, new_AGEMA_signal_29341, new_AGEMA_signal_29338, new_AGEMA_signal_29335}), .clk (clk), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968]}), .c ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_29356, new_AGEMA_signal_29353, new_AGEMA_signal_29350, new_AGEMA_signal_29347}), .clk (clk), .r ({Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_29368, new_AGEMA_signal_29365, new_AGEMA_signal_29362, new_AGEMA_signal_29359}), .clk (clk), .r ({Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992]}), .c ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_29380, new_AGEMA_signal_29377, new_AGEMA_signal_29374, new_AGEMA_signal_29371}), .clk (clk), .r ({Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010], Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004]}), .c ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_29392, new_AGEMA_signal_29389, new_AGEMA_signal_29386, new_AGEMA_signal_29383}), .clk (clk), .r ({Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016]}), .c ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, new_AGEMA_signal_10777, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_29404, new_AGEMA_signal_29401, new_AGEMA_signal_29398, new_AGEMA_signal_29395}), .clk (clk), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028]}), .c ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_29416, new_AGEMA_signal_29413, new_AGEMA_signal_29410, new_AGEMA_signal_29407}), .clk (clk), .r ({Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_29428, new_AGEMA_signal_29425, new_AGEMA_signal_29422, new_AGEMA_signal_29419}), .clk (clk), .r ({Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052]}), .c ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, new_AGEMA_signal_10072, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_29440, new_AGEMA_signal_29437, new_AGEMA_signal_29434, new_AGEMA_signal_29431}), .clk (clk), .r ({Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070], Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064]}), .c ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_29452, new_AGEMA_signal_29449, new_AGEMA_signal_29446, new_AGEMA_signal_29443}), .clk (clk), .r ({Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076]}), .c ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_29464, new_AGEMA_signal_29461, new_AGEMA_signal_29458, new_AGEMA_signal_29455}), .clk (clk), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088]}), .c ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, new_AGEMA_signal_10078, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_29476, new_AGEMA_signal_29473, new_AGEMA_signal_29470, new_AGEMA_signal_29467}), .clk (clk), .r ({Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_29488, new_AGEMA_signal_29485, new_AGEMA_signal_29482, new_AGEMA_signal_29479}), .clk (clk), .r ({Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112]}), .c ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_29500, new_AGEMA_signal_29497, new_AGEMA_signal_29494, new_AGEMA_signal_29491}), .clk (clk), .r ({Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130], Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124]}), .c ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, new_AGEMA_signal_10789, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, new_AGEMA_signal_10777, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, new_AGEMA_signal_10771, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, new_AGEMA_signal_11446, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, new_AGEMA_signal_11446, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, new_AGEMA_signal_10078, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, new_AGEMA_signal_10798, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, new_AGEMA_signal_12598, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, new_AGEMA_signal_11449, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, new_AGEMA_signal_11452, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, new_AGEMA_signal_12601, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, new_AGEMA_signal_10072, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, new_AGEMA_signal_11455, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, new_AGEMA_signal_11458, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, new_AGEMA_signal_10789, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, new_AGEMA_signal_12022, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_12606, new_AGEMA_signal_12605, new_AGEMA_signal_12604, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, new_AGEMA_signal_12607, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, new_AGEMA_signal_10798, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, new_AGEMA_signal_12025, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, new_AGEMA_signal_11458, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, new_AGEMA_signal_12028, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, new_AGEMA_signal_11452, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, new_AGEMA_signal_12610, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, new_AGEMA_signal_12613, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_12618, new_AGEMA_signal_12617, new_AGEMA_signal_12616, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, new_AGEMA_signal_12619, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, new_AGEMA_signal_11449, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, new_AGEMA_signal_12622, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, new_AGEMA_signal_11455, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, new_AGEMA_signal_12625, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, new_AGEMA_signal_12610, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, new_AGEMA_signal_12601, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_12618, new_AGEMA_signal_12617, new_AGEMA_signal_12616, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, new_AGEMA_signal_12022, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, new_AGEMA_signal_12622, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, new_AGEMA_signal_12607, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_12606, new_AGEMA_signal_12605, new_AGEMA_signal_12604, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, new_AGEMA_signal_12025, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, new_AGEMA_signal_12613, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, new_AGEMA_signal_12625, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, new_AGEMA_signal_12598, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, new_AGEMA_signal_12619, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, new_AGEMA_signal_12028, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_29512, new_AGEMA_signal_29509, new_AGEMA_signal_29506, new_AGEMA_signal_29503}), .clk (clk), .r ({Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136]}), .c ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_29524, new_AGEMA_signal_29521, new_AGEMA_signal_29518, new_AGEMA_signal_29515}), .clk (clk), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148]}), .c ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_29536, new_AGEMA_signal_29533, new_AGEMA_signal_29530, new_AGEMA_signal_29527}), .clk (clk), .r ({Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_29548, new_AGEMA_signal_29545, new_AGEMA_signal_29542, new_AGEMA_signal_29539}), .clk (clk), .r ({Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172]}), .c ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, new_AGEMA_signal_10807, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_29560, new_AGEMA_signal_29557, new_AGEMA_signal_29554, new_AGEMA_signal_29551}), .clk (clk), .r ({Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190], Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184]}), .c ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_29572, new_AGEMA_signal_29569, new_AGEMA_signal_29566, new_AGEMA_signal_29563}), .clk (clk), .r ({Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196]}), .c ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_29584, new_AGEMA_signal_29581, new_AGEMA_signal_29578, new_AGEMA_signal_29575}), .clk (clk), .r ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208]}), .c ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_29596, new_AGEMA_signal_29593, new_AGEMA_signal_29590, new_AGEMA_signal_29587}), .clk (clk), .r ({Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .c ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_29608, new_AGEMA_signal_29605, new_AGEMA_signal_29602, new_AGEMA_signal_29599}), .clk (clk), .r ({Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232]}), .c ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, new_AGEMA_signal_10813, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_29620, new_AGEMA_signal_29617, new_AGEMA_signal_29614, new_AGEMA_signal_29611}), .clk (clk), .r ({Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250], Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244]}), .c ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_29632, new_AGEMA_signal_29629, new_AGEMA_signal_29626, new_AGEMA_signal_29623}), .clk (clk), .r ({Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256]}), .c ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_29644, new_AGEMA_signal_29641, new_AGEMA_signal_29638, new_AGEMA_signal_29635}), .clk (clk), .r ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268]}), .c ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, new_AGEMA_signal_10108, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_29656, new_AGEMA_signal_29653, new_AGEMA_signal_29650, new_AGEMA_signal_29647}), .clk (clk), .r ({Fresh[5291], Fresh[5290], Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .c ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_29668, new_AGEMA_signal_29665, new_AGEMA_signal_29662, new_AGEMA_signal_29659}), .clk (clk), .r ({Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300], Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292]}), .c ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, new_AGEMA_signal_10111, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_29680, new_AGEMA_signal_29677, new_AGEMA_signal_29674, new_AGEMA_signal_29671}), .clk (clk), .r ({Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310], Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304]}), .c ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, new_AGEMA_signal_10114, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_29692, new_AGEMA_signal_29689, new_AGEMA_signal_29686, new_AGEMA_signal_29683}), .clk (clk), .r ({Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320], Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316]}), .c ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_29704, new_AGEMA_signal_29701, new_AGEMA_signal_29698, new_AGEMA_signal_29695}), .clk (clk), .r ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330], Fresh[5329], Fresh[5328]}), .c ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_29716, new_AGEMA_signal_29713, new_AGEMA_signal_29710, new_AGEMA_signal_29707}), .clk (clk), .r ({Fresh[5351], Fresh[5350], Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .c ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, new_AGEMA_signal_10825, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, new_AGEMA_signal_10813, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, new_AGEMA_signal_10807, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, new_AGEMA_signal_11476, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, new_AGEMA_signal_11476, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, new_AGEMA_signal_10111, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, new_AGEMA_signal_10114, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, new_AGEMA_signal_10834, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, new_AGEMA_signal_12631, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, new_AGEMA_signal_11479, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, new_AGEMA_signal_11482, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, new_AGEMA_signal_12634, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, new_AGEMA_signal_10108, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, new_AGEMA_signal_11485, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, new_AGEMA_signal_11488, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, new_AGEMA_signal_10825, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, new_AGEMA_signal_12049, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, new_AGEMA_signal_12637, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_12642, new_AGEMA_signal_12641, new_AGEMA_signal_12640, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, new_AGEMA_signal_10834, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, new_AGEMA_signal_12052, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, new_AGEMA_signal_11488, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, new_AGEMA_signal_12055, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, new_AGEMA_signal_11482, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, new_AGEMA_signal_12643, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, new_AGEMA_signal_12646, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, new_AGEMA_signal_12649, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_12654, new_AGEMA_signal_12653, new_AGEMA_signal_12652, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, new_AGEMA_signal_11479, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, new_AGEMA_signal_12655, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, new_AGEMA_signal_11485, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, new_AGEMA_signal_12658, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, new_AGEMA_signal_12643, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, new_AGEMA_signal_12634, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, new_AGEMA_signal_12649, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, new_AGEMA_signal_12049, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, new_AGEMA_signal_12655, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12642, new_AGEMA_signal_12641, new_AGEMA_signal_12640, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, new_AGEMA_signal_12637, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, new_AGEMA_signal_12052, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, new_AGEMA_signal_12646, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, new_AGEMA_signal_12658, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, new_AGEMA_signal_12631, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_12654, new_AGEMA_signal_12653, new_AGEMA_signal_12652, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, new_AGEMA_signal_12055, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_29728, new_AGEMA_signal_29725, new_AGEMA_signal_29722, new_AGEMA_signal_29719}), .clk (clk), .r ({Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360], Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352]}), .c ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_29740, new_AGEMA_signal_29737, new_AGEMA_signal_29734, new_AGEMA_signal_29731}), .clk (clk), .r ({Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370], Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364]}), .c ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_29752, new_AGEMA_signal_29749, new_AGEMA_signal_29746, new_AGEMA_signal_29743}), .clk (clk), .r ({Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380], Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376]}), .c ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_29764, new_AGEMA_signal_29761, new_AGEMA_signal_29758, new_AGEMA_signal_29755}), .clk (clk), .r ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390], Fresh[5389], Fresh[5388]}), .c ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, new_AGEMA_signal_10843, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_29776, new_AGEMA_signal_29773, new_AGEMA_signal_29770, new_AGEMA_signal_29767}), .clk (clk), .r ({Fresh[5411], Fresh[5410], Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .c ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_29788, new_AGEMA_signal_29785, new_AGEMA_signal_29782, new_AGEMA_signal_29779}), .clk (clk), .r ({Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420], Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412]}), .c ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_29800, new_AGEMA_signal_29797, new_AGEMA_signal_29794, new_AGEMA_signal_29791}), .clk (clk), .r ({Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430], Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424]}), .c ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_29812, new_AGEMA_signal_29809, new_AGEMA_signal_29806, new_AGEMA_signal_29803}), .clk (clk), .r ({Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440], Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436]}), .c ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_29824, new_AGEMA_signal_29821, new_AGEMA_signal_29818, new_AGEMA_signal_29815}), .clk (clk), .r ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450], Fresh[5449], Fresh[5448]}), .c ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, new_AGEMA_signal_10849, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_29836, new_AGEMA_signal_29833, new_AGEMA_signal_29830, new_AGEMA_signal_29827}), .clk (clk), .r ({Fresh[5471], Fresh[5470], Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .c ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_29848, new_AGEMA_signal_29845, new_AGEMA_signal_29842, new_AGEMA_signal_29839}), .clk (clk), .r ({Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480], Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472]}), .c ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_29860, new_AGEMA_signal_29857, new_AGEMA_signal_29854, new_AGEMA_signal_29851}), .clk (clk), .r ({Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490], Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484]}), .c ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, new_AGEMA_signal_10144, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_29872, new_AGEMA_signal_29869, new_AGEMA_signal_29866, new_AGEMA_signal_29863}), .clk (clk), .r ({Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500], Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496]}), .c ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_29884, new_AGEMA_signal_29881, new_AGEMA_signal_29878, new_AGEMA_signal_29875}), .clk (clk), .r ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510], Fresh[5509], Fresh[5508]}), .c ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_29896, new_AGEMA_signal_29893, new_AGEMA_signal_29890, new_AGEMA_signal_29887}), .clk (clk), .r ({Fresh[5531], Fresh[5530], Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .c ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, new_AGEMA_signal_10150, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_29908, new_AGEMA_signal_29905, new_AGEMA_signal_29902, new_AGEMA_signal_29899}), .clk (clk), .r ({Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540], Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532]}), .c ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_29920, new_AGEMA_signal_29917, new_AGEMA_signal_29914, new_AGEMA_signal_29911}), .clk (clk), .r ({Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550], Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544]}), .c ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_29932, new_AGEMA_signal_29929, new_AGEMA_signal_29926, new_AGEMA_signal_29923}), .clk (clk), .r ({Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560], Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556]}), .c ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, new_AGEMA_signal_10861, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, new_AGEMA_signal_10849, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, new_AGEMA_signal_10843, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, new_AGEMA_signal_11506, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, new_AGEMA_signal_11506, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, new_AGEMA_signal_10150, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, new_AGEMA_signal_10870, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_12666, new_AGEMA_signal_12665, new_AGEMA_signal_12664, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, new_AGEMA_signal_11509, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, new_AGEMA_signal_11512, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, new_AGEMA_signal_12667, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, new_AGEMA_signal_10144, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, new_AGEMA_signal_11515, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, new_AGEMA_signal_11518, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, new_AGEMA_signal_10861, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, new_AGEMA_signal_12076, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, new_AGEMA_signal_12670, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, new_AGEMA_signal_12673, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, new_AGEMA_signal_10870, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, new_AGEMA_signal_12079, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, new_AGEMA_signal_11518, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, new_AGEMA_signal_12082, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, new_AGEMA_signal_11512, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_12678, new_AGEMA_signal_12677, new_AGEMA_signal_12676, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, new_AGEMA_signal_12679, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, new_AGEMA_signal_12682, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, new_AGEMA_signal_12685, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, new_AGEMA_signal_11509, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_12690, new_AGEMA_signal_12689, new_AGEMA_signal_12688, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, new_AGEMA_signal_11515, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, new_AGEMA_signal_12691, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12678, new_AGEMA_signal_12677, new_AGEMA_signal_12676, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, new_AGEMA_signal_12667, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, new_AGEMA_signal_12682, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, new_AGEMA_signal_12076, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_12690, new_AGEMA_signal_12689, new_AGEMA_signal_12688, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, new_AGEMA_signal_12673, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, new_AGEMA_signal_12670, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, new_AGEMA_signal_12079, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, new_AGEMA_signal_12679, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, new_AGEMA_signal_12691, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_12666, new_AGEMA_signal_12665, new_AGEMA_signal_12664, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, new_AGEMA_signal_12685, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, new_AGEMA_signal_12082, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_29944, new_AGEMA_signal_29941, new_AGEMA_signal_29938, new_AGEMA_signal_29935}), .clk (clk), .r ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570], Fresh[5569], Fresh[5568]}), .c ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_29956, new_AGEMA_signal_29953, new_AGEMA_signal_29950, new_AGEMA_signal_29947}), .clk (clk), .r ({Fresh[5591], Fresh[5590], Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .c ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, new_AGEMA_signal_10165, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_29968, new_AGEMA_signal_29965, new_AGEMA_signal_29962, new_AGEMA_signal_29959}), .clk (clk), .r ({Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600], Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592]}), .c ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_29980, new_AGEMA_signal_29977, new_AGEMA_signal_29974, new_AGEMA_signal_29971}), .clk (clk), .r ({Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610], Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604]}), .c ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, new_AGEMA_signal_10879, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_29992, new_AGEMA_signal_29989, new_AGEMA_signal_29986, new_AGEMA_signal_29983}), .clk (clk), .r ({Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620], Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616]}), .c ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_30004, new_AGEMA_signal_30001, new_AGEMA_signal_29998, new_AGEMA_signal_29995}), .clk (clk), .r ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630], Fresh[5629], Fresh[5628]}), .c ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_30016, new_AGEMA_signal_30013, new_AGEMA_signal_30010, new_AGEMA_signal_30007}), .clk (clk), .r ({Fresh[5651], Fresh[5650], Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .c ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_30028, new_AGEMA_signal_30025, new_AGEMA_signal_30022, new_AGEMA_signal_30019}), .clk (clk), .r ({Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660], Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652]}), .c ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_30040, new_AGEMA_signal_30037, new_AGEMA_signal_30034, new_AGEMA_signal_30031}), .clk (clk), .r ({Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670], Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664]}), .c ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, new_AGEMA_signal_10885, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_30052, new_AGEMA_signal_30049, new_AGEMA_signal_30046, new_AGEMA_signal_30043}), .clk (clk), .r ({Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680], Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676]}), .c ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_30064, new_AGEMA_signal_30061, new_AGEMA_signal_30058, new_AGEMA_signal_30055}), .clk (clk), .r ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690], Fresh[5689], Fresh[5688]}), .c ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_30076, new_AGEMA_signal_30073, new_AGEMA_signal_30070, new_AGEMA_signal_30067}), .clk (clk), .r ({Fresh[5711], Fresh[5710], Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .c ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, new_AGEMA_signal_10180, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_30088, new_AGEMA_signal_30085, new_AGEMA_signal_30082, new_AGEMA_signal_30079}), .clk (clk), .r ({Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720], Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712]}), .c ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_30100, new_AGEMA_signal_30097, new_AGEMA_signal_30094, new_AGEMA_signal_30091}), .clk (clk), .r ({Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730], Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724]}), .c ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, new_AGEMA_signal_10183, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_30112, new_AGEMA_signal_30109, new_AGEMA_signal_30106, new_AGEMA_signal_30103}), .clk (clk), .r ({Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740], Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736]}), .c ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, new_AGEMA_signal_10186, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_30124, new_AGEMA_signal_30121, new_AGEMA_signal_30118, new_AGEMA_signal_30115}), .clk (clk), .r ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750], Fresh[5749], Fresh[5748]}), .c ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_30136, new_AGEMA_signal_30133, new_AGEMA_signal_30130, new_AGEMA_signal_30127}), .clk (clk), .r ({Fresh[5771], Fresh[5770], Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .c ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_30148, new_AGEMA_signal_30145, new_AGEMA_signal_30142, new_AGEMA_signal_30139}), .clk (clk), .r ({Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780], Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772]}), .c ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, new_AGEMA_signal_10897, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, new_AGEMA_signal_10165, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, new_AGEMA_signal_10885, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, new_AGEMA_signal_10879, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, new_AGEMA_signal_11536, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, new_AGEMA_signal_11536, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, new_AGEMA_signal_10183, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, new_AGEMA_signal_10186, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, new_AGEMA_signal_10906, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, new_AGEMA_signal_12697, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, new_AGEMA_signal_11539, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, new_AGEMA_signal_11542, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_12702, new_AGEMA_signal_12701, new_AGEMA_signal_12700, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, new_AGEMA_signal_10180, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, new_AGEMA_signal_11545, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, new_AGEMA_signal_11548, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, new_AGEMA_signal_10897, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, new_AGEMA_signal_12103, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, new_AGEMA_signal_12703, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, new_AGEMA_signal_12706, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, new_AGEMA_signal_10906, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_12108, new_AGEMA_signal_12107, new_AGEMA_signal_12106, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, new_AGEMA_signal_11548, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, new_AGEMA_signal_12109, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, new_AGEMA_signal_11542, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, new_AGEMA_signal_12709, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_12714, new_AGEMA_signal_12713, new_AGEMA_signal_12712, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, new_AGEMA_signal_12715, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, new_AGEMA_signal_12718, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, new_AGEMA_signal_11539, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, new_AGEMA_signal_12721, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, new_AGEMA_signal_11545, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_12726, new_AGEMA_signal_12725, new_AGEMA_signal_12724, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, new_AGEMA_signal_12709, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_12702, new_AGEMA_signal_12701, new_AGEMA_signal_12700, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, new_AGEMA_signal_12715, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, new_AGEMA_signal_12103, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, new_AGEMA_signal_12721, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, new_AGEMA_signal_12706, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, new_AGEMA_signal_12703, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_12108, new_AGEMA_signal_12107, new_AGEMA_signal_12106, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_12714, new_AGEMA_signal_12713, new_AGEMA_signal_12712, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_12726, new_AGEMA_signal_12725, new_AGEMA_signal_12724, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, new_AGEMA_signal_12697, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, new_AGEMA_signal_12718, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, new_AGEMA_signal_12109, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_30160, new_AGEMA_signal_30157, new_AGEMA_signal_30154, new_AGEMA_signal_30151}), .clk (clk), .r ({Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790], Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784]}), .c ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_30172, new_AGEMA_signal_30169, new_AGEMA_signal_30166, new_AGEMA_signal_30163}), .clk (clk), .r ({Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800], Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796]}), .c ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, new_AGEMA_signal_10201, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_30184, new_AGEMA_signal_30181, new_AGEMA_signal_30178, new_AGEMA_signal_30175}), .clk (clk), .r ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810], Fresh[5809], Fresh[5808]}), .c ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_30196, new_AGEMA_signal_30193, new_AGEMA_signal_30190, new_AGEMA_signal_30187}), .clk (clk), .r ({Fresh[5831], Fresh[5830], Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .c ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, new_AGEMA_signal_10915, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_30208, new_AGEMA_signal_30205, new_AGEMA_signal_30202, new_AGEMA_signal_30199}), .clk (clk), .r ({Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840], Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832]}), .c ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_30220, new_AGEMA_signal_30217, new_AGEMA_signal_30214, new_AGEMA_signal_30211}), .clk (clk), .r ({Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850], Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844]}), .c ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_30232, new_AGEMA_signal_30229, new_AGEMA_signal_30226, new_AGEMA_signal_30223}), .clk (clk), .r ({Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860], Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856]}), .c ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_30244, new_AGEMA_signal_30241, new_AGEMA_signal_30238, new_AGEMA_signal_30235}), .clk (clk), .r ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870], Fresh[5869], Fresh[5868]}), .c ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_30256, new_AGEMA_signal_30253, new_AGEMA_signal_30250, new_AGEMA_signal_30247}), .clk (clk), .r ({Fresh[5891], Fresh[5890], Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .c ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, new_AGEMA_signal_10921, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_30268, new_AGEMA_signal_30265, new_AGEMA_signal_30262, new_AGEMA_signal_30259}), .clk (clk), .r ({Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900], Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892]}), .c ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_30280, new_AGEMA_signal_30277, new_AGEMA_signal_30274, new_AGEMA_signal_30271}), .clk (clk), .r ({Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910], Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904]}), .c ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_30292, new_AGEMA_signal_30289, new_AGEMA_signal_30286, new_AGEMA_signal_30283}), .clk (clk), .r ({Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920], Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916]}), .c ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, new_AGEMA_signal_10216, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_30304, new_AGEMA_signal_30301, new_AGEMA_signal_30298, new_AGEMA_signal_30295}), .clk (clk), .r ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930], Fresh[5929], Fresh[5928]}), .c ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_30316, new_AGEMA_signal_30313, new_AGEMA_signal_30310, new_AGEMA_signal_30307}), .clk (clk), .r ({Fresh[5951], Fresh[5950], Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .c ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, new_AGEMA_signal_10219, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_30328, new_AGEMA_signal_30325, new_AGEMA_signal_30322, new_AGEMA_signal_30319}), .clk (clk), .r ({Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960], Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952]}), .c ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, new_AGEMA_signal_10222, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_30340, new_AGEMA_signal_30337, new_AGEMA_signal_30334, new_AGEMA_signal_30331}), .clk (clk), .r ({Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970], Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964]}), .c ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_30352, new_AGEMA_signal_30349, new_AGEMA_signal_30346, new_AGEMA_signal_30343}), .clk (clk), .r ({Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980], Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976]}), .c ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_30364, new_AGEMA_signal_30361, new_AGEMA_signal_30358, new_AGEMA_signal_30355}), .clk (clk), .r ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990], Fresh[5989], Fresh[5988]}), .c ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, new_AGEMA_signal_10933, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, new_AGEMA_signal_10201, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, new_AGEMA_signal_10921, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, new_AGEMA_signal_10915, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, new_AGEMA_signal_11566, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, new_AGEMA_signal_11566, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, new_AGEMA_signal_10219, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, new_AGEMA_signal_10222, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, new_AGEMA_signal_10942, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, new_AGEMA_signal_12730, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, new_AGEMA_signal_11569, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, new_AGEMA_signal_11572, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, new_AGEMA_signal_12733, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, new_AGEMA_signal_10216, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, new_AGEMA_signal_11575, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, new_AGEMA_signal_11578, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, new_AGEMA_signal_10933, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_12132, new_AGEMA_signal_12131, new_AGEMA_signal_12130, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_12738, new_AGEMA_signal_12737, new_AGEMA_signal_12736, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, new_AGEMA_signal_12739, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, new_AGEMA_signal_10942, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, new_AGEMA_signal_12133, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, new_AGEMA_signal_11578, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, new_AGEMA_signal_12136, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, new_AGEMA_signal_11572, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, new_AGEMA_signal_12742, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, new_AGEMA_signal_12745, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_12750, new_AGEMA_signal_12749, new_AGEMA_signal_12748, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, new_AGEMA_signal_12751, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, new_AGEMA_signal_11569, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, new_AGEMA_signal_12754, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, new_AGEMA_signal_11575, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, new_AGEMA_signal_12757, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, new_AGEMA_signal_12742, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, new_AGEMA_signal_12733, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_12750, new_AGEMA_signal_12749, new_AGEMA_signal_12748, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_12132, new_AGEMA_signal_12131, new_AGEMA_signal_12130, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, new_AGEMA_signal_12754, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, new_AGEMA_signal_12739, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_12738, new_AGEMA_signal_12737, new_AGEMA_signal_12736, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, new_AGEMA_signal_12133, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, new_AGEMA_signal_12745, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, new_AGEMA_signal_12757, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, new_AGEMA_signal_12730, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, new_AGEMA_signal_12751, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, new_AGEMA_signal_12136, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_30376, new_AGEMA_signal_30373, new_AGEMA_signal_30370, new_AGEMA_signal_30367}), .clk (clk), .r ({Fresh[6011], Fresh[6010], Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .c ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_30388, new_AGEMA_signal_30385, new_AGEMA_signal_30382, new_AGEMA_signal_30379}), .clk (clk), .r ({Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020], Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012]}), .c ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, new_AGEMA_signal_10237, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_30400, new_AGEMA_signal_30397, new_AGEMA_signal_30394, new_AGEMA_signal_30391}), .clk (clk), .r ({Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030], Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024]}), .c ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_30412, new_AGEMA_signal_30409, new_AGEMA_signal_30406, new_AGEMA_signal_30403}), .clk (clk), .r ({Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040], Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036]}), .c ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, new_AGEMA_signal_10951, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_30424, new_AGEMA_signal_30421, new_AGEMA_signal_30418, new_AGEMA_signal_30415}), .clk (clk), .r ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050], Fresh[6049], Fresh[6048]}), .c ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_30436, new_AGEMA_signal_30433, new_AGEMA_signal_30430, new_AGEMA_signal_30427}), .clk (clk), .r ({Fresh[6071], Fresh[6070], Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .c ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_30448, new_AGEMA_signal_30445, new_AGEMA_signal_30442, new_AGEMA_signal_30439}), .clk (clk), .r ({Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080], Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072]}), .c ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_30460, new_AGEMA_signal_30457, new_AGEMA_signal_30454, new_AGEMA_signal_30451}), .clk (clk), .r ({Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090], Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084]}), .c ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_30472, new_AGEMA_signal_30469, new_AGEMA_signal_30466, new_AGEMA_signal_30463}), .clk (clk), .r ({Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100], Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096]}), .c ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, new_AGEMA_signal_10957, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_30484, new_AGEMA_signal_30481, new_AGEMA_signal_30478, new_AGEMA_signal_30475}), .clk (clk), .r ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110], Fresh[6109], Fresh[6108]}), .c ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_30496, new_AGEMA_signal_30493, new_AGEMA_signal_30490, new_AGEMA_signal_30487}), .clk (clk), .r ({Fresh[6131], Fresh[6130], Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .c ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_30508, new_AGEMA_signal_30505, new_AGEMA_signal_30502, new_AGEMA_signal_30499}), .clk (clk), .r ({Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140], Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132]}), .c ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, new_AGEMA_signal_10252, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_30520, new_AGEMA_signal_30517, new_AGEMA_signal_30514, new_AGEMA_signal_30511}), .clk (clk), .r ({Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150], Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144]}), .c ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_30532, new_AGEMA_signal_30529, new_AGEMA_signal_30526, new_AGEMA_signal_30523}), .clk (clk), .r ({Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160], Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156]}), .c ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, new_AGEMA_signal_10255, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_30544, new_AGEMA_signal_30541, new_AGEMA_signal_30538, new_AGEMA_signal_30535}), .clk (clk), .r ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170], Fresh[6169], Fresh[6168]}), .c ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, new_AGEMA_signal_10258, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_30556, new_AGEMA_signal_30553, new_AGEMA_signal_30550, new_AGEMA_signal_30547}), .clk (clk), .r ({Fresh[6191], Fresh[6190], Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .c ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_30568, new_AGEMA_signal_30565, new_AGEMA_signal_30562, new_AGEMA_signal_30559}), .clk (clk), .r ({Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200], Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192]}), .c ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_30580, new_AGEMA_signal_30577, new_AGEMA_signal_30574, new_AGEMA_signal_30571}), .clk (clk), .r ({Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210], Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204]}), .c ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, new_AGEMA_signal_10969, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, new_AGEMA_signal_10237, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, new_AGEMA_signal_10957, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, new_AGEMA_signal_10951, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, new_AGEMA_signal_11596, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, new_AGEMA_signal_11596, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, new_AGEMA_signal_10255, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, new_AGEMA_signal_10258, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, new_AGEMA_signal_10978, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, new_AGEMA_signal_12763, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, new_AGEMA_signal_11599, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, new_AGEMA_signal_11602, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, new_AGEMA_signal_12766, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, new_AGEMA_signal_10252, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, new_AGEMA_signal_11605, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, new_AGEMA_signal_11608, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, new_AGEMA_signal_10969, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, new_AGEMA_signal_12157, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, new_AGEMA_signal_12769, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_12774, new_AGEMA_signal_12773, new_AGEMA_signal_12772, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, new_AGEMA_signal_10978, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, new_AGEMA_signal_12160, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, new_AGEMA_signal_11608, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, new_AGEMA_signal_12163, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, new_AGEMA_signal_11602, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, new_AGEMA_signal_12775, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, new_AGEMA_signal_12778, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, new_AGEMA_signal_12781, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_12786, new_AGEMA_signal_12785, new_AGEMA_signal_12784, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, new_AGEMA_signal_11599, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, new_AGEMA_signal_12787, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, new_AGEMA_signal_11605, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, new_AGEMA_signal_12790, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, new_AGEMA_signal_12775, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, new_AGEMA_signal_12766, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, new_AGEMA_signal_12781, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, new_AGEMA_signal_12157, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, new_AGEMA_signal_12787, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12774, new_AGEMA_signal_12773, new_AGEMA_signal_12772, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, new_AGEMA_signal_12769, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, new_AGEMA_signal_12160, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, new_AGEMA_signal_12778, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, new_AGEMA_signal_12790, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, new_AGEMA_signal_12763, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_12786, new_AGEMA_signal_12785, new_AGEMA_signal_12784, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, new_AGEMA_signal_12163, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_30592, new_AGEMA_signal_30589, new_AGEMA_signal_30586, new_AGEMA_signal_30583}), .clk (clk), .r ({Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220], Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216]}), .c ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_30604, new_AGEMA_signal_30601, new_AGEMA_signal_30598, new_AGEMA_signal_30595}), .clk (clk), .r ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230], Fresh[6229], Fresh[6228]}), .c ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, new_AGEMA_signal_10273, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_30616, new_AGEMA_signal_30613, new_AGEMA_signal_30610, new_AGEMA_signal_30607}), .clk (clk), .r ({Fresh[6251], Fresh[6250], Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .c ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_30628, new_AGEMA_signal_30625, new_AGEMA_signal_30622, new_AGEMA_signal_30619}), .clk (clk), .r ({Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260], Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252]}), .c ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, new_AGEMA_signal_10987, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_30640, new_AGEMA_signal_30637, new_AGEMA_signal_30634, new_AGEMA_signal_30631}), .clk (clk), .r ({Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270], Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264]}), .c ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_30652, new_AGEMA_signal_30649, new_AGEMA_signal_30646, new_AGEMA_signal_30643}), .clk (clk), .r ({Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280], Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276]}), .c ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_30664, new_AGEMA_signal_30661, new_AGEMA_signal_30658, new_AGEMA_signal_30655}), .clk (clk), .r ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290], Fresh[6289], Fresh[6288]}), .c ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_30676, new_AGEMA_signal_30673, new_AGEMA_signal_30670, new_AGEMA_signal_30667}), .clk (clk), .r ({Fresh[6311], Fresh[6310], Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .c ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_30688, new_AGEMA_signal_30685, new_AGEMA_signal_30682, new_AGEMA_signal_30679}), .clk (clk), .r ({Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320], Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312]}), .c ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, new_AGEMA_signal_10993, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_30700, new_AGEMA_signal_30697, new_AGEMA_signal_30694, new_AGEMA_signal_30691}), .clk (clk), .r ({Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330], Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324]}), .c ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_30712, new_AGEMA_signal_30709, new_AGEMA_signal_30706, new_AGEMA_signal_30703}), .clk (clk), .r ({Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340], Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336]}), .c ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_30724, new_AGEMA_signal_30721, new_AGEMA_signal_30718, new_AGEMA_signal_30715}), .clk (clk), .r ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350], Fresh[6349], Fresh[6348]}), .c ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, new_AGEMA_signal_10288, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_30736, new_AGEMA_signal_30733, new_AGEMA_signal_30730, new_AGEMA_signal_30727}), .clk (clk), .r ({Fresh[6371], Fresh[6370], Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .c ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_30748, new_AGEMA_signal_30745, new_AGEMA_signal_30742, new_AGEMA_signal_30739}), .clk (clk), .r ({Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380], Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372]}), .c ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, new_AGEMA_signal_10291, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_30760, new_AGEMA_signal_30757, new_AGEMA_signal_30754, new_AGEMA_signal_30751}), .clk (clk), .r ({Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390], Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384]}), .c ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, new_AGEMA_signal_10294, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_30772, new_AGEMA_signal_30769, new_AGEMA_signal_30766, new_AGEMA_signal_30763}), .clk (clk), .r ({Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400], Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396]}), .c ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_30784, new_AGEMA_signal_30781, new_AGEMA_signal_30778, new_AGEMA_signal_30775}), .clk (clk), .r ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410], Fresh[6409], Fresh[6408]}), .c ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_30796, new_AGEMA_signal_30793, new_AGEMA_signal_30790, new_AGEMA_signal_30787}), .clk (clk), .r ({Fresh[6431], Fresh[6430], Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .c ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, new_AGEMA_signal_11005, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, new_AGEMA_signal_10273, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, new_AGEMA_signal_10993, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, new_AGEMA_signal_10987, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, new_AGEMA_signal_11626, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, new_AGEMA_signal_11626, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, new_AGEMA_signal_10291, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, new_AGEMA_signal_10294, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, new_AGEMA_signal_11014, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_12798, new_AGEMA_signal_12797, new_AGEMA_signal_12796, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, new_AGEMA_signal_11629, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, new_AGEMA_signal_11632, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, new_AGEMA_signal_12799, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, new_AGEMA_signal_10288, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, new_AGEMA_signal_11635, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, new_AGEMA_signal_11638, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, new_AGEMA_signal_11005, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, new_AGEMA_signal_12184, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, new_AGEMA_signal_12802, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, new_AGEMA_signal_12805, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, new_AGEMA_signal_11014, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, new_AGEMA_signal_12187, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, new_AGEMA_signal_11638, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_12192, new_AGEMA_signal_12191, new_AGEMA_signal_12190, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, new_AGEMA_signal_11632, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_12810, new_AGEMA_signal_12809, new_AGEMA_signal_12808, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, new_AGEMA_signal_12811, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, new_AGEMA_signal_12814, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, new_AGEMA_signal_12817, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, new_AGEMA_signal_11629, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_12822, new_AGEMA_signal_12821, new_AGEMA_signal_12820, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, new_AGEMA_signal_11635, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, new_AGEMA_signal_12823, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12810, new_AGEMA_signal_12809, new_AGEMA_signal_12808, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, new_AGEMA_signal_12799, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, new_AGEMA_signal_12814, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, new_AGEMA_signal_12184, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_12822, new_AGEMA_signal_12821, new_AGEMA_signal_12820, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, new_AGEMA_signal_12805, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, new_AGEMA_signal_12802, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, new_AGEMA_signal_12187, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, new_AGEMA_signal_12811, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, new_AGEMA_signal_12823, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_12798, new_AGEMA_signal_12797, new_AGEMA_signal_12796, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, new_AGEMA_signal_12817, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12192, new_AGEMA_signal_12191, new_AGEMA_signal_12190, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_30808, new_AGEMA_signal_30805, new_AGEMA_signal_30802, new_AGEMA_signal_30799}), .clk (clk), .r ({Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440], Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432]}), .c ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_30820, new_AGEMA_signal_30817, new_AGEMA_signal_30814, new_AGEMA_signal_30811}), .clk (clk), .r ({Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450], Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444]}), .c ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, new_AGEMA_signal_10309, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_30832, new_AGEMA_signal_30829, new_AGEMA_signal_30826, new_AGEMA_signal_30823}), .clk (clk), .r ({Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460], Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456]}), .c ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_30844, new_AGEMA_signal_30841, new_AGEMA_signal_30838, new_AGEMA_signal_30835}), .clk (clk), .r ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470], Fresh[6469], Fresh[6468]}), .c ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, new_AGEMA_signal_11023, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_30856, new_AGEMA_signal_30853, new_AGEMA_signal_30850, new_AGEMA_signal_30847}), .clk (clk), .r ({Fresh[6491], Fresh[6490], Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .c ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_30868, new_AGEMA_signal_30865, new_AGEMA_signal_30862, new_AGEMA_signal_30859}), .clk (clk), .r ({Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500], Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492]}), .c ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_30880, new_AGEMA_signal_30877, new_AGEMA_signal_30874, new_AGEMA_signal_30871}), .clk (clk), .r ({Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510], Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504]}), .c ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_30892, new_AGEMA_signal_30889, new_AGEMA_signal_30886, new_AGEMA_signal_30883}), .clk (clk), .r ({Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520], Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516]}), .c ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_30904, new_AGEMA_signal_30901, new_AGEMA_signal_30898, new_AGEMA_signal_30895}), .clk (clk), .r ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530], Fresh[6529], Fresh[6528]}), .c ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, new_AGEMA_signal_11029, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_30916, new_AGEMA_signal_30913, new_AGEMA_signal_30910, new_AGEMA_signal_30907}), .clk (clk), .r ({Fresh[6551], Fresh[6550], Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .c ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_30928, new_AGEMA_signal_30925, new_AGEMA_signal_30922, new_AGEMA_signal_30919}), .clk (clk), .r ({Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560], Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552]}), .c ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_30940, new_AGEMA_signal_30937, new_AGEMA_signal_30934, new_AGEMA_signal_30931}), .clk (clk), .r ({Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570], Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564]}), .c ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, new_AGEMA_signal_10324, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_30952, new_AGEMA_signal_30949, new_AGEMA_signal_30946, new_AGEMA_signal_30943}), .clk (clk), .r ({Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580], Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576]}), .c ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_30964, new_AGEMA_signal_30961, new_AGEMA_signal_30958, new_AGEMA_signal_30955}), .clk (clk), .r ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590], Fresh[6589], Fresh[6588]}), .c ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, new_AGEMA_signal_10327, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_30976, new_AGEMA_signal_30973, new_AGEMA_signal_30970, new_AGEMA_signal_30967}), .clk (clk), .r ({Fresh[6611], Fresh[6610], Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .c ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, new_AGEMA_signal_10330, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_30988, new_AGEMA_signal_30985, new_AGEMA_signal_30982, new_AGEMA_signal_30979}), .clk (clk), .r ({Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620], Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612]}), .c ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_31000, new_AGEMA_signal_30997, new_AGEMA_signal_30994, new_AGEMA_signal_30991}), .clk (clk), .r ({Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630], Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624]}), .c ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_31012, new_AGEMA_signal_31009, new_AGEMA_signal_31006, new_AGEMA_signal_31003}), .clk (clk), .r ({Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640], Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636]}), .c ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, new_AGEMA_signal_11041, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, new_AGEMA_signal_10309, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, new_AGEMA_signal_11029, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, new_AGEMA_signal_11023, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_11658, new_AGEMA_signal_11657, new_AGEMA_signal_11656, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_11658, new_AGEMA_signal_11657, new_AGEMA_signal_11656, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, new_AGEMA_signal_10327, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, new_AGEMA_signal_10330, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, new_AGEMA_signal_11050, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, new_AGEMA_signal_12829, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, new_AGEMA_signal_11659, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, new_AGEMA_signal_11662, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_12834, new_AGEMA_signal_12833, new_AGEMA_signal_12832, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, new_AGEMA_signal_10324, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, new_AGEMA_signal_11665, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_11670, new_AGEMA_signal_11669, new_AGEMA_signal_11668, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, new_AGEMA_signal_11041, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, new_AGEMA_signal_12211, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, new_AGEMA_signal_12835, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, new_AGEMA_signal_12838, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, new_AGEMA_signal_11050, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, new_AGEMA_signal_12214, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_11670, new_AGEMA_signal_11669, new_AGEMA_signal_11668, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, new_AGEMA_signal_12217, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, new_AGEMA_signal_11662, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, new_AGEMA_signal_12841, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_12846, new_AGEMA_signal_12845, new_AGEMA_signal_12844, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, new_AGEMA_signal_12847, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, new_AGEMA_signal_12850, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, new_AGEMA_signal_11659, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, new_AGEMA_signal_12853, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, new_AGEMA_signal_11665, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_12858, new_AGEMA_signal_12857, new_AGEMA_signal_12856, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, new_AGEMA_signal_12841, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_12834, new_AGEMA_signal_12833, new_AGEMA_signal_12832, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, new_AGEMA_signal_12847, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, new_AGEMA_signal_12211, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, new_AGEMA_signal_12853, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, new_AGEMA_signal_12838, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, new_AGEMA_signal_12835, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, new_AGEMA_signal_12214, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_12846, new_AGEMA_signal_12845, new_AGEMA_signal_12844, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_12858, new_AGEMA_signal_12857, new_AGEMA_signal_12856, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, new_AGEMA_signal_12829, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, new_AGEMA_signal_12850, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, new_AGEMA_signal_12217, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_31024, new_AGEMA_signal_31021, new_AGEMA_signal_31018, new_AGEMA_signal_31015}), .clk (clk), .r ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650], Fresh[6649], Fresh[6648]}), .c ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_31036, new_AGEMA_signal_31033, new_AGEMA_signal_31030, new_AGEMA_signal_31027}), .clk (clk), .r ({Fresh[6671], Fresh[6670], Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .c ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, new_AGEMA_signal_10345, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_31048, new_AGEMA_signal_31045, new_AGEMA_signal_31042, new_AGEMA_signal_31039}), .clk (clk), .r ({Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680], Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672]}), .c ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_31060, new_AGEMA_signal_31057, new_AGEMA_signal_31054, new_AGEMA_signal_31051}), .clk (clk), .r ({Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690], Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684]}), .c ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, new_AGEMA_signal_11059, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_31072, new_AGEMA_signal_31069, new_AGEMA_signal_31066, new_AGEMA_signal_31063}), .clk (clk), .r ({Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700], Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696]}), .c ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_31084, new_AGEMA_signal_31081, new_AGEMA_signal_31078, new_AGEMA_signal_31075}), .clk (clk), .r ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710], Fresh[6709], Fresh[6708]}), .c ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_31096, new_AGEMA_signal_31093, new_AGEMA_signal_31090, new_AGEMA_signal_31087}), .clk (clk), .r ({Fresh[6731], Fresh[6730], Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720]}), .c ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_31108, new_AGEMA_signal_31105, new_AGEMA_signal_31102, new_AGEMA_signal_31099}), .clk (clk), .r ({Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740], Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732]}), .c ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_31120, new_AGEMA_signal_31117, new_AGEMA_signal_31114, new_AGEMA_signal_31111}), .clk (clk), .r ({Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750], Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744]}), .c ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, new_AGEMA_signal_11065, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_31132, new_AGEMA_signal_31129, new_AGEMA_signal_31126, new_AGEMA_signal_31123}), .clk (clk), .r ({Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760], Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756]}), .c ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_31144, new_AGEMA_signal_31141, new_AGEMA_signal_31138, new_AGEMA_signal_31135}), .clk (clk), .r ({Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770], Fresh[6769], Fresh[6768]}), .c ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_31156, new_AGEMA_signal_31153, new_AGEMA_signal_31150, new_AGEMA_signal_31147}), .clk (clk), .r ({Fresh[6791], Fresh[6790], Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780]}), .c ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, new_AGEMA_signal_10360, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_31168, new_AGEMA_signal_31165, new_AGEMA_signal_31162, new_AGEMA_signal_31159}), .clk (clk), .r ({Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800], Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792]}), .c ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_31180, new_AGEMA_signal_31177, new_AGEMA_signal_31174, new_AGEMA_signal_31171}), .clk (clk), .r ({Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810], Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804]}), .c ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, new_AGEMA_signal_10363, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_31192, new_AGEMA_signal_31189, new_AGEMA_signal_31186, new_AGEMA_signal_31183}), .clk (clk), .r ({Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820], Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816]}), .c ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, new_AGEMA_signal_10366, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_31204, new_AGEMA_signal_31201, new_AGEMA_signal_31198, new_AGEMA_signal_31195}), .clk (clk), .r ({Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830], Fresh[6829], Fresh[6828]}), .c ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_31216, new_AGEMA_signal_31213, new_AGEMA_signal_31210, new_AGEMA_signal_31207}), .clk (clk), .r ({Fresh[6851], Fresh[6850], Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840]}), .c ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_31228, new_AGEMA_signal_31225, new_AGEMA_signal_31222, new_AGEMA_signal_31219}), .clk (clk), .r ({Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860], Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852]}), .c ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, new_AGEMA_signal_11077, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, new_AGEMA_signal_10345, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, new_AGEMA_signal_11065, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, new_AGEMA_signal_11059, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, new_AGEMA_signal_11686, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, new_AGEMA_signal_11686, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, new_AGEMA_signal_10363, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, new_AGEMA_signal_10366, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, new_AGEMA_signal_11086, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_12864, new_AGEMA_signal_12863, new_AGEMA_signal_12862, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, new_AGEMA_signal_11689, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_11694, new_AGEMA_signal_11693, new_AGEMA_signal_11692, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, new_AGEMA_signal_12865, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, new_AGEMA_signal_10360, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, new_AGEMA_signal_11695, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, new_AGEMA_signal_11698, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, new_AGEMA_signal_11077, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, new_AGEMA_signal_12238, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_12870, new_AGEMA_signal_12869, new_AGEMA_signal_12868, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, new_AGEMA_signal_12871, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, new_AGEMA_signal_11086, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, new_AGEMA_signal_12241, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, new_AGEMA_signal_11698, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, new_AGEMA_signal_12244, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_11694, new_AGEMA_signal_11693, new_AGEMA_signal_11692, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_12876, new_AGEMA_signal_12875, new_AGEMA_signal_12874, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, new_AGEMA_signal_12877, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_12882, new_AGEMA_signal_12881, new_AGEMA_signal_12880, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, new_AGEMA_signal_12883, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, new_AGEMA_signal_11689, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_12888, new_AGEMA_signal_12887, new_AGEMA_signal_12886, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, new_AGEMA_signal_11695, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, new_AGEMA_signal_12889, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12876, new_AGEMA_signal_12875, new_AGEMA_signal_12874, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, new_AGEMA_signal_12865, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_12882, new_AGEMA_signal_12881, new_AGEMA_signal_12880, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, new_AGEMA_signal_12238, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_12888, new_AGEMA_signal_12887, new_AGEMA_signal_12886, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, new_AGEMA_signal_12871, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_12870, new_AGEMA_signal_12869, new_AGEMA_signal_12868, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, new_AGEMA_signal_12241, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, new_AGEMA_signal_12877, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, new_AGEMA_signal_12889, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_12864, new_AGEMA_signal_12863, new_AGEMA_signal_12862, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, new_AGEMA_signal_12883, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, new_AGEMA_signal_12244, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_31240, new_AGEMA_signal_31237, new_AGEMA_signal_31234, new_AGEMA_signal_31231}), .clk (clk), .r ({Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870], Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864]}), .c ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_31252, new_AGEMA_signal_31249, new_AGEMA_signal_31246, new_AGEMA_signal_31243}), .clk (clk), .r ({Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880], Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876]}), .c ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, new_AGEMA_signal_10381, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_31264, new_AGEMA_signal_31261, new_AGEMA_signal_31258, new_AGEMA_signal_31255}), .clk (clk), .r ({Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890], Fresh[6889], Fresh[6888]}), .c ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_31276, new_AGEMA_signal_31273, new_AGEMA_signal_31270, new_AGEMA_signal_31267}), .clk (clk), .r ({Fresh[6911], Fresh[6910], Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900]}), .c ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, new_AGEMA_signal_11095, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_31288, new_AGEMA_signal_31285, new_AGEMA_signal_31282, new_AGEMA_signal_31279}), .clk (clk), .r ({Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920], Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912]}), .c ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_31300, new_AGEMA_signal_31297, new_AGEMA_signal_31294, new_AGEMA_signal_31291}), .clk (clk), .r ({Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930], Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924]}), .c ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_31312, new_AGEMA_signal_31309, new_AGEMA_signal_31306, new_AGEMA_signal_31303}), .clk (clk), .r ({Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940], Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936]}), .c ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_31324, new_AGEMA_signal_31321, new_AGEMA_signal_31318, new_AGEMA_signal_31315}), .clk (clk), .r ({Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950], Fresh[6949], Fresh[6948]}), .c ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_31336, new_AGEMA_signal_31333, new_AGEMA_signal_31330, new_AGEMA_signal_31327}), .clk (clk), .r ({Fresh[6971], Fresh[6970], Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960]}), .c ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, new_AGEMA_signal_11101, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_31348, new_AGEMA_signal_31345, new_AGEMA_signal_31342, new_AGEMA_signal_31339}), .clk (clk), .r ({Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980], Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972]}), .c ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_31360, new_AGEMA_signal_31357, new_AGEMA_signal_31354, new_AGEMA_signal_31351}), .clk (clk), .r ({Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990], Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984]}), .c ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_31372, new_AGEMA_signal_31369, new_AGEMA_signal_31366, new_AGEMA_signal_31363}), .clk (clk), .r ({Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000], Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996]}), .c ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, new_AGEMA_signal_10396, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_31384, new_AGEMA_signal_31381, new_AGEMA_signal_31378, new_AGEMA_signal_31375}), .clk (clk), .r ({Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010], Fresh[7009], Fresh[7008]}), .c ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_31396, new_AGEMA_signal_31393, new_AGEMA_signal_31390, new_AGEMA_signal_31387}), .clk (clk), .r ({Fresh[7031], Fresh[7030], Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020]}), .c ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, new_AGEMA_signal_10399, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_31408, new_AGEMA_signal_31405, new_AGEMA_signal_31402, new_AGEMA_signal_31399}), .clk (clk), .r ({Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040], Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032]}), .c ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, new_AGEMA_signal_10402, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_31420, new_AGEMA_signal_31417, new_AGEMA_signal_31414, new_AGEMA_signal_31411}), .clk (clk), .r ({Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050], Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044]}), .c ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_31432, new_AGEMA_signal_31429, new_AGEMA_signal_31426, new_AGEMA_signal_31423}), .clk (clk), .r ({Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060], Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056]}), .c ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_31444, new_AGEMA_signal_31441, new_AGEMA_signal_31438, new_AGEMA_signal_31435}), .clk (clk), .r ({Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070], Fresh[7069], Fresh[7068]}), .c ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, new_AGEMA_signal_11113, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, new_AGEMA_signal_10381, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, new_AGEMA_signal_11101, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, new_AGEMA_signal_11095, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_11718, new_AGEMA_signal_11717, new_AGEMA_signal_11716, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_11718, new_AGEMA_signal_11717, new_AGEMA_signal_11716, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, new_AGEMA_signal_10399, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, new_AGEMA_signal_10402, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, new_AGEMA_signal_11122, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, new_AGEMA_signal_12895, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, new_AGEMA_signal_11719, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, new_AGEMA_signal_11722, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_12900, new_AGEMA_signal_12899, new_AGEMA_signal_12898, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, new_AGEMA_signal_10396, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, new_AGEMA_signal_11725, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_11730, new_AGEMA_signal_11729, new_AGEMA_signal_11728, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, new_AGEMA_signal_11113, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, new_AGEMA_signal_12265, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, new_AGEMA_signal_12901, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_12906, new_AGEMA_signal_12905, new_AGEMA_signal_12904, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, new_AGEMA_signal_11122, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, new_AGEMA_signal_12268, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_11730, new_AGEMA_signal_11729, new_AGEMA_signal_11728, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, new_AGEMA_signal_12271, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, new_AGEMA_signal_11722, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, new_AGEMA_signal_12907, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_12912, new_AGEMA_signal_12911, new_AGEMA_signal_12910, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, new_AGEMA_signal_12913, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_12918, new_AGEMA_signal_12917, new_AGEMA_signal_12916, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, new_AGEMA_signal_11719, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, new_AGEMA_signal_12919, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, new_AGEMA_signal_11725, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_12924, new_AGEMA_signal_12923, new_AGEMA_signal_12922, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, new_AGEMA_signal_12907, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_12900, new_AGEMA_signal_12899, new_AGEMA_signal_12898, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, new_AGEMA_signal_12913, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, new_AGEMA_signal_12265, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, new_AGEMA_signal_12919, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12906, new_AGEMA_signal_12905, new_AGEMA_signal_12904, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, new_AGEMA_signal_12901, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, new_AGEMA_signal_12268, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_12912, new_AGEMA_signal_12911, new_AGEMA_signal_12910, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_12924, new_AGEMA_signal_12923, new_AGEMA_signal_12922, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, new_AGEMA_signal_12895, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_12918, new_AGEMA_signal_12917, new_AGEMA_signal_12916, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, new_AGEMA_signal_12271, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_31456, new_AGEMA_signal_31453, new_AGEMA_signal_31450, new_AGEMA_signal_31447}), .clk (clk), .r ({Fresh[7091], Fresh[7090], Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080]}), .c ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_31468, new_AGEMA_signal_31465, new_AGEMA_signal_31462, new_AGEMA_signal_31459}), .clk (clk), .r ({Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100], Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092]}), .c ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, new_AGEMA_signal_10417, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_31480, new_AGEMA_signal_31477, new_AGEMA_signal_31474, new_AGEMA_signal_31471}), .clk (clk), .r ({Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110], Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104]}), .c ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_31492, new_AGEMA_signal_31489, new_AGEMA_signal_31486, new_AGEMA_signal_31483}), .clk (clk), .r ({Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120], Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116]}), .c ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, new_AGEMA_signal_11131, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_31504, new_AGEMA_signal_31501, new_AGEMA_signal_31498, new_AGEMA_signal_31495}), .clk (clk), .r ({Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130], Fresh[7129], Fresh[7128]}), .c ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_31516, new_AGEMA_signal_31513, new_AGEMA_signal_31510, new_AGEMA_signal_31507}), .clk (clk), .r ({Fresh[7151], Fresh[7150], Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140]}), .c ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_31528, new_AGEMA_signal_31525, new_AGEMA_signal_31522, new_AGEMA_signal_31519}), .clk (clk), .r ({Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160], Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152]}), .c ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_31540, new_AGEMA_signal_31537, new_AGEMA_signal_31534, new_AGEMA_signal_31531}), .clk (clk), .r ({Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170], Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164]}), .c ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_31552, new_AGEMA_signal_31549, new_AGEMA_signal_31546, new_AGEMA_signal_31543}), .clk (clk), .r ({Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180], Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176]}), .c ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, new_AGEMA_signal_11137, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_31564, new_AGEMA_signal_31561, new_AGEMA_signal_31558, new_AGEMA_signal_31555}), .clk (clk), .r ({Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190], Fresh[7189], Fresh[7188]}), .c ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_31576, new_AGEMA_signal_31573, new_AGEMA_signal_31570, new_AGEMA_signal_31567}), .clk (clk), .r ({Fresh[7211], Fresh[7210], Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200]}), .c ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_31588, new_AGEMA_signal_31585, new_AGEMA_signal_31582, new_AGEMA_signal_31579}), .clk (clk), .r ({Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220], Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212]}), .c ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, new_AGEMA_signal_10432, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_31600, new_AGEMA_signal_31597, new_AGEMA_signal_31594, new_AGEMA_signal_31591}), .clk (clk), .r ({Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230], Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224]}), .c ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_31612, new_AGEMA_signal_31609, new_AGEMA_signal_31606, new_AGEMA_signal_31603}), .clk (clk), .r ({Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240], Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236]}), .c ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, new_AGEMA_signal_10435, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_31624, new_AGEMA_signal_31621, new_AGEMA_signal_31618, new_AGEMA_signal_31615}), .clk (clk), .r ({Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250], Fresh[7249], Fresh[7248]}), .c ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, new_AGEMA_signal_10438, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_31636, new_AGEMA_signal_31633, new_AGEMA_signal_31630, new_AGEMA_signal_31627}), .clk (clk), .r ({Fresh[7271], Fresh[7270], Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260]}), .c ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_31648, new_AGEMA_signal_31645, new_AGEMA_signal_31642, new_AGEMA_signal_31639}), .clk (clk), .r ({Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280], Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272]}), .c ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_31660, new_AGEMA_signal_31657, new_AGEMA_signal_31654, new_AGEMA_signal_31651}), .clk (clk), .r ({Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290], Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284]}), .c ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, new_AGEMA_signal_11149, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, new_AGEMA_signal_10417, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, new_AGEMA_signal_11137, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, new_AGEMA_signal_11131, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, new_AGEMA_signal_11746, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, new_AGEMA_signal_11746, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, new_AGEMA_signal_10435, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, new_AGEMA_signal_10438, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, new_AGEMA_signal_11158, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_12930, new_AGEMA_signal_12929, new_AGEMA_signal_12928, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, new_AGEMA_signal_11749, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_11754, new_AGEMA_signal_11753, new_AGEMA_signal_11752, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, new_AGEMA_signal_12931, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, new_AGEMA_signal_10432, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, new_AGEMA_signal_11755, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, new_AGEMA_signal_11758, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, new_AGEMA_signal_11149, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, new_AGEMA_signal_12292, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_12936, new_AGEMA_signal_12935, new_AGEMA_signal_12934, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, new_AGEMA_signal_12937, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, new_AGEMA_signal_11158, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, new_AGEMA_signal_12295, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, new_AGEMA_signal_11758, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, new_AGEMA_signal_12298, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_11754, new_AGEMA_signal_11753, new_AGEMA_signal_11752, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_12942, new_AGEMA_signal_12941, new_AGEMA_signal_12940, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, new_AGEMA_signal_12943, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_12948, new_AGEMA_signal_12947, new_AGEMA_signal_12946, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, new_AGEMA_signal_12949, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, new_AGEMA_signal_11749, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_12954, new_AGEMA_signal_12953, new_AGEMA_signal_12952, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, new_AGEMA_signal_11755, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, new_AGEMA_signal_12955, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12942, new_AGEMA_signal_12941, new_AGEMA_signal_12940, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, new_AGEMA_signal_12931, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_12948, new_AGEMA_signal_12947, new_AGEMA_signal_12946, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, new_AGEMA_signal_12292, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_12954, new_AGEMA_signal_12953, new_AGEMA_signal_12952, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, new_AGEMA_signal_12937, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_12936, new_AGEMA_signal_12935, new_AGEMA_signal_12934, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, new_AGEMA_signal_12295, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, new_AGEMA_signal_12943, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, new_AGEMA_signal_12955, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_12930, new_AGEMA_signal_12929, new_AGEMA_signal_12928, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, new_AGEMA_signal_12949, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, new_AGEMA_signal_12298, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_14811, new_AGEMA_signal_14810, new_AGEMA_signal_14809, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_15714, new_AGEMA_signal_15713, new_AGEMA_signal_15712, MixColumnsOutput[105]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_14811, new_AGEMA_signal_14810, new_AGEMA_signal_14809, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, new_AGEMA_signal_14137, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_14814, new_AGEMA_signal_14813, new_AGEMA_signal_14812, MixColumnsOutput[104]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .c ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, new_AGEMA_signal_14137, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_14142, new_AGEMA_signal_14141, new_AGEMA_signal_14140, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_14817, new_AGEMA_signal_14816, new_AGEMA_signal_14815, MixColumnsOutput[103]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_14142, new_AGEMA_signal_14141, new_AGEMA_signal_14140, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, new_AGEMA_signal_14143, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_14820, new_AGEMA_signal_14819, new_AGEMA_signal_14818, MixColumnsOutput[102]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, new_AGEMA_signal_14143, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_14148, new_AGEMA_signal_14147, new_AGEMA_signal_14146, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_14823, new_AGEMA_signal_14822, new_AGEMA_signal_14821, MixColumnsOutput[101]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_14148, new_AGEMA_signal_14147, new_AGEMA_signal_14146, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_14826, new_AGEMA_signal_14825, new_AGEMA_signal_14824, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, new_AGEMA_signal_15715, MixColumnsOutput[100]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_14826, new_AGEMA_signal_14825, new_AGEMA_signal_14824, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, new_AGEMA_signal_14827, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_15720, new_AGEMA_signal_15719, new_AGEMA_signal_15718, MixColumnsOutput[99]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .c ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, new_AGEMA_signal_14827, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, new_AGEMA_signal_14149, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_14832, new_AGEMA_signal_14831, new_AGEMA_signal_14830, MixColumnsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, new_AGEMA_signal_14149, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_14154, new_AGEMA_signal_14153, new_AGEMA_signal_14152, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, new_AGEMA_signal_14833, MixColumnsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_14154, new_AGEMA_signal_14153, new_AGEMA_signal_14152, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, new_AGEMA_signal_14155, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_14838, new_AGEMA_signal_14837, new_AGEMA_signal_14836, MixColumnsOutput[98]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .c ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, new_AGEMA_signal_14155, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_14160, new_AGEMA_signal_14159, new_AGEMA_signal_14158, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, new_AGEMA_signal_14839, MixColumnsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_14160, new_AGEMA_signal_14159, new_AGEMA_signal_14158, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_14844, new_AGEMA_signal_14843, new_AGEMA_signal_14842, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, new_AGEMA_signal_15721, MixColumnsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, new_AGEMA_signal_13567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_14844, new_AGEMA_signal_14843, new_AGEMA_signal_14842, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, new_AGEMA_signal_14845, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_15726, new_AGEMA_signal_15725, new_AGEMA_signal_15724, MixColumnsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .b ({new_AGEMA_signal_13572, new_AGEMA_signal_13571, new_AGEMA_signal_13570, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .b ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, new_AGEMA_signal_14845, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, new_AGEMA_signal_14167, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_14850, new_AGEMA_signal_14849, new_AGEMA_signal_14848, MixColumnsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .b ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, new_AGEMA_signal_14167, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, new_AGEMA_signal_14851, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_15729, new_AGEMA_signal_15728, new_AGEMA_signal_15727, MixColumnsOutput[121]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, new_AGEMA_signal_14851, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_14172, new_AGEMA_signal_14171, new_AGEMA_signal_14170, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_14856, new_AGEMA_signal_14855, new_AGEMA_signal_14854, MixColumnsOutput[120]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_14172, new_AGEMA_signal_14171, new_AGEMA_signal_14170, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, new_AGEMA_signal_14173, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, new_AGEMA_signal_14857, MixColumnsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, new_AGEMA_signal_14173, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_14178, new_AGEMA_signal_14177, new_AGEMA_signal_14176, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_14862, new_AGEMA_signal_14861, new_AGEMA_signal_14860, MixColumnsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_14178, new_AGEMA_signal_14177, new_AGEMA_signal_14176, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, new_AGEMA_signal_14179, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_14865, new_AGEMA_signal_14864, new_AGEMA_signal_14863, MixColumnsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, new_AGEMA_signal_14179, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_14868, new_AGEMA_signal_14867, new_AGEMA_signal_14866, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_15732, new_AGEMA_signal_15731, new_AGEMA_signal_15730, MixColumnsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_13578, new_AGEMA_signal_13577, new_AGEMA_signal_13576, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_14868, new_AGEMA_signal_14867, new_AGEMA_signal_14866, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_14871, new_AGEMA_signal_14870, new_AGEMA_signal_14869, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_15735, new_AGEMA_signal_15734, new_AGEMA_signal_15733, MixColumnsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, new_AGEMA_signal_13573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_14871, new_AGEMA_signal_14870, new_AGEMA_signal_14869, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_13602, new_AGEMA_signal_13601, new_AGEMA_signal_13600, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_14874, new_AGEMA_signal_14873, new_AGEMA_signal_14872, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_15738, new_AGEMA_signal_15737, new_AGEMA_signal_15736, MixColumnsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .b ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, new_AGEMA_signal_13579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .b ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_14874, new_AGEMA_signal_14873, new_AGEMA_signal_14872, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_14196, new_AGEMA_signal_14195, new_AGEMA_signal_14194, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_14877, new_AGEMA_signal_14876, new_AGEMA_signal_14875, MixColumnsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .b ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_14196, new_AGEMA_signal_14195, new_AGEMA_signal_14194, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_14880, new_AGEMA_signal_14879, new_AGEMA_signal_14878, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, new_AGEMA_signal_15739, MixColumnsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_13584, new_AGEMA_signal_13583, new_AGEMA_signal_13582, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_14880, new_AGEMA_signal_14879, new_AGEMA_signal_14878, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, new_AGEMA_signal_13591, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, new_AGEMA_signal_14203, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_14883, new_AGEMA_signal_14882, new_AGEMA_signal_14881, MixColumnsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .b ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, new_AGEMA_signal_14203, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_14208, new_AGEMA_signal_14207, new_AGEMA_signal_14206, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_14886, new_AGEMA_signal_14885, new_AGEMA_signal_14884, MixColumnsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_14208, new_AGEMA_signal_14207, new_AGEMA_signal_14206, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, new_AGEMA_signal_14209, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_14889, new_AGEMA_signal_14888, new_AGEMA_signal_14887, MixColumnsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, new_AGEMA_signal_14209, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_14214, new_AGEMA_signal_14213, new_AGEMA_signal_14212, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_14892, new_AGEMA_signal_14891, new_AGEMA_signal_14890, MixColumnsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_14214, new_AGEMA_signal_14213, new_AGEMA_signal_14212, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_14895, new_AGEMA_signal_14894, new_AGEMA_signal_14893, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_15744, new_AGEMA_signal_15743, new_AGEMA_signal_15742, MixColumnsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, new_AGEMA_signal_13585, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_14895, new_AGEMA_signal_14894, new_AGEMA_signal_14893, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_13596, new_AGEMA_signal_13595, new_AGEMA_signal_13594, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_14898, new_AGEMA_signal_14897, new_AGEMA_signal_14896, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, new_AGEMA_signal_15745, MixColumnsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .b ({new_AGEMA_signal_13590, new_AGEMA_signal_13589, new_AGEMA_signal_13588, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .c ({new_AGEMA_signal_14898, new_AGEMA_signal_14897, new_AGEMA_signal_14896, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, new_AGEMA_signal_13597, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .c ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, new_AGEMA_signal_14227, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, new_AGEMA_signal_14899, MixColumnsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .c ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, new_AGEMA_signal_14227, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .c ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_14232, new_AGEMA_signal_14231, new_AGEMA_signal_14230, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .c ({new_AGEMA_signal_14904, new_AGEMA_signal_14903, new_AGEMA_signal_14902, MixColumnsOutput[96]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_14232, new_AGEMA_signal_14231, new_AGEMA_signal_14230, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .c ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .c ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, new_AGEMA_signal_13567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .c ({new_AGEMA_signal_13572, new_AGEMA_signal_13571, new_AGEMA_signal_13570, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .c ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, new_AGEMA_signal_13573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .c ({new_AGEMA_signal_13578, new_AGEMA_signal_13577, new_AGEMA_signal_13576, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .c ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, new_AGEMA_signal_13579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .c ({new_AGEMA_signal_13584, new_AGEMA_signal_13583, new_AGEMA_signal_13582, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .c ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, new_AGEMA_signal_13585, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .c ({new_AGEMA_signal_13590, new_AGEMA_signal_13589, new_AGEMA_signal_13588, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .c ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, new_AGEMA_signal_13591, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .c ({new_AGEMA_signal_13596, new_AGEMA_signal_13595, new_AGEMA_signal_13594, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .c ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, new_AGEMA_signal_13597, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_13602, new_AGEMA_signal_13601, new_AGEMA_signal_13600, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_14907, new_AGEMA_signal_14906, new_AGEMA_signal_14905, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_15750, new_AGEMA_signal_15749, new_AGEMA_signal_15748, MixColumnsOutput[73]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_14907, new_AGEMA_signal_14906, new_AGEMA_signal_14905, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, new_AGEMA_signal_14233, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_14910, new_AGEMA_signal_14909, new_AGEMA_signal_14908, MixColumnsOutput[72]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .c ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, new_AGEMA_signal_14233, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_14238, new_AGEMA_signal_14237, new_AGEMA_signal_14236, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, new_AGEMA_signal_14911, MixColumnsOutput[71]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_14238, new_AGEMA_signal_14237, new_AGEMA_signal_14236, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, new_AGEMA_signal_14239, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_14916, new_AGEMA_signal_14915, new_AGEMA_signal_14914, MixColumnsOutput[70]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, new_AGEMA_signal_14239, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_14244, new_AGEMA_signal_14243, new_AGEMA_signal_14242, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, new_AGEMA_signal_14917, MixColumnsOutput[69]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_14244, new_AGEMA_signal_14243, new_AGEMA_signal_14242, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_14922, new_AGEMA_signal_14921, new_AGEMA_signal_14920, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_15753, new_AGEMA_signal_15752, new_AGEMA_signal_15751, MixColumnsOutput[68]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_14922, new_AGEMA_signal_14921, new_AGEMA_signal_14920, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, new_AGEMA_signal_14923, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_15756, new_AGEMA_signal_15755, new_AGEMA_signal_15754, MixColumnsOutput[67]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .c ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, new_AGEMA_signal_14923, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, new_AGEMA_signal_14245, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_14928, new_AGEMA_signal_14927, new_AGEMA_signal_14926, MixColumnsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, new_AGEMA_signal_14245, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_14250, new_AGEMA_signal_14249, new_AGEMA_signal_14248, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, new_AGEMA_signal_14929, MixColumnsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_14250, new_AGEMA_signal_14249, new_AGEMA_signal_14248, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, new_AGEMA_signal_14251, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_14934, new_AGEMA_signal_14933, new_AGEMA_signal_14932, MixColumnsOutput[66]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .c ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, new_AGEMA_signal_14251, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_14256, new_AGEMA_signal_14255, new_AGEMA_signal_14254, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_14937, new_AGEMA_signal_14936, new_AGEMA_signal_14935, MixColumnsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_14256, new_AGEMA_signal_14255, new_AGEMA_signal_14254, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_14940, new_AGEMA_signal_14939, new_AGEMA_signal_14938, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, new_AGEMA_signal_15757, MixColumnsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, new_AGEMA_signal_13663, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_14940, new_AGEMA_signal_14939, new_AGEMA_signal_14938, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_14943, new_AGEMA_signal_14942, new_AGEMA_signal_14941, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_15762, new_AGEMA_signal_15761, new_AGEMA_signal_15760, MixColumnsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .b ({new_AGEMA_signal_13668, new_AGEMA_signal_13667, new_AGEMA_signal_13666, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .b ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_14943, new_AGEMA_signal_14942, new_AGEMA_signal_14941, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, new_AGEMA_signal_14263, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_14946, new_AGEMA_signal_14945, new_AGEMA_signal_14944, MixColumnsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .b ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, new_AGEMA_signal_14263, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_14949, new_AGEMA_signal_14948, new_AGEMA_signal_14947, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_15765, new_AGEMA_signal_15764, new_AGEMA_signal_15763, MixColumnsOutput[89]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_14949, new_AGEMA_signal_14948, new_AGEMA_signal_14947, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_14268, new_AGEMA_signal_14267, new_AGEMA_signal_14266, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_14952, new_AGEMA_signal_14951, new_AGEMA_signal_14950, MixColumnsOutput[88]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_14268, new_AGEMA_signal_14267, new_AGEMA_signal_14266, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, new_AGEMA_signal_14269, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, new_AGEMA_signal_14953, MixColumnsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, new_AGEMA_signal_14269, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_14274, new_AGEMA_signal_14273, new_AGEMA_signal_14272, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_14958, new_AGEMA_signal_14957, new_AGEMA_signal_14956, MixColumnsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_14274, new_AGEMA_signal_14273, new_AGEMA_signal_14272, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, new_AGEMA_signal_14275, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, new_AGEMA_signal_14959, MixColumnsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, new_AGEMA_signal_14275, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_14964, new_AGEMA_signal_14963, new_AGEMA_signal_14962, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_15768, new_AGEMA_signal_15767, new_AGEMA_signal_15766, MixColumnsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_13674, new_AGEMA_signal_13673, new_AGEMA_signal_13672, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_14964, new_AGEMA_signal_14963, new_AGEMA_signal_14962, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, new_AGEMA_signal_14965, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_15771, new_AGEMA_signal_15770, new_AGEMA_signal_15769, MixColumnsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, new_AGEMA_signal_13669, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, new_AGEMA_signal_14965, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_13698, new_AGEMA_signal_13697, new_AGEMA_signal_13696, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_14970, new_AGEMA_signal_14969, new_AGEMA_signal_14968, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_15774, new_AGEMA_signal_15773, new_AGEMA_signal_15772, MixColumnsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .b ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, new_AGEMA_signal_13675, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .b ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_14970, new_AGEMA_signal_14969, new_AGEMA_signal_14968, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_14292, new_AGEMA_signal_14291, new_AGEMA_signal_14290, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, new_AGEMA_signal_14971, MixColumnsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .b ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_14292, new_AGEMA_signal_14291, new_AGEMA_signal_14290, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_14976, new_AGEMA_signal_14975, new_AGEMA_signal_14974, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_15777, new_AGEMA_signal_15776, new_AGEMA_signal_15775, MixColumnsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_13680, new_AGEMA_signal_13679, new_AGEMA_signal_13678, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_14976, new_AGEMA_signal_14975, new_AGEMA_signal_14974, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, new_AGEMA_signal_13687, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, new_AGEMA_signal_14299, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, new_AGEMA_signal_14977, MixColumnsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .b ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, new_AGEMA_signal_14299, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_14304, new_AGEMA_signal_14303, new_AGEMA_signal_14302, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_14982, new_AGEMA_signal_14981, new_AGEMA_signal_14980, MixColumnsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_14304, new_AGEMA_signal_14303, new_AGEMA_signal_14302, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, new_AGEMA_signal_14305, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_14985, new_AGEMA_signal_14984, new_AGEMA_signal_14983, MixColumnsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, new_AGEMA_signal_14305, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_14310, new_AGEMA_signal_14309, new_AGEMA_signal_14308, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_14988, new_AGEMA_signal_14987, new_AGEMA_signal_14986, MixColumnsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_14310, new_AGEMA_signal_14309, new_AGEMA_signal_14308, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_14991, new_AGEMA_signal_14990, new_AGEMA_signal_14989, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_15780, new_AGEMA_signal_15779, new_AGEMA_signal_15778, MixColumnsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, new_AGEMA_signal_13681, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_14991, new_AGEMA_signal_14990, new_AGEMA_signal_14989, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_13692, new_AGEMA_signal_13691, new_AGEMA_signal_13690, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_14994, new_AGEMA_signal_14993, new_AGEMA_signal_14992, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_15783, new_AGEMA_signal_15782, new_AGEMA_signal_15781, MixColumnsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .b ({new_AGEMA_signal_13686, new_AGEMA_signal_13685, new_AGEMA_signal_13684, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .c ({new_AGEMA_signal_14994, new_AGEMA_signal_14993, new_AGEMA_signal_14992, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, new_AGEMA_signal_13693, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .c ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, new_AGEMA_signal_14323, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, new_AGEMA_signal_14995, MixColumnsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .c ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, new_AGEMA_signal_14323, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .c ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_14328, new_AGEMA_signal_14327, new_AGEMA_signal_14326, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .c ({new_AGEMA_signal_15000, new_AGEMA_signal_14999, new_AGEMA_signal_14998, MixColumnsOutput[64]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_14328, new_AGEMA_signal_14327, new_AGEMA_signal_14326, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .c ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .c ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, new_AGEMA_signal_13663, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .c ({new_AGEMA_signal_13668, new_AGEMA_signal_13667, new_AGEMA_signal_13666, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .c ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, new_AGEMA_signal_13669, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .c ({new_AGEMA_signal_13674, new_AGEMA_signal_13673, new_AGEMA_signal_13672, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .c ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, new_AGEMA_signal_13675, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .c ({new_AGEMA_signal_13680, new_AGEMA_signal_13679, new_AGEMA_signal_13678, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .c ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, new_AGEMA_signal_13681, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .c ({new_AGEMA_signal_13686, new_AGEMA_signal_13685, new_AGEMA_signal_13684, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .c ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, new_AGEMA_signal_13687, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .c ({new_AGEMA_signal_13692, new_AGEMA_signal_13691, new_AGEMA_signal_13690, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .c ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, new_AGEMA_signal_13693, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_13698, new_AGEMA_signal_13697, new_AGEMA_signal_13696, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, new_AGEMA_signal_15001, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_15786, new_AGEMA_signal_15785, new_AGEMA_signal_15784, MixColumnsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, new_AGEMA_signal_15001, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, new_AGEMA_signal_14329, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_15006, new_AGEMA_signal_15005, new_AGEMA_signal_15004, MixColumnsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .c ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, new_AGEMA_signal_14329, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_14334, new_AGEMA_signal_14333, new_AGEMA_signal_14332, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, new_AGEMA_signal_15007, MixColumnsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_14334, new_AGEMA_signal_14333, new_AGEMA_signal_14332, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, new_AGEMA_signal_14335, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_15012, new_AGEMA_signal_15011, new_AGEMA_signal_15010, MixColumnsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, new_AGEMA_signal_14335, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_14340, new_AGEMA_signal_14339, new_AGEMA_signal_14338, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, new_AGEMA_signal_15013, MixColumnsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_14340, new_AGEMA_signal_14339, new_AGEMA_signal_14338, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_15018, new_AGEMA_signal_15017, new_AGEMA_signal_15016, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_15789, new_AGEMA_signal_15788, new_AGEMA_signal_15787, MixColumnsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_15018, new_AGEMA_signal_15017, new_AGEMA_signal_15016, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, new_AGEMA_signal_15019, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_15792, new_AGEMA_signal_15791, new_AGEMA_signal_15790, MixColumnsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .c ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, new_AGEMA_signal_15019, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, new_AGEMA_signal_14341, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_15024, new_AGEMA_signal_15023, new_AGEMA_signal_15022, MixColumnsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, new_AGEMA_signal_14341, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_14346, new_AGEMA_signal_14345, new_AGEMA_signal_14344, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, new_AGEMA_signal_15025, MixColumnsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_14346, new_AGEMA_signal_14345, new_AGEMA_signal_14344, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, new_AGEMA_signal_14347, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_15030, new_AGEMA_signal_15029, new_AGEMA_signal_15028, MixColumnsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .c ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, new_AGEMA_signal_14347, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_14352, new_AGEMA_signal_14351, new_AGEMA_signal_14350, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, new_AGEMA_signal_15031, MixColumnsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_14352, new_AGEMA_signal_14351, new_AGEMA_signal_14350, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_15036, new_AGEMA_signal_15035, new_AGEMA_signal_15034, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_15795, new_AGEMA_signal_15794, new_AGEMA_signal_15793, MixColumnsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, new_AGEMA_signal_13759, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_15036, new_AGEMA_signal_15035, new_AGEMA_signal_15034, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_15039, new_AGEMA_signal_15038, new_AGEMA_signal_15037, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_15798, new_AGEMA_signal_15797, new_AGEMA_signal_15796, MixColumnsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .b ({new_AGEMA_signal_13764, new_AGEMA_signal_13763, new_AGEMA_signal_13762, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .b ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_15039, new_AGEMA_signal_15038, new_AGEMA_signal_15037, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, new_AGEMA_signal_14359, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_15042, new_AGEMA_signal_15041, new_AGEMA_signal_15040, MixColumnsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .b ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, new_AGEMA_signal_14359, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, new_AGEMA_signal_15043, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, new_AGEMA_signal_15799, MixColumnsOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, new_AGEMA_signal_15043, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_14364, new_AGEMA_signal_14363, new_AGEMA_signal_14362, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_15048, new_AGEMA_signal_15047, new_AGEMA_signal_15046, MixColumnsOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_14364, new_AGEMA_signal_14363, new_AGEMA_signal_14362, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, new_AGEMA_signal_14365, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, new_AGEMA_signal_15049, MixColumnsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, new_AGEMA_signal_14365, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_14370, new_AGEMA_signal_14369, new_AGEMA_signal_14368, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_15054, new_AGEMA_signal_15053, new_AGEMA_signal_15052, MixColumnsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_14370, new_AGEMA_signal_14369, new_AGEMA_signal_14368, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, new_AGEMA_signal_14371, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, new_AGEMA_signal_15055, MixColumnsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, new_AGEMA_signal_14371, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_15060, new_AGEMA_signal_15059, new_AGEMA_signal_15058, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_15804, new_AGEMA_signal_15803, new_AGEMA_signal_15802, MixColumnsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_13770, new_AGEMA_signal_13769, new_AGEMA_signal_13768, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_15060, new_AGEMA_signal_15059, new_AGEMA_signal_15058, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, new_AGEMA_signal_15061, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, new_AGEMA_signal_15805, MixColumnsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, new_AGEMA_signal_13765, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, new_AGEMA_signal_15061, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_13794, new_AGEMA_signal_13793, new_AGEMA_signal_13792, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_15066, new_AGEMA_signal_15065, new_AGEMA_signal_15064, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_15810, new_AGEMA_signal_15809, new_AGEMA_signal_15808, MixColumnsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .b ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, new_AGEMA_signal_13771, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .b ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_15066, new_AGEMA_signal_15065, new_AGEMA_signal_15064, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_14388, new_AGEMA_signal_14387, new_AGEMA_signal_14386, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, new_AGEMA_signal_15067, MixColumnsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .b ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_14388, new_AGEMA_signal_14387, new_AGEMA_signal_14386, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_15072, new_AGEMA_signal_15071, new_AGEMA_signal_15070, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, new_AGEMA_signal_15811, MixColumnsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_13776, new_AGEMA_signal_13775, new_AGEMA_signal_13774, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_15072, new_AGEMA_signal_15071, new_AGEMA_signal_15070, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, new_AGEMA_signal_13783, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_14397, new_AGEMA_signal_14396, new_AGEMA_signal_14395, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, new_AGEMA_signal_15073, MixColumnsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .b ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_14397, new_AGEMA_signal_14396, new_AGEMA_signal_14395, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_14400, new_AGEMA_signal_14399, new_AGEMA_signal_14398, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_15078, new_AGEMA_signal_15077, new_AGEMA_signal_15076, MixColumnsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_14400, new_AGEMA_signal_14399, new_AGEMA_signal_14398, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_14403, new_AGEMA_signal_14402, new_AGEMA_signal_14401, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, new_AGEMA_signal_15079, MixColumnsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_14403, new_AGEMA_signal_14402, new_AGEMA_signal_14401, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_14406, new_AGEMA_signal_14405, new_AGEMA_signal_14404, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_15084, new_AGEMA_signal_15083, new_AGEMA_signal_15082, MixColumnsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_14406, new_AGEMA_signal_14405, new_AGEMA_signal_14404, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, new_AGEMA_signal_15085, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_15816, new_AGEMA_signal_15815, new_AGEMA_signal_15814, MixColumnsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, new_AGEMA_signal_13777, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, new_AGEMA_signal_15085, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_13788, new_AGEMA_signal_13787, new_AGEMA_signal_13786, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_15090, new_AGEMA_signal_15089, new_AGEMA_signal_15088, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, new_AGEMA_signal_15817, MixColumnsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .b ({new_AGEMA_signal_13782, new_AGEMA_signal_13781, new_AGEMA_signal_13780, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .c ({new_AGEMA_signal_15090, new_AGEMA_signal_15089, new_AGEMA_signal_15088, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, new_AGEMA_signal_13789, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .c ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, new_AGEMA_signal_14419, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, new_AGEMA_signal_15091, MixColumnsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .c ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, new_AGEMA_signal_14419, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .c ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_14424, new_AGEMA_signal_14423, new_AGEMA_signal_14422, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .c ({new_AGEMA_signal_15096, new_AGEMA_signal_15095, new_AGEMA_signal_15094, MixColumnsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_14424, new_AGEMA_signal_14423, new_AGEMA_signal_14422, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .c ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .c ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, new_AGEMA_signal_13759, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .c ({new_AGEMA_signal_13764, new_AGEMA_signal_13763, new_AGEMA_signal_13762, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .c ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, new_AGEMA_signal_13765, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .c ({new_AGEMA_signal_13770, new_AGEMA_signal_13769, new_AGEMA_signal_13768, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .c ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, new_AGEMA_signal_13771, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .c ({new_AGEMA_signal_13776, new_AGEMA_signal_13775, new_AGEMA_signal_13774, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .c ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, new_AGEMA_signal_13777, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .c ({new_AGEMA_signal_13782, new_AGEMA_signal_13781, new_AGEMA_signal_13780, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .c ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, new_AGEMA_signal_13783, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .c ({new_AGEMA_signal_13788, new_AGEMA_signal_13787, new_AGEMA_signal_13786, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .c ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, new_AGEMA_signal_13789, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_13794, new_AGEMA_signal_13793, new_AGEMA_signal_13792, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_15099, new_AGEMA_signal_15098, new_AGEMA_signal_15097, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_15822, new_AGEMA_signal_15821, new_AGEMA_signal_15820, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_15099, new_AGEMA_signal_15098, new_AGEMA_signal_15097, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, new_AGEMA_signal_14425, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_15102, new_AGEMA_signal_15101, new_AGEMA_signal_15100, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .c ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, new_AGEMA_signal_14425, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_14430, new_AGEMA_signal_14429, new_AGEMA_signal_14428, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, new_AGEMA_signal_15103, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_14430, new_AGEMA_signal_14429, new_AGEMA_signal_14428, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, new_AGEMA_signal_14431, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_15108, new_AGEMA_signal_15107, new_AGEMA_signal_15106, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, new_AGEMA_signal_14431, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_14436, new_AGEMA_signal_14435, new_AGEMA_signal_14434, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, new_AGEMA_signal_15109, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_14436, new_AGEMA_signal_14435, new_AGEMA_signal_14434, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_15114, new_AGEMA_signal_15113, new_AGEMA_signal_15112, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, new_AGEMA_signal_15823, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_15114, new_AGEMA_signal_15113, new_AGEMA_signal_15112, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, new_AGEMA_signal_15115, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_15828, new_AGEMA_signal_15827, new_AGEMA_signal_15826, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .c ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, new_AGEMA_signal_15115, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, new_AGEMA_signal_14437, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_15120, new_AGEMA_signal_15119, new_AGEMA_signal_15118, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, new_AGEMA_signal_14437, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_14442, new_AGEMA_signal_14441, new_AGEMA_signal_14440, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, new_AGEMA_signal_15121, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_14442, new_AGEMA_signal_14441, new_AGEMA_signal_14440, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, new_AGEMA_signal_14443, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_15126, new_AGEMA_signal_15125, new_AGEMA_signal_15124, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .c ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, new_AGEMA_signal_14443, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_14448, new_AGEMA_signal_14447, new_AGEMA_signal_14446, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, new_AGEMA_signal_15127, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_14448, new_AGEMA_signal_14447, new_AGEMA_signal_14446, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_15132, new_AGEMA_signal_15131, new_AGEMA_signal_15130, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, new_AGEMA_signal_15829, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, new_AGEMA_signal_13855, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_15132, new_AGEMA_signal_15131, new_AGEMA_signal_15130, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, new_AGEMA_signal_15133, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_15834, new_AGEMA_signal_15833, new_AGEMA_signal_15832, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .b ({new_AGEMA_signal_13860, new_AGEMA_signal_13859, new_AGEMA_signal_13858, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .b ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, new_AGEMA_signal_15133, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, new_AGEMA_signal_14455, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_15138, new_AGEMA_signal_15137, new_AGEMA_signal_15136, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .b ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, new_AGEMA_signal_14455, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, new_AGEMA_signal_15139, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, new_AGEMA_signal_15835, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, new_AGEMA_signal_15139, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_14460, new_AGEMA_signal_14459, new_AGEMA_signal_14458, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_15144, new_AGEMA_signal_15143, new_AGEMA_signal_15142, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_14460, new_AGEMA_signal_14459, new_AGEMA_signal_14458, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, new_AGEMA_signal_14461, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, new_AGEMA_signal_15145, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, new_AGEMA_signal_14461, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_14466, new_AGEMA_signal_14465, new_AGEMA_signal_14464, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_15150, new_AGEMA_signal_15149, new_AGEMA_signal_15148, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_14466, new_AGEMA_signal_14465, new_AGEMA_signal_14464, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, new_AGEMA_signal_14467, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, new_AGEMA_signal_15151, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, new_AGEMA_signal_14467, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_15156, new_AGEMA_signal_15155, new_AGEMA_signal_15154, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_15840, new_AGEMA_signal_15839, new_AGEMA_signal_15838, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_13866, new_AGEMA_signal_13865, new_AGEMA_signal_13864, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_15156, new_AGEMA_signal_15155, new_AGEMA_signal_15154, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_15159, new_AGEMA_signal_15158, new_AGEMA_signal_15157, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, new_AGEMA_signal_15841, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, new_AGEMA_signal_13861, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_15159, new_AGEMA_signal_15158, new_AGEMA_signal_15157, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_13890, new_AGEMA_signal_13889, new_AGEMA_signal_13888, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_15162, new_AGEMA_signal_15161, new_AGEMA_signal_15160, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_15846, new_AGEMA_signal_15845, new_AGEMA_signal_15844, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .b ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, new_AGEMA_signal_13867, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .b ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_15162, new_AGEMA_signal_15161, new_AGEMA_signal_15160, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_14484, new_AGEMA_signal_14483, new_AGEMA_signal_14482, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, new_AGEMA_signal_15163, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .b ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_14484, new_AGEMA_signal_14483, new_AGEMA_signal_14482, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_15168, new_AGEMA_signal_15167, new_AGEMA_signal_15166, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, new_AGEMA_signal_15847, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_13872, new_AGEMA_signal_13871, new_AGEMA_signal_13870, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_15168, new_AGEMA_signal_15167, new_AGEMA_signal_15166, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, new_AGEMA_signal_13879, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, new_AGEMA_signal_14491, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, new_AGEMA_signal_15169, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .b ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, new_AGEMA_signal_14491, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_14496, new_AGEMA_signal_14495, new_AGEMA_signal_14494, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_15174, new_AGEMA_signal_15173, new_AGEMA_signal_15172, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_14496, new_AGEMA_signal_14495, new_AGEMA_signal_14494, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, new_AGEMA_signal_14497, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_15177, new_AGEMA_signal_15176, new_AGEMA_signal_15175, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, new_AGEMA_signal_14497, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_14502, new_AGEMA_signal_14501, new_AGEMA_signal_14500, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_15180, new_AGEMA_signal_15179, new_AGEMA_signal_15178, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_14502, new_AGEMA_signal_14501, new_AGEMA_signal_14500, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_15183, new_AGEMA_signal_15182, new_AGEMA_signal_15181, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_15852, new_AGEMA_signal_15851, new_AGEMA_signal_15850, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, new_AGEMA_signal_13873, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_15183, new_AGEMA_signal_15182, new_AGEMA_signal_15181, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_13884, new_AGEMA_signal_13883, new_AGEMA_signal_13882, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_15186, new_AGEMA_signal_15185, new_AGEMA_signal_15184, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_15855, new_AGEMA_signal_15854, new_AGEMA_signal_15853, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .b ({new_AGEMA_signal_13878, new_AGEMA_signal_13877, new_AGEMA_signal_13876, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .c ({new_AGEMA_signal_15186, new_AGEMA_signal_15185, new_AGEMA_signal_15184, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, new_AGEMA_signal_13885, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .c ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, new_AGEMA_signal_14515, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, new_AGEMA_signal_15187, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .c ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, new_AGEMA_signal_14515, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .c ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_14520, new_AGEMA_signal_14519, new_AGEMA_signal_14518, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .c ({new_AGEMA_signal_15192, new_AGEMA_signal_15191, new_AGEMA_signal_15190, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_14520, new_AGEMA_signal_14519, new_AGEMA_signal_14518, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .c ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .c ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, new_AGEMA_signal_13855, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .c ({new_AGEMA_signal_13860, new_AGEMA_signal_13859, new_AGEMA_signal_13858, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .c ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, new_AGEMA_signal_13861, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .c ({new_AGEMA_signal_13866, new_AGEMA_signal_13865, new_AGEMA_signal_13864, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .c ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, new_AGEMA_signal_13867, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .c ({new_AGEMA_signal_13872, new_AGEMA_signal_13871, new_AGEMA_signal_13870, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .c ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, new_AGEMA_signal_13873, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .c ({new_AGEMA_signal_13878, new_AGEMA_signal_13877, new_AGEMA_signal_13876, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .c ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, new_AGEMA_signal_13879, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .c ({new_AGEMA_signal_13884, new_AGEMA_signal_13883, new_AGEMA_signal_13882, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .c ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, new_AGEMA_signal_13885, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_13890, new_AGEMA_signal_13889, new_AGEMA_signal_13888, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14808, new_AGEMA_signal_14807, new_AGEMA_signal_14806, KeyExpansionOutput[0]}), .a ({new_AGEMA_signal_31676, new_AGEMA_signal_31672, new_AGEMA_signal_31668, new_AGEMA_signal_31664}), .c ({new_AGEMA_signal_15198, new_AGEMA_signal_15197, new_AGEMA_signal_15196, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15444, new_AGEMA_signal_15443, new_AGEMA_signal_15442, KeyExpansionOutput[1]}), .a ({new_AGEMA_signal_31692, new_AGEMA_signal_31688, new_AGEMA_signal_31684, new_AGEMA_signal_31680}), .c ({new_AGEMA_signal_15861, new_AGEMA_signal_15860, new_AGEMA_signal_15859, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15411, new_AGEMA_signal_15410, new_AGEMA_signal_15409, KeyExpansionOutput[2]}), .a ({new_AGEMA_signal_31708, new_AGEMA_signal_31704, new_AGEMA_signal_31700, new_AGEMA_signal_31696}), .c ({new_AGEMA_signal_15867, new_AGEMA_signal_15866, new_AGEMA_signal_15865, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15402, new_AGEMA_signal_15401, new_AGEMA_signal_15400, KeyExpansionOutput[3]}), .a ({new_AGEMA_signal_31724, new_AGEMA_signal_31720, new_AGEMA_signal_31716, new_AGEMA_signal_31712}), .c ({new_AGEMA_signal_15873, new_AGEMA_signal_15872, new_AGEMA_signal_15871, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15399, new_AGEMA_signal_15398, new_AGEMA_signal_15397, KeyExpansionOutput[4]}), .a ({new_AGEMA_signal_31740, new_AGEMA_signal_31736, new_AGEMA_signal_31732, new_AGEMA_signal_31728}), .c ({new_AGEMA_signal_15879, new_AGEMA_signal_15878, new_AGEMA_signal_15877, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15396, new_AGEMA_signal_15395, new_AGEMA_signal_15394, KeyExpansionOutput[5]}), .a ({new_AGEMA_signal_31756, new_AGEMA_signal_31752, new_AGEMA_signal_31748, new_AGEMA_signal_31744}), .c ({new_AGEMA_signal_15885, new_AGEMA_signal_15884, new_AGEMA_signal_15883, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15393, new_AGEMA_signal_15392, new_AGEMA_signal_15391, KeyExpansionOutput[6]}), .a ({new_AGEMA_signal_31772, new_AGEMA_signal_31768, new_AGEMA_signal_31764, new_AGEMA_signal_31760}), .c ({new_AGEMA_signal_15891, new_AGEMA_signal_15890, new_AGEMA_signal_15889, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15390, new_AGEMA_signal_15389, new_AGEMA_signal_15388, KeyExpansionOutput[7]}), .a ({new_AGEMA_signal_31788, new_AGEMA_signal_31784, new_AGEMA_signal_31780, new_AGEMA_signal_31776}), .c ({new_AGEMA_signal_15897, new_AGEMA_signal_15896, new_AGEMA_signal_15895, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, new_AGEMA_signal_14713, KeyExpansionOutput[8]}), .a ({new_AGEMA_signal_31804, new_AGEMA_signal_31800, new_AGEMA_signal_31796, new_AGEMA_signal_31792}), .c ({new_AGEMA_signal_15204, new_AGEMA_signal_15203, new_AGEMA_signal_15202, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15387, new_AGEMA_signal_15386, new_AGEMA_signal_15385, KeyExpansionOutput[9]}), .a ({new_AGEMA_signal_31820, new_AGEMA_signal_31816, new_AGEMA_signal_31812, new_AGEMA_signal_31808}), .c ({new_AGEMA_signal_15903, new_AGEMA_signal_15902, new_AGEMA_signal_15901, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15471, new_AGEMA_signal_15470, new_AGEMA_signal_15469, KeyExpansionOutput[10]}), .a ({new_AGEMA_signal_31836, new_AGEMA_signal_31832, new_AGEMA_signal_31828, new_AGEMA_signal_31824}), .c ({new_AGEMA_signal_15909, new_AGEMA_signal_15908, new_AGEMA_signal_15907, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15468, new_AGEMA_signal_15467, new_AGEMA_signal_15466, KeyExpansionOutput[11]}), .a ({new_AGEMA_signal_31852, new_AGEMA_signal_31848, new_AGEMA_signal_31844, new_AGEMA_signal_31840}), .c ({new_AGEMA_signal_15915, new_AGEMA_signal_15914, new_AGEMA_signal_15913, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15465, new_AGEMA_signal_15464, new_AGEMA_signal_15463, KeyExpansionOutput[12]}), .a ({new_AGEMA_signal_31868, new_AGEMA_signal_31864, new_AGEMA_signal_31860, new_AGEMA_signal_31856}), .c ({new_AGEMA_signal_15921, new_AGEMA_signal_15920, new_AGEMA_signal_15919, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15462, new_AGEMA_signal_15461, new_AGEMA_signal_15460, KeyExpansionOutput[13]}), .a ({new_AGEMA_signal_31884, new_AGEMA_signal_31880, new_AGEMA_signal_31876, new_AGEMA_signal_31872}), .c ({new_AGEMA_signal_15927, new_AGEMA_signal_15926, new_AGEMA_signal_15925, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15459, new_AGEMA_signal_15458, new_AGEMA_signal_15457, KeyExpansionOutput[14]}), .a ({new_AGEMA_signal_31900, new_AGEMA_signal_31896, new_AGEMA_signal_31892, new_AGEMA_signal_31888}), .c ({new_AGEMA_signal_15933, new_AGEMA_signal_15932, new_AGEMA_signal_15931, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15456, new_AGEMA_signal_15455, new_AGEMA_signal_15454, KeyExpansionOutput[15]}), .a ({new_AGEMA_signal_31916, new_AGEMA_signal_31912, new_AGEMA_signal_31908, new_AGEMA_signal_31904}), .c ({new_AGEMA_signal_15939, new_AGEMA_signal_15938, new_AGEMA_signal_15937, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, new_AGEMA_signal_14785, KeyExpansionOutput[16]}), .a ({new_AGEMA_signal_31932, new_AGEMA_signal_31928, new_AGEMA_signal_31924, new_AGEMA_signal_31920}), .c ({new_AGEMA_signal_15210, new_AGEMA_signal_15209, new_AGEMA_signal_15208, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15453, new_AGEMA_signal_15452, new_AGEMA_signal_15451, KeyExpansionOutput[17]}), .a ({new_AGEMA_signal_31948, new_AGEMA_signal_31944, new_AGEMA_signal_31940, new_AGEMA_signal_31936}), .c ({new_AGEMA_signal_15945, new_AGEMA_signal_15944, new_AGEMA_signal_15943, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15450, new_AGEMA_signal_15449, new_AGEMA_signal_15448, KeyExpansionOutput[18]}), .a ({new_AGEMA_signal_31964, new_AGEMA_signal_31960, new_AGEMA_signal_31956, new_AGEMA_signal_31952}), .c ({new_AGEMA_signal_15951, new_AGEMA_signal_15950, new_AGEMA_signal_15949, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15447, new_AGEMA_signal_15446, new_AGEMA_signal_15445, KeyExpansionOutput[19]}), .a ({new_AGEMA_signal_31980, new_AGEMA_signal_31976, new_AGEMA_signal_31972, new_AGEMA_signal_31968}), .c ({new_AGEMA_signal_15957, new_AGEMA_signal_15956, new_AGEMA_signal_15955, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15441, new_AGEMA_signal_15440, new_AGEMA_signal_15439, KeyExpansionOutput[20]}), .a ({new_AGEMA_signal_31996, new_AGEMA_signal_31992, new_AGEMA_signal_31988, new_AGEMA_signal_31984}), .c ({new_AGEMA_signal_15963, new_AGEMA_signal_15962, new_AGEMA_signal_15961, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15438, new_AGEMA_signal_15437, new_AGEMA_signal_15436, KeyExpansionOutput[21]}), .a ({new_AGEMA_signal_32012, new_AGEMA_signal_32008, new_AGEMA_signal_32004, new_AGEMA_signal_32000}), .c ({new_AGEMA_signal_15969, new_AGEMA_signal_15968, new_AGEMA_signal_15967, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15435, new_AGEMA_signal_15434, new_AGEMA_signal_15433, KeyExpansionOutput[22]}), .a ({new_AGEMA_signal_32028, new_AGEMA_signal_32024, new_AGEMA_signal_32020, new_AGEMA_signal_32016}), .c ({new_AGEMA_signal_15975, new_AGEMA_signal_15974, new_AGEMA_signal_15973, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15432, new_AGEMA_signal_15431, new_AGEMA_signal_15430, KeyExpansionOutput[23]}), .a ({new_AGEMA_signal_32044, new_AGEMA_signal_32040, new_AGEMA_signal_32036, new_AGEMA_signal_32032}), .c ({new_AGEMA_signal_15981, new_AGEMA_signal_15980, new_AGEMA_signal_15979, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15429, new_AGEMA_signal_15428, new_AGEMA_signal_15427, KeyExpansionOutput[24]}), .a ({new_AGEMA_signal_32060, new_AGEMA_signal_32056, new_AGEMA_signal_32052, new_AGEMA_signal_32048}), .c ({new_AGEMA_signal_15987, new_AGEMA_signal_15986, new_AGEMA_signal_15985, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16050, new_AGEMA_signal_16049, new_AGEMA_signal_16048, KeyExpansionOutput[25]}), .a ({new_AGEMA_signal_32076, new_AGEMA_signal_32072, new_AGEMA_signal_32068, new_AGEMA_signal_32064}), .c ({new_AGEMA_signal_16680, new_AGEMA_signal_16679, new_AGEMA_signal_16678, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, new_AGEMA_signal_16045, KeyExpansionOutput[26]}), .a ({new_AGEMA_signal_32092, new_AGEMA_signal_32088, new_AGEMA_signal_32084, new_AGEMA_signal_32080}), .c ({new_AGEMA_signal_16686, new_AGEMA_signal_16685, new_AGEMA_signal_16684, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16044, new_AGEMA_signal_16043, new_AGEMA_signal_16042, KeyExpansionOutput[27]}), .a ({new_AGEMA_signal_32108, new_AGEMA_signal_32104, new_AGEMA_signal_32100, new_AGEMA_signal_32096}), .c ({new_AGEMA_signal_16692, new_AGEMA_signal_16691, new_AGEMA_signal_16690, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, new_AGEMA_signal_16039, KeyExpansionOutput[28]}), .a ({new_AGEMA_signal_32124, new_AGEMA_signal_32120, new_AGEMA_signal_32116, new_AGEMA_signal_32112}), .c ({new_AGEMA_signal_16698, new_AGEMA_signal_16697, new_AGEMA_signal_16696, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16038, new_AGEMA_signal_16037, new_AGEMA_signal_16036, KeyExpansionOutput[29]}), .a ({new_AGEMA_signal_32140, new_AGEMA_signal_32136, new_AGEMA_signal_32132, new_AGEMA_signal_32128}), .c ({new_AGEMA_signal_16704, new_AGEMA_signal_16703, new_AGEMA_signal_16702, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16035, new_AGEMA_signal_16034, new_AGEMA_signal_16033, KeyExpansionOutput[30]}), .a ({new_AGEMA_signal_32156, new_AGEMA_signal_32152, new_AGEMA_signal_32148, new_AGEMA_signal_32144}), .c ({new_AGEMA_signal_16710, new_AGEMA_signal_16709, new_AGEMA_signal_16708, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_16032, new_AGEMA_signal_16031, new_AGEMA_signal_16030, KeyExpansionOutput[31]}), .a ({new_AGEMA_signal_32172, new_AGEMA_signal_32168, new_AGEMA_signal_32164, new_AGEMA_signal_32160}), .c ({new_AGEMA_signal_16716, new_AGEMA_signal_16715, new_AGEMA_signal_16714, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}), .a ({new_AGEMA_signal_32188, new_AGEMA_signal_32184, new_AGEMA_signal_32180, new_AGEMA_signal_32176}), .c ({new_AGEMA_signal_14526, new_AGEMA_signal_14525, new_AGEMA_signal_14524, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}), .a ({new_AGEMA_signal_32204, new_AGEMA_signal_32200, new_AGEMA_signal_32196, new_AGEMA_signal_32192}), .c ({new_AGEMA_signal_15216, new_AGEMA_signal_15215, new_AGEMA_signal_15214, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}), .a ({new_AGEMA_signal_32220, new_AGEMA_signal_32216, new_AGEMA_signal_32212, new_AGEMA_signal_32208}), .c ({new_AGEMA_signal_15222, new_AGEMA_signal_15221, new_AGEMA_signal_15220, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}), .a ({new_AGEMA_signal_32236, new_AGEMA_signal_32232, new_AGEMA_signal_32228, new_AGEMA_signal_32224}), .c ({new_AGEMA_signal_15228, new_AGEMA_signal_15227, new_AGEMA_signal_15226, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}), .a ({new_AGEMA_signal_32252, new_AGEMA_signal_32248, new_AGEMA_signal_32244, new_AGEMA_signal_32240}), .c ({new_AGEMA_signal_15234, new_AGEMA_signal_15233, new_AGEMA_signal_15232, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}), .a ({new_AGEMA_signal_32268, new_AGEMA_signal_32264, new_AGEMA_signal_32260, new_AGEMA_signal_32256}), .c ({new_AGEMA_signal_15240, new_AGEMA_signal_15239, new_AGEMA_signal_15238, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}), .a ({new_AGEMA_signal_32284, new_AGEMA_signal_32280, new_AGEMA_signal_32276, new_AGEMA_signal_32272}), .c ({new_AGEMA_signal_15246, new_AGEMA_signal_15245, new_AGEMA_signal_15244, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}), .a ({new_AGEMA_signal_32300, new_AGEMA_signal_32296, new_AGEMA_signal_32292, new_AGEMA_signal_32288}), .c ({new_AGEMA_signal_15252, new_AGEMA_signal_15251, new_AGEMA_signal_15250, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}), .a ({new_AGEMA_signal_32316, new_AGEMA_signal_32312, new_AGEMA_signal_32308, new_AGEMA_signal_32304}), .c ({new_AGEMA_signal_14532, new_AGEMA_signal_14531, new_AGEMA_signal_14530, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}), .a ({new_AGEMA_signal_32332, new_AGEMA_signal_32328, new_AGEMA_signal_32324, new_AGEMA_signal_32320}), .c ({new_AGEMA_signal_15258, new_AGEMA_signal_15257, new_AGEMA_signal_15256, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}), .a ({new_AGEMA_signal_32348, new_AGEMA_signal_32344, new_AGEMA_signal_32340, new_AGEMA_signal_32336}), .c ({new_AGEMA_signal_15264, new_AGEMA_signal_15263, new_AGEMA_signal_15262, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}), .a ({new_AGEMA_signal_32364, new_AGEMA_signal_32360, new_AGEMA_signal_32356, new_AGEMA_signal_32352}), .c ({new_AGEMA_signal_15270, new_AGEMA_signal_15269, new_AGEMA_signal_15268, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}), .a ({new_AGEMA_signal_32380, new_AGEMA_signal_32376, new_AGEMA_signal_32372, new_AGEMA_signal_32368}), .c ({new_AGEMA_signal_15276, new_AGEMA_signal_15275, new_AGEMA_signal_15274, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}), .a ({new_AGEMA_signal_32396, new_AGEMA_signal_32392, new_AGEMA_signal_32388, new_AGEMA_signal_32384}), .c ({new_AGEMA_signal_15282, new_AGEMA_signal_15281, new_AGEMA_signal_15280, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}), .a ({new_AGEMA_signal_32412, new_AGEMA_signal_32408, new_AGEMA_signal_32404, new_AGEMA_signal_32400}), .c ({new_AGEMA_signal_15288, new_AGEMA_signal_15287, new_AGEMA_signal_15286, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}), .a ({new_AGEMA_signal_32428, new_AGEMA_signal_32424, new_AGEMA_signal_32420, new_AGEMA_signal_32416}), .c ({new_AGEMA_signal_15294, new_AGEMA_signal_15293, new_AGEMA_signal_15292, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}), .a ({new_AGEMA_signal_32444, new_AGEMA_signal_32440, new_AGEMA_signal_32436, new_AGEMA_signal_32432}), .c ({new_AGEMA_signal_14538, new_AGEMA_signal_14537, new_AGEMA_signal_14536, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}), .a ({new_AGEMA_signal_32460, new_AGEMA_signal_32456, new_AGEMA_signal_32452, new_AGEMA_signal_32448}), .c ({new_AGEMA_signal_15300, new_AGEMA_signal_15299, new_AGEMA_signal_15298, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}), .a ({new_AGEMA_signal_32476, new_AGEMA_signal_32472, new_AGEMA_signal_32468, new_AGEMA_signal_32464}), .c ({new_AGEMA_signal_15306, new_AGEMA_signal_15305, new_AGEMA_signal_15304, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}), .a ({new_AGEMA_signal_32492, new_AGEMA_signal_32488, new_AGEMA_signal_32484, new_AGEMA_signal_32480}), .c ({new_AGEMA_signal_15312, new_AGEMA_signal_15311, new_AGEMA_signal_15310, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}), .a ({new_AGEMA_signal_32508, new_AGEMA_signal_32504, new_AGEMA_signal_32500, new_AGEMA_signal_32496}), .c ({new_AGEMA_signal_15318, new_AGEMA_signal_15317, new_AGEMA_signal_15316, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}), .a ({new_AGEMA_signal_32524, new_AGEMA_signal_32520, new_AGEMA_signal_32516, new_AGEMA_signal_32512}), .c ({new_AGEMA_signal_15324, new_AGEMA_signal_15323, new_AGEMA_signal_15322, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}), .a ({new_AGEMA_signal_32540, new_AGEMA_signal_32536, new_AGEMA_signal_32532, new_AGEMA_signal_32528}), .c ({new_AGEMA_signal_15330, new_AGEMA_signal_15329, new_AGEMA_signal_15328, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}), .a ({new_AGEMA_signal_32556, new_AGEMA_signal_32552, new_AGEMA_signal_32548, new_AGEMA_signal_32544}), .c ({new_AGEMA_signal_15336, new_AGEMA_signal_15335, new_AGEMA_signal_15334, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}), .a ({new_AGEMA_signal_32572, new_AGEMA_signal_32568, new_AGEMA_signal_32564, new_AGEMA_signal_32560}), .c ({new_AGEMA_signal_15342, new_AGEMA_signal_15341, new_AGEMA_signal_15340, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}), .a ({new_AGEMA_signal_32588, new_AGEMA_signal_32584, new_AGEMA_signal_32580, new_AGEMA_signal_32576}), .c ({new_AGEMA_signal_15993, new_AGEMA_signal_15992, new_AGEMA_signal_15991, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}), .a ({new_AGEMA_signal_32604, new_AGEMA_signal_32600, new_AGEMA_signal_32596, new_AGEMA_signal_32592}), .c ({new_AGEMA_signal_15999, new_AGEMA_signal_15998, new_AGEMA_signal_15997, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}), .a ({new_AGEMA_signal_32620, new_AGEMA_signal_32616, new_AGEMA_signal_32612, new_AGEMA_signal_32608}), .c ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, new_AGEMA_signal_16003, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}), .a ({new_AGEMA_signal_32636, new_AGEMA_signal_32632, new_AGEMA_signal_32628, new_AGEMA_signal_32624}), .c ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, new_AGEMA_signal_16009, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}), .a ({new_AGEMA_signal_32652, new_AGEMA_signal_32648, new_AGEMA_signal_32644, new_AGEMA_signal_32640}), .c ({new_AGEMA_signal_16017, new_AGEMA_signal_16016, new_AGEMA_signal_16015, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}), .a ({new_AGEMA_signal_32668, new_AGEMA_signal_32664, new_AGEMA_signal_32660, new_AGEMA_signal_32656}), .c ({new_AGEMA_signal_16023, new_AGEMA_signal_16022, new_AGEMA_signal_16021, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}), .a ({new_AGEMA_signal_32684, new_AGEMA_signal_32680, new_AGEMA_signal_32676, new_AGEMA_signal_32672}), .c ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, new_AGEMA_signal_16027, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}), .a ({new_AGEMA_signal_32700, new_AGEMA_signal_32696, new_AGEMA_signal_32692, new_AGEMA_signal_32688}), .c ({new_AGEMA_signal_13896, new_AGEMA_signal_13895, new_AGEMA_signal_13894, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}), .a ({new_AGEMA_signal_32716, new_AGEMA_signal_32712, new_AGEMA_signal_32708, new_AGEMA_signal_32704}), .c ({new_AGEMA_signal_14544, new_AGEMA_signal_14543, new_AGEMA_signal_14542, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}), .a ({new_AGEMA_signal_32732, new_AGEMA_signal_32728, new_AGEMA_signal_32724, new_AGEMA_signal_32720}), .c ({new_AGEMA_signal_14550, new_AGEMA_signal_14549, new_AGEMA_signal_14548, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}), .a ({new_AGEMA_signal_32748, new_AGEMA_signal_32744, new_AGEMA_signal_32740, new_AGEMA_signal_32736}), .c ({new_AGEMA_signal_14556, new_AGEMA_signal_14555, new_AGEMA_signal_14554, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}), .a ({new_AGEMA_signal_32764, new_AGEMA_signal_32760, new_AGEMA_signal_32756, new_AGEMA_signal_32752}), .c ({new_AGEMA_signal_14562, new_AGEMA_signal_14561, new_AGEMA_signal_14560, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}), .a ({new_AGEMA_signal_32780, new_AGEMA_signal_32776, new_AGEMA_signal_32772, new_AGEMA_signal_32768}), .c ({new_AGEMA_signal_14568, new_AGEMA_signal_14567, new_AGEMA_signal_14566, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}), .a ({new_AGEMA_signal_32796, new_AGEMA_signal_32792, new_AGEMA_signal_32788, new_AGEMA_signal_32784}), .c ({new_AGEMA_signal_14574, new_AGEMA_signal_14573, new_AGEMA_signal_14572, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}), .a ({new_AGEMA_signal_32812, new_AGEMA_signal_32808, new_AGEMA_signal_32804, new_AGEMA_signal_32800}), .c ({new_AGEMA_signal_14580, new_AGEMA_signal_14579, new_AGEMA_signal_14578, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}), .a ({new_AGEMA_signal_32828, new_AGEMA_signal_32824, new_AGEMA_signal_32820, new_AGEMA_signal_32816}), .c ({new_AGEMA_signal_13902, new_AGEMA_signal_13901, new_AGEMA_signal_13900, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}), .a ({new_AGEMA_signal_32844, new_AGEMA_signal_32840, new_AGEMA_signal_32836, new_AGEMA_signal_32832}), .c ({new_AGEMA_signal_14586, new_AGEMA_signal_14585, new_AGEMA_signal_14584, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}), .a ({new_AGEMA_signal_32860, new_AGEMA_signal_32856, new_AGEMA_signal_32852, new_AGEMA_signal_32848}), .c ({new_AGEMA_signal_14592, new_AGEMA_signal_14591, new_AGEMA_signal_14590, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}), .a ({new_AGEMA_signal_32876, new_AGEMA_signal_32872, new_AGEMA_signal_32868, new_AGEMA_signal_32864}), .c ({new_AGEMA_signal_14598, new_AGEMA_signal_14597, new_AGEMA_signal_14596, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}), .a ({new_AGEMA_signal_32892, new_AGEMA_signal_32888, new_AGEMA_signal_32884, new_AGEMA_signal_32880}), .c ({new_AGEMA_signal_14604, new_AGEMA_signal_14603, new_AGEMA_signal_14602, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}), .a ({new_AGEMA_signal_32908, new_AGEMA_signal_32904, new_AGEMA_signal_32900, new_AGEMA_signal_32896}), .c ({new_AGEMA_signal_14610, new_AGEMA_signal_14609, new_AGEMA_signal_14608, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}), .a ({new_AGEMA_signal_32924, new_AGEMA_signal_32920, new_AGEMA_signal_32916, new_AGEMA_signal_32912}), .c ({new_AGEMA_signal_14616, new_AGEMA_signal_14615, new_AGEMA_signal_14614, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}), .a ({new_AGEMA_signal_32940, new_AGEMA_signal_32936, new_AGEMA_signal_32932, new_AGEMA_signal_32928}), .c ({new_AGEMA_signal_14622, new_AGEMA_signal_14621, new_AGEMA_signal_14620, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}), .a ({new_AGEMA_signal_32956, new_AGEMA_signal_32952, new_AGEMA_signal_32948, new_AGEMA_signal_32944}), .c ({new_AGEMA_signal_13908, new_AGEMA_signal_13907, new_AGEMA_signal_13906, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}), .a ({new_AGEMA_signal_32972, new_AGEMA_signal_32968, new_AGEMA_signal_32964, new_AGEMA_signal_32960}), .c ({new_AGEMA_signal_14628, new_AGEMA_signal_14627, new_AGEMA_signal_14626, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}), .a ({new_AGEMA_signal_32988, new_AGEMA_signal_32984, new_AGEMA_signal_32980, new_AGEMA_signal_32976}), .c ({new_AGEMA_signal_14634, new_AGEMA_signal_14633, new_AGEMA_signal_14632, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}), .a ({new_AGEMA_signal_33004, new_AGEMA_signal_33000, new_AGEMA_signal_32996, new_AGEMA_signal_32992}), .c ({new_AGEMA_signal_14640, new_AGEMA_signal_14639, new_AGEMA_signal_14638, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}), .a ({new_AGEMA_signal_33020, new_AGEMA_signal_33016, new_AGEMA_signal_33012, new_AGEMA_signal_33008}), .c ({new_AGEMA_signal_14646, new_AGEMA_signal_14645, new_AGEMA_signal_14644, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}), .a ({new_AGEMA_signal_33036, new_AGEMA_signal_33032, new_AGEMA_signal_33028, new_AGEMA_signal_33024}), .c ({new_AGEMA_signal_14652, new_AGEMA_signal_14651, new_AGEMA_signal_14650, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}), .a ({new_AGEMA_signal_33052, new_AGEMA_signal_33048, new_AGEMA_signal_33044, new_AGEMA_signal_33040}), .c ({new_AGEMA_signal_14658, new_AGEMA_signal_14657, new_AGEMA_signal_14656, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}), .a ({new_AGEMA_signal_33068, new_AGEMA_signal_33064, new_AGEMA_signal_33060, new_AGEMA_signal_33056}), .c ({new_AGEMA_signal_14664, new_AGEMA_signal_14663, new_AGEMA_signal_14662, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}), .a ({new_AGEMA_signal_33084, new_AGEMA_signal_33080, new_AGEMA_signal_33076, new_AGEMA_signal_33072}), .c ({new_AGEMA_signal_14670, new_AGEMA_signal_14669, new_AGEMA_signal_14668, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}), .a ({new_AGEMA_signal_33100, new_AGEMA_signal_33096, new_AGEMA_signal_33092, new_AGEMA_signal_33088}), .c ({new_AGEMA_signal_15348, new_AGEMA_signal_15347, new_AGEMA_signal_15346, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}), .a ({new_AGEMA_signal_33116, new_AGEMA_signal_33112, new_AGEMA_signal_33108, new_AGEMA_signal_33104}), .c ({new_AGEMA_signal_15354, new_AGEMA_signal_15353, new_AGEMA_signal_15352, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}), .a ({new_AGEMA_signal_33132, new_AGEMA_signal_33128, new_AGEMA_signal_33124, new_AGEMA_signal_33120}), .c ({new_AGEMA_signal_15360, new_AGEMA_signal_15359, new_AGEMA_signal_15358, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}), .a ({new_AGEMA_signal_33148, new_AGEMA_signal_33144, new_AGEMA_signal_33140, new_AGEMA_signal_33136}), .c ({new_AGEMA_signal_15366, new_AGEMA_signal_15365, new_AGEMA_signal_15364, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}), .a ({new_AGEMA_signal_33164, new_AGEMA_signal_33160, new_AGEMA_signal_33156, new_AGEMA_signal_33152}), .c ({new_AGEMA_signal_15372, new_AGEMA_signal_15371, new_AGEMA_signal_15370, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}), .a ({new_AGEMA_signal_33180, new_AGEMA_signal_33176, new_AGEMA_signal_33172, new_AGEMA_signal_33168}), .c ({new_AGEMA_signal_15378, new_AGEMA_signal_15377, new_AGEMA_signal_15376, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}), .a ({new_AGEMA_signal_33196, new_AGEMA_signal_33192, new_AGEMA_signal_33188, new_AGEMA_signal_33184}), .c ({new_AGEMA_signal_15384, new_AGEMA_signal_15383, new_AGEMA_signal_15382, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}), .a ({new_AGEMA_signal_33212, new_AGEMA_signal_33208, new_AGEMA_signal_33204, new_AGEMA_signal_33200}), .c ({new_AGEMA_signal_13398, new_AGEMA_signal_13397, new_AGEMA_signal_13396, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}), .a ({new_AGEMA_signal_33228, new_AGEMA_signal_33224, new_AGEMA_signal_33220, new_AGEMA_signal_33216}), .c ({new_AGEMA_signal_13914, new_AGEMA_signal_13913, new_AGEMA_signal_13912, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}), .a ({new_AGEMA_signal_33244, new_AGEMA_signal_33240, new_AGEMA_signal_33236, new_AGEMA_signal_33232}), .c ({new_AGEMA_signal_13920, new_AGEMA_signal_13919, new_AGEMA_signal_13918, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}), .a ({new_AGEMA_signal_33260, new_AGEMA_signal_33256, new_AGEMA_signal_33252, new_AGEMA_signal_33248}), .c ({new_AGEMA_signal_13926, new_AGEMA_signal_13925, new_AGEMA_signal_13924, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}), .a ({new_AGEMA_signal_33276, new_AGEMA_signal_33272, new_AGEMA_signal_33268, new_AGEMA_signal_33264}), .c ({new_AGEMA_signal_13932, new_AGEMA_signal_13931, new_AGEMA_signal_13930, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}), .a ({new_AGEMA_signal_33292, new_AGEMA_signal_33288, new_AGEMA_signal_33284, new_AGEMA_signal_33280}), .c ({new_AGEMA_signal_13938, new_AGEMA_signal_13937, new_AGEMA_signal_13936, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}), .a ({new_AGEMA_signal_33308, new_AGEMA_signal_33304, new_AGEMA_signal_33300, new_AGEMA_signal_33296}), .c ({new_AGEMA_signal_13944, new_AGEMA_signal_13943, new_AGEMA_signal_13942, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}), .a ({new_AGEMA_signal_33324, new_AGEMA_signal_33320, new_AGEMA_signal_33316, new_AGEMA_signal_33312}), .c ({new_AGEMA_signal_13950, new_AGEMA_signal_13949, new_AGEMA_signal_13948, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}), .a ({new_AGEMA_signal_33340, new_AGEMA_signal_33336, new_AGEMA_signal_33332, new_AGEMA_signal_33328}), .c ({new_AGEMA_signal_13404, new_AGEMA_signal_13403, new_AGEMA_signal_13402, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}), .a ({new_AGEMA_signal_33356, new_AGEMA_signal_33352, new_AGEMA_signal_33348, new_AGEMA_signal_33344}), .c ({new_AGEMA_signal_13956, new_AGEMA_signal_13955, new_AGEMA_signal_13954, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}), .a ({new_AGEMA_signal_33372, new_AGEMA_signal_33368, new_AGEMA_signal_33364, new_AGEMA_signal_33360}), .c ({new_AGEMA_signal_13962, new_AGEMA_signal_13961, new_AGEMA_signal_13960, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}), .a ({new_AGEMA_signal_33388, new_AGEMA_signal_33384, new_AGEMA_signal_33380, new_AGEMA_signal_33376}), .c ({new_AGEMA_signal_13968, new_AGEMA_signal_13967, new_AGEMA_signal_13966, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}), .a ({new_AGEMA_signal_33404, new_AGEMA_signal_33400, new_AGEMA_signal_33396, new_AGEMA_signal_33392}), .c ({new_AGEMA_signal_13974, new_AGEMA_signal_13973, new_AGEMA_signal_13972, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}), .a ({new_AGEMA_signal_33420, new_AGEMA_signal_33416, new_AGEMA_signal_33412, new_AGEMA_signal_33408}), .c ({new_AGEMA_signal_13980, new_AGEMA_signal_13979, new_AGEMA_signal_13978, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}), .a ({new_AGEMA_signal_33436, new_AGEMA_signal_33432, new_AGEMA_signal_33428, new_AGEMA_signal_33424}), .c ({new_AGEMA_signal_13986, new_AGEMA_signal_13985, new_AGEMA_signal_13984, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}), .a ({new_AGEMA_signal_33452, new_AGEMA_signal_33448, new_AGEMA_signal_33444, new_AGEMA_signal_33440}), .c ({new_AGEMA_signal_13992, new_AGEMA_signal_13991, new_AGEMA_signal_13990, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}), .a ({new_AGEMA_signal_33468, new_AGEMA_signal_33464, new_AGEMA_signal_33460, new_AGEMA_signal_33456}), .c ({new_AGEMA_signal_13410, new_AGEMA_signal_13409, new_AGEMA_signal_13408, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}), .a ({new_AGEMA_signal_33484, new_AGEMA_signal_33480, new_AGEMA_signal_33476, new_AGEMA_signal_33472}), .c ({new_AGEMA_signal_13998, new_AGEMA_signal_13997, new_AGEMA_signal_13996, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}), .a ({new_AGEMA_signal_33500, new_AGEMA_signal_33496, new_AGEMA_signal_33492, new_AGEMA_signal_33488}), .c ({new_AGEMA_signal_14004, new_AGEMA_signal_14003, new_AGEMA_signal_14002, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}), .a ({new_AGEMA_signal_33516, new_AGEMA_signal_33512, new_AGEMA_signal_33508, new_AGEMA_signal_33504}), .c ({new_AGEMA_signal_14010, new_AGEMA_signal_14009, new_AGEMA_signal_14008, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}), .a ({new_AGEMA_signal_33532, new_AGEMA_signal_33528, new_AGEMA_signal_33524, new_AGEMA_signal_33520}), .c ({new_AGEMA_signal_14016, new_AGEMA_signal_14015, new_AGEMA_signal_14014, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}), .a ({new_AGEMA_signal_33548, new_AGEMA_signal_33544, new_AGEMA_signal_33540, new_AGEMA_signal_33536}), .c ({new_AGEMA_signal_14022, new_AGEMA_signal_14021, new_AGEMA_signal_14020, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}), .a ({new_AGEMA_signal_33564, new_AGEMA_signal_33560, new_AGEMA_signal_33556, new_AGEMA_signal_33552}), .c ({new_AGEMA_signal_14028, new_AGEMA_signal_14027, new_AGEMA_signal_14026, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}), .a ({new_AGEMA_signal_33580, new_AGEMA_signal_33576, new_AGEMA_signal_33572, new_AGEMA_signal_33568}), .c ({new_AGEMA_signal_14034, new_AGEMA_signal_14033, new_AGEMA_signal_14032, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}), .a ({new_AGEMA_signal_33596, new_AGEMA_signal_33592, new_AGEMA_signal_33588, new_AGEMA_signal_33584}), .c ({new_AGEMA_signal_14040, new_AGEMA_signal_14039, new_AGEMA_signal_14038, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}), .a ({new_AGEMA_signal_33612, new_AGEMA_signal_33608, new_AGEMA_signal_33604, new_AGEMA_signal_33600}), .c ({new_AGEMA_signal_14676, new_AGEMA_signal_14675, new_AGEMA_signal_14674, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}), .a ({new_AGEMA_signal_33628, new_AGEMA_signal_33624, new_AGEMA_signal_33620, new_AGEMA_signal_33616}), .c ({new_AGEMA_signal_14682, new_AGEMA_signal_14681, new_AGEMA_signal_14680, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}), .a ({new_AGEMA_signal_33644, new_AGEMA_signal_33640, new_AGEMA_signal_33636, new_AGEMA_signal_33632}), .c ({new_AGEMA_signal_14688, new_AGEMA_signal_14687, new_AGEMA_signal_14686, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}), .a ({new_AGEMA_signal_33660, new_AGEMA_signal_33656, new_AGEMA_signal_33652, new_AGEMA_signal_33648}), .c ({new_AGEMA_signal_14694, new_AGEMA_signal_14693, new_AGEMA_signal_14692, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}), .a ({new_AGEMA_signal_33676, new_AGEMA_signal_33672, new_AGEMA_signal_33668, new_AGEMA_signal_33664}), .c ({new_AGEMA_signal_14700, new_AGEMA_signal_14699, new_AGEMA_signal_14698, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}), .a ({new_AGEMA_signal_33692, new_AGEMA_signal_33688, new_AGEMA_signal_33684, new_AGEMA_signal_33680}), .c ({new_AGEMA_signal_14706, new_AGEMA_signal_14705, new_AGEMA_signal_14704, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_26156), .b ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}), .a ({new_AGEMA_signal_33708, new_AGEMA_signal_33704, new_AGEMA_signal_33700, new_AGEMA_signal_33696}), .c ({new_AGEMA_signal_14712, new_AGEMA_signal_14711, new_AGEMA_signal_14710, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_33724, new_AGEMA_signal_33720, new_AGEMA_signal_33716, new_AGEMA_signal_33712}), .b ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_15387, new_AGEMA_signal_15386, new_AGEMA_signal_15385, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_33740, new_AGEMA_signal_33736, new_AGEMA_signal_33732, new_AGEMA_signal_33728}), .b ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, new_AGEMA_signal_14713, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_33756, new_AGEMA_signal_33752, new_AGEMA_signal_33748, new_AGEMA_signal_33744}), .b ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_15390, new_AGEMA_signal_15389, new_AGEMA_signal_15388, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_33772, new_AGEMA_signal_33768, new_AGEMA_signal_33764, new_AGEMA_signal_33760}), .b ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_15393, new_AGEMA_signal_15392, new_AGEMA_signal_15391, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_33788, new_AGEMA_signal_33784, new_AGEMA_signal_33780, new_AGEMA_signal_33776}), .b ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_15396, new_AGEMA_signal_15395, new_AGEMA_signal_15394, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_33804, new_AGEMA_signal_33800, new_AGEMA_signal_33796, new_AGEMA_signal_33792}), .b ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_15399, new_AGEMA_signal_15398, new_AGEMA_signal_15397, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_33820, new_AGEMA_signal_33816, new_AGEMA_signal_33812, new_AGEMA_signal_33808}), .b ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_33836, new_AGEMA_signal_33832, new_AGEMA_signal_33828, new_AGEMA_signal_33824}), .b ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_33852, new_AGEMA_signal_33848, new_AGEMA_signal_33844, new_AGEMA_signal_33840}), .b ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_33868, new_AGEMA_signal_33864, new_AGEMA_signal_33860, new_AGEMA_signal_33856}), .b ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_33884, new_AGEMA_signal_33880, new_AGEMA_signal_33876, new_AGEMA_signal_33872}), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_15402, new_AGEMA_signal_15401, new_AGEMA_signal_15400, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_33900, new_AGEMA_signal_33896, new_AGEMA_signal_33892, new_AGEMA_signal_33888}), .b ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_33916, new_AGEMA_signal_33912, new_AGEMA_signal_33908, new_AGEMA_signal_33904}), .b ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_33932, new_AGEMA_signal_33928, new_AGEMA_signal_33924, new_AGEMA_signal_33920}), .b ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_33948, new_AGEMA_signal_33944, new_AGEMA_signal_33940, new_AGEMA_signal_33936}), .b ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_33964, new_AGEMA_signal_33960, new_AGEMA_signal_33956, new_AGEMA_signal_33952}), .b ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_33980, new_AGEMA_signal_33976, new_AGEMA_signal_33972, new_AGEMA_signal_33968}), .b ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_33996, new_AGEMA_signal_33992, new_AGEMA_signal_33988, new_AGEMA_signal_33984}), .b ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_34012, new_AGEMA_signal_34008, new_AGEMA_signal_34004, new_AGEMA_signal_34000}), .b ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_34028, new_AGEMA_signal_34024, new_AGEMA_signal_34020, new_AGEMA_signal_34016}), .b ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_34044, new_AGEMA_signal_34040, new_AGEMA_signal_34036, new_AGEMA_signal_34032}), .b ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_34060, new_AGEMA_signal_34056, new_AGEMA_signal_34052, new_AGEMA_signal_34048}), .b ({new_AGEMA_signal_13050, new_AGEMA_signal_13049, new_AGEMA_signal_13048, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_34076, new_AGEMA_signal_34072, new_AGEMA_signal_34068, new_AGEMA_signal_34064}), .b ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_16032, new_AGEMA_signal_16031, new_AGEMA_signal_16030, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_34092, new_AGEMA_signal_34088, new_AGEMA_signal_34084, new_AGEMA_signal_34080}), .b ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_34108, new_AGEMA_signal_34104, new_AGEMA_signal_34100, new_AGEMA_signal_34096}), .b ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_34124, new_AGEMA_signal_34120, new_AGEMA_signal_34116, new_AGEMA_signal_34112}), .b ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_16035, new_AGEMA_signal_16034, new_AGEMA_signal_16033, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_34140, new_AGEMA_signal_34136, new_AGEMA_signal_34132, new_AGEMA_signal_34128}), .b ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_34156, new_AGEMA_signal_34152, new_AGEMA_signal_34148, new_AGEMA_signal_34144}), .b ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_34172, new_AGEMA_signal_34168, new_AGEMA_signal_34164, new_AGEMA_signal_34160}), .b ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_15411, new_AGEMA_signal_15410, new_AGEMA_signal_15409, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_34188, new_AGEMA_signal_34184, new_AGEMA_signal_34180, new_AGEMA_signal_34176}), .b ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_34204, new_AGEMA_signal_34200, new_AGEMA_signal_34196, new_AGEMA_signal_34192}), .b ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_34220, new_AGEMA_signal_34216, new_AGEMA_signal_34212, new_AGEMA_signal_34208}), .b ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, new_AGEMA_signal_13051, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_34236, new_AGEMA_signal_34232, new_AGEMA_signal_34228, new_AGEMA_signal_34224}), .b ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_16038, new_AGEMA_signal_16037, new_AGEMA_signal_16036, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_34252, new_AGEMA_signal_34248, new_AGEMA_signal_34244, new_AGEMA_signal_34240}), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_34268, new_AGEMA_signal_34264, new_AGEMA_signal_34260, new_AGEMA_signal_34256}), .b ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_34284, new_AGEMA_signal_34280, new_AGEMA_signal_34276, new_AGEMA_signal_34272}), .b ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, new_AGEMA_signal_16039, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_34300, new_AGEMA_signal_34296, new_AGEMA_signal_34292, new_AGEMA_signal_34288}), .b ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_34316, new_AGEMA_signal_34312, new_AGEMA_signal_34308, new_AGEMA_signal_34304}), .b ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_34332, new_AGEMA_signal_34328, new_AGEMA_signal_34324, new_AGEMA_signal_34320}), .b ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_16044, new_AGEMA_signal_16043, new_AGEMA_signal_16042, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_34348, new_AGEMA_signal_34344, new_AGEMA_signal_34340, new_AGEMA_signal_34336}), .b ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_34364, new_AGEMA_signal_34360, new_AGEMA_signal_34356, new_AGEMA_signal_34352}), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_34380, new_AGEMA_signal_34376, new_AGEMA_signal_34372, new_AGEMA_signal_34368}), .b ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, new_AGEMA_signal_16045, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_34396, new_AGEMA_signal_34392, new_AGEMA_signal_34388, new_AGEMA_signal_34384}), .b ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_34412, new_AGEMA_signal_34408, new_AGEMA_signal_34404, new_AGEMA_signal_34400}), .b ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_34428, new_AGEMA_signal_34424, new_AGEMA_signal_34420, new_AGEMA_signal_34416}), .b ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_16050, new_AGEMA_signal_16049, new_AGEMA_signal_16048, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_34444, new_AGEMA_signal_34440, new_AGEMA_signal_34436, new_AGEMA_signal_34432}), .b ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_34460, new_AGEMA_signal_34456, new_AGEMA_signal_34452, new_AGEMA_signal_34448}), .b ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_34476, new_AGEMA_signal_34472, new_AGEMA_signal_34468, new_AGEMA_signal_34464}), .b ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_15429, new_AGEMA_signal_15428, new_AGEMA_signal_15427, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_34492, new_AGEMA_signal_34488, new_AGEMA_signal_34484, new_AGEMA_signal_34480}), .b ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_34508, new_AGEMA_signal_34504, new_AGEMA_signal_34500, new_AGEMA_signal_34496}), .b ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_34524, new_AGEMA_signal_34520, new_AGEMA_signal_34516, new_AGEMA_signal_34512}), .b ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_15432, new_AGEMA_signal_15431, new_AGEMA_signal_15430, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_34540, new_AGEMA_signal_34536, new_AGEMA_signal_34532, new_AGEMA_signal_34528}), .b ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_34556, new_AGEMA_signal_34552, new_AGEMA_signal_34548, new_AGEMA_signal_34544}), .b ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_34572, new_AGEMA_signal_34568, new_AGEMA_signal_34564, new_AGEMA_signal_34560}), .b ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_15435, new_AGEMA_signal_15434, new_AGEMA_signal_15433, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_34588, new_AGEMA_signal_34584, new_AGEMA_signal_34580, new_AGEMA_signal_34576}), .b ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_34604, new_AGEMA_signal_34600, new_AGEMA_signal_34596, new_AGEMA_signal_34592}), .b ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_34620, new_AGEMA_signal_34616, new_AGEMA_signal_34612, new_AGEMA_signal_34608}), .b ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_15438, new_AGEMA_signal_15437, new_AGEMA_signal_15436, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_34636, new_AGEMA_signal_34632, new_AGEMA_signal_34628, new_AGEMA_signal_34624}), .b ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_34652, new_AGEMA_signal_34648, new_AGEMA_signal_34644, new_AGEMA_signal_34640}), .b ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_34668, new_AGEMA_signal_34664, new_AGEMA_signal_34660, new_AGEMA_signal_34656}), .b ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_15441, new_AGEMA_signal_15440, new_AGEMA_signal_15439, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_34684, new_AGEMA_signal_34680, new_AGEMA_signal_34676, new_AGEMA_signal_34672}), .b ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_34700, new_AGEMA_signal_34696, new_AGEMA_signal_34692, new_AGEMA_signal_34688}), .b ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_34716, new_AGEMA_signal_34712, new_AGEMA_signal_34708, new_AGEMA_signal_34704}), .b ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_15444, new_AGEMA_signal_15443, new_AGEMA_signal_15442, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_34732, new_AGEMA_signal_34728, new_AGEMA_signal_34724, new_AGEMA_signal_34720}), .b ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_34748, new_AGEMA_signal_34744, new_AGEMA_signal_34740, new_AGEMA_signal_34736}), .b ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_34764, new_AGEMA_signal_34760, new_AGEMA_signal_34756, new_AGEMA_signal_34752}), .b ({new_AGEMA_signal_13056, new_AGEMA_signal_13055, new_AGEMA_signal_13054, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_34780, new_AGEMA_signal_34776, new_AGEMA_signal_34772, new_AGEMA_signal_34768}), .b ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_15447, new_AGEMA_signal_15446, new_AGEMA_signal_15445, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_34796, new_AGEMA_signal_34792, new_AGEMA_signal_34788, new_AGEMA_signal_34784}), .b ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_34812, new_AGEMA_signal_34808, new_AGEMA_signal_34804, new_AGEMA_signal_34800}), .b ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_34828, new_AGEMA_signal_34824, new_AGEMA_signal_34820, new_AGEMA_signal_34816}), .b ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_15450, new_AGEMA_signal_15449, new_AGEMA_signal_15448, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_34844, new_AGEMA_signal_34840, new_AGEMA_signal_34836, new_AGEMA_signal_34832}), .b ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_34860, new_AGEMA_signal_34856, new_AGEMA_signal_34852, new_AGEMA_signal_34848}), .b ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_34876, new_AGEMA_signal_34872, new_AGEMA_signal_34868, new_AGEMA_signal_34864}), .b ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_15453, new_AGEMA_signal_15452, new_AGEMA_signal_15451, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_34892, new_AGEMA_signal_34888, new_AGEMA_signal_34884, new_AGEMA_signal_34880}), .b ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_34908, new_AGEMA_signal_34904, new_AGEMA_signal_34900, new_AGEMA_signal_34896}), .b ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_34924, new_AGEMA_signal_34920, new_AGEMA_signal_34916, new_AGEMA_signal_34912}), .b ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, new_AGEMA_signal_14785, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_34940, new_AGEMA_signal_34936, new_AGEMA_signal_34932, new_AGEMA_signal_34928}), .b ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_34956, new_AGEMA_signal_34952, new_AGEMA_signal_34948, new_AGEMA_signal_34944}), .b ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_34972, new_AGEMA_signal_34968, new_AGEMA_signal_34964, new_AGEMA_signal_34960}), .b ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_15456, new_AGEMA_signal_15455, new_AGEMA_signal_15454, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_34988, new_AGEMA_signal_34984, new_AGEMA_signal_34980, new_AGEMA_signal_34976}), .b ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_35004, new_AGEMA_signal_35000, new_AGEMA_signal_34996, new_AGEMA_signal_34992}), .b ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_35020, new_AGEMA_signal_35016, new_AGEMA_signal_35012, new_AGEMA_signal_35008}), .b ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_15459, new_AGEMA_signal_15458, new_AGEMA_signal_15457, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_35036, new_AGEMA_signal_35032, new_AGEMA_signal_35028, new_AGEMA_signal_35024}), .b ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_35052, new_AGEMA_signal_35048, new_AGEMA_signal_35044, new_AGEMA_signal_35040}), .b ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_35068, new_AGEMA_signal_35064, new_AGEMA_signal_35060, new_AGEMA_signal_35056}), .b ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_15462, new_AGEMA_signal_15461, new_AGEMA_signal_15460, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_35084, new_AGEMA_signal_35080, new_AGEMA_signal_35076, new_AGEMA_signal_35072}), .b ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_35100, new_AGEMA_signal_35096, new_AGEMA_signal_35092, new_AGEMA_signal_35088}), .b ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_35116, new_AGEMA_signal_35112, new_AGEMA_signal_35108, new_AGEMA_signal_35104}), .b ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_15465, new_AGEMA_signal_15464, new_AGEMA_signal_15463, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_35132, new_AGEMA_signal_35128, new_AGEMA_signal_35124, new_AGEMA_signal_35120}), .b ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_35148, new_AGEMA_signal_35144, new_AGEMA_signal_35140, new_AGEMA_signal_35136}), .b ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_35164, new_AGEMA_signal_35160, new_AGEMA_signal_35156, new_AGEMA_signal_35152}), .b ({new_AGEMA_signal_13488, new_AGEMA_signal_13487, new_AGEMA_signal_13486, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_35180, new_AGEMA_signal_35176, new_AGEMA_signal_35172, new_AGEMA_signal_35168}), .b ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, new_AGEMA_signal_13489, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_35196, new_AGEMA_signal_35192, new_AGEMA_signal_35188, new_AGEMA_signal_35184}), .b ({new_AGEMA_signal_13494, new_AGEMA_signal_13493, new_AGEMA_signal_13492, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_35212, new_AGEMA_signal_35208, new_AGEMA_signal_35204, new_AGEMA_signal_35200}), .b ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, new_AGEMA_signal_13495, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_35228, new_AGEMA_signal_35224, new_AGEMA_signal_35220, new_AGEMA_signal_35216}), .b ({new_AGEMA_signal_13500, new_AGEMA_signal_13499, new_AGEMA_signal_13498, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_35244, new_AGEMA_signal_35240, new_AGEMA_signal_35236, new_AGEMA_signal_35232}), .b ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, new_AGEMA_signal_13501, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_35260, new_AGEMA_signal_35256, new_AGEMA_signal_35252, new_AGEMA_signal_35248}), .b ({new_AGEMA_signal_13506, new_AGEMA_signal_13505, new_AGEMA_signal_13504, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_35276, new_AGEMA_signal_35272, new_AGEMA_signal_35268, new_AGEMA_signal_35264}), .b ({new_AGEMA_signal_12972, new_AGEMA_signal_12971, new_AGEMA_signal_12970, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_35292, new_AGEMA_signal_35288, new_AGEMA_signal_35284, new_AGEMA_signal_35280}), .b ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_15468, new_AGEMA_signal_15467, new_AGEMA_signal_15466, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_35308, new_AGEMA_signal_35304, new_AGEMA_signal_35300, new_AGEMA_signal_35296}), .b ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_35324, new_AGEMA_signal_35320, new_AGEMA_signal_35316, new_AGEMA_signal_35312}), .b ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_35340, new_AGEMA_signal_35336, new_AGEMA_signal_35332, new_AGEMA_signal_35328}), .b ({new_AGEMA_signal_12996, new_AGEMA_signal_12995, new_AGEMA_signal_12994, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_35356, new_AGEMA_signal_35352, new_AGEMA_signal_35348, new_AGEMA_signal_35344}), .b ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, new_AGEMA_signal_12997, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_35372, new_AGEMA_signal_35368, new_AGEMA_signal_35364, new_AGEMA_signal_35360}), .b ({new_AGEMA_signal_13002, new_AGEMA_signal_13001, new_AGEMA_signal_13000, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_35388, new_AGEMA_signal_35384, new_AGEMA_signal_35380, new_AGEMA_signal_35376}), .b ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, new_AGEMA_signal_13003, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_35404, new_AGEMA_signal_35400, new_AGEMA_signal_35396, new_AGEMA_signal_35392}), .b ({new_AGEMA_signal_13008, new_AGEMA_signal_13007, new_AGEMA_signal_13006, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_35420, new_AGEMA_signal_35416, new_AGEMA_signal_35412, new_AGEMA_signal_35408}), .b ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, new_AGEMA_signal_13009, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_35436, new_AGEMA_signal_35432, new_AGEMA_signal_35428, new_AGEMA_signal_35424}), .b ({new_AGEMA_signal_13014, new_AGEMA_signal_13013, new_AGEMA_signal_13012, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_35452, new_AGEMA_signal_35448, new_AGEMA_signal_35444, new_AGEMA_signal_35440}), .b ({new_AGEMA_signal_12366, new_AGEMA_signal_12365, new_AGEMA_signal_12364, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_35468, new_AGEMA_signal_35464, new_AGEMA_signal_35460, new_AGEMA_signal_35456}), .b ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, new_AGEMA_signal_13015, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_35484, new_AGEMA_signal_35480, new_AGEMA_signal_35476, new_AGEMA_signal_35472}), .b ({new_AGEMA_signal_13020, new_AGEMA_signal_13019, new_AGEMA_signal_13018, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_35500, new_AGEMA_signal_35496, new_AGEMA_signal_35492, new_AGEMA_signal_35488}), .b ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_15471, new_AGEMA_signal_15470, new_AGEMA_signal_15469, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_35516, new_AGEMA_signal_35512, new_AGEMA_signal_35508, new_AGEMA_signal_35504}), .b ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_35532, new_AGEMA_signal_35528, new_AGEMA_signal_35524, new_AGEMA_signal_35520}), .b ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_35548, new_AGEMA_signal_35544, new_AGEMA_signal_35540, new_AGEMA_signal_35536}), .b ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, new_AGEMA_signal_13021, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_35564, new_AGEMA_signal_35560, new_AGEMA_signal_35556, new_AGEMA_signal_35552}), .b ({new_AGEMA_signal_13026, new_AGEMA_signal_13025, new_AGEMA_signal_13024, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_35580, new_AGEMA_signal_35576, new_AGEMA_signal_35572, new_AGEMA_signal_35568}), .b ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, new_AGEMA_signal_13027, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_35596, new_AGEMA_signal_35592, new_AGEMA_signal_35588, new_AGEMA_signal_35584}), .b ({new_AGEMA_signal_13032, new_AGEMA_signal_13031, new_AGEMA_signal_13030, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_35612, new_AGEMA_signal_35608, new_AGEMA_signal_35604, new_AGEMA_signal_35600}), .b ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, new_AGEMA_signal_13033, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_35628, new_AGEMA_signal_35624, new_AGEMA_signal_35620, new_AGEMA_signal_35616}), .b ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, new_AGEMA_signal_12397, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_35644, new_AGEMA_signal_35640, new_AGEMA_signal_35636, new_AGEMA_signal_35632}), .b ({new_AGEMA_signal_13038, new_AGEMA_signal_13037, new_AGEMA_signal_13036, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_35660, new_AGEMA_signal_35656, new_AGEMA_signal_35652, new_AGEMA_signal_35648}), .b ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, new_AGEMA_signal_13039, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_35676, new_AGEMA_signal_35672, new_AGEMA_signal_35668, new_AGEMA_signal_35664}), .b ({new_AGEMA_signal_13044, new_AGEMA_signal_13043, new_AGEMA_signal_13042, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_35692, new_AGEMA_signal_35688, new_AGEMA_signal_35684, new_AGEMA_signal_35680}), .b ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, new_AGEMA_signal_13045, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_35708, new_AGEMA_signal_35704, new_AGEMA_signal_35700, new_AGEMA_signal_35696}), .b ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_14808, new_AGEMA_signal_14807, new_AGEMA_signal_14806, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_35724, new_AGEMA_signal_35720, new_AGEMA_signal_35716, new_AGEMA_signal_35712}), .b ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_35740, new_AGEMA_signal_35736, new_AGEMA_signal_35732, new_AGEMA_signal_35728}), .b ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_35756, new_AGEMA_signal_35752, new_AGEMA_signal_35748, new_AGEMA_signal_35744}), .b ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, new_AGEMA_signal_12430, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, new_AGEMA_signal_12973, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35760}), .c ({new_AGEMA_signal_13488, new_AGEMA_signal_13487, new_AGEMA_signal_13486, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_12978, new_AGEMA_signal_12977, new_AGEMA_signal_12976, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35764}), .c ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, new_AGEMA_signal_13489, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, new_AGEMA_signal_12979, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35768}), .c ({new_AGEMA_signal_13494, new_AGEMA_signal_13493, new_AGEMA_signal_13492, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_12984, new_AGEMA_signal_12983, new_AGEMA_signal_12982, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35772}), .c ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, new_AGEMA_signal_13495, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, new_AGEMA_signal_12985, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35776}), .c ({new_AGEMA_signal_13500, new_AGEMA_signal_13499, new_AGEMA_signal_13498, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_12990, new_AGEMA_signal_12989, new_AGEMA_signal_12988, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35780}), .c ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, new_AGEMA_signal_13501, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, new_AGEMA_signal_12991, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35784}), .c ({new_AGEMA_signal_13506, new_AGEMA_signal_13505, new_AGEMA_signal_13504, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, new_AGEMA_signal_12331, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_35788}), .c ({new_AGEMA_signal_12972, new_AGEMA_signal_12971, new_AGEMA_signal_12970, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_35800, new_AGEMA_signal_35797, new_AGEMA_signal_35794, new_AGEMA_signal_35791}), .clk (clk), .r ({Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300], Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296]}), .c ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_35812, new_AGEMA_signal_35809, new_AGEMA_signal_35806, new_AGEMA_signal_35803}), .clk (clk), .r ({Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310], Fresh[7309], Fresh[7308]}), .c ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_34923, new_AGEMA_signal_34919, new_AGEMA_signal_34915, new_AGEMA_signal_34911}), .clk (clk), .r ({Fresh[7331], Fresh[7330], Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320]}), .c ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_35824, new_AGEMA_signal_35821, new_AGEMA_signal_35818, new_AGEMA_signal_35815}), .clk (clk), .r ({Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340], Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332]}), .c ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_35836, new_AGEMA_signal_35833, new_AGEMA_signal_35830, new_AGEMA_signal_35827}), .clk (clk), .r ({Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350], Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344]}), .c ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_35848, new_AGEMA_signal_35845, new_AGEMA_signal_35842, new_AGEMA_signal_35839}), .clk (clk), .r ({Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360], Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356]}), .c ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_35860, new_AGEMA_signal_35857, new_AGEMA_signal_35854, new_AGEMA_signal_35851}), .clk (clk), .r ({Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370], Fresh[7369], Fresh[7368]}), .c ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_35872, new_AGEMA_signal_35869, new_AGEMA_signal_35866, new_AGEMA_signal_35863}), .clk (clk), .r ({Fresh[7391], Fresh[7390], Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380]}), .c ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_35884, new_AGEMA_signal_35881, new_AGEMA_signal_35878, new_AGEMA_signal_35875}), .clk (clk), .r ({Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400], Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392]}), .c ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, new_AGEMA_signal_10453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_35896, new_AGEMA_signal_35893, new_AGEMA_signal_35890, new_AGEMA_signal_35887}), .clk (clk), .r ({Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410], Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404]}), .c ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_35908, new_AGEMA_signal_35905, new_AGEMA_signal_35902, new_AGEMA_signal_35899}), .clk (clk), .r ({Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420], Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416]}), .c ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_35920, new_AGEMA_signal_35917, new_AGEMA_signal_35914, new_AGEMA_signal_35911}), .clk (clk), .r ({Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430], Fresh[7429], Fresh[7428]}), .c ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, new_AGEMA_signal_9748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_35932, new_AGEMA_signal_35929, new_AGEMA_signal_35926, new_AGEMA_signal_35923}), .clk (clk), .r ({Fresh[7451], Fresh[7450], Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440]}), .c ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_35944, new_AGEMA_signal_35941, new_AGEMA_signal_35938, new_AGEMA_signal_35935}), .clk (clk), .r ({Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460], Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452]}), .c ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_35956, new_AGEMA_signal_35953, new_AGEMA_signal_35950, new_AGEMA_signal_35947}), .clk (clk), .r ({Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470], Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464]}), .c ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, new_AGEMA_signal_9754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_35968, new_AGEMA_signal_35965, new_AGEMA_signal_35962, new_AGEMA_signal_35959}), .clk (clk), .r ({Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480], Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476]}), .c ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_35980, new_AGEMA_signal_35977, new_AGEMA_signal_35974, new_AGEMA_signal_35971}), .clk (clk), .r ({Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490], Fresh[7489], Fresh[7488]}), .c ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_35992, new_AGEMA_signal_35989, new_AGEMA_signal_35986, new_AGEMA_signal_35983}), .clk (clk), .r ({Fresh[7511], Fresh[7510], Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500]}), .c ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, new_AGEMA_signal_10453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, new_AGEMA_signal_11176, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, new_AGEMA_signal_11176, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, new_AGEMA_signal_9754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, new_AGEMA_signal_10474, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, new_AGEMA_signal_12301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, new_AGEMA_signal_11179, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, new_AGEMA_signal_11182, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, new_AGEMA_signal_12304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, new_AGEMA_signal_9748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, new_AGEMA_signal_11185, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, new_AGEMA_signal_11188, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, new_AGEMA_signal_12307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, new_AGEMA_signal_12310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, new_AGEMA_signal_10474, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, new_AGEMA_signal_11782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, new_AGEMA_signal_11188, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, new_AGEMA_signal_11182, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, new_AGEMA_signal_12313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12318, new_AGEMA_signal_12317, new_AGEMA_signal_12316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, new_AGEMA_signal_12319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, new_AGEMA_signal_12322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, new_AGEMA_signal_11179, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, new_AGEMA_signal_12325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, new_AGEMA_signal_11185, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_12330, new_AGEMA_signal_12329, new_AGEMA_signal_12328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, new_AGEMA_signal_12313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, new_AGEMA_signal_12973, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, new_AGEMA_signal_12304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, new_AGEMA_signal_12319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_12978, new_AGEMA_signal_12977, new_AGEMA_signal_12976, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, new_AGEMA_signal_12325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, new_AGEMA_signal_12979, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, new_AGEMA_signal_12310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_12984, new_AGEMA_signal_12983, new_AGEMA_signal_12982, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, new_AGEMA_signal_12307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, new_AGEMA_signal_11782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, new_AGEMA_signal_12985, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_12318, new_AGEMA_signal_12317, new_AGEMA_signal_12316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_12330, new_AGEMA_signal_12329, new_AGEMA_signal_12328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_12990, new_AGEMA_signal_12989, new_AGEMA_signal_12988, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, new_AGEMA_signal_12301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, new_AGEMA_signal_12322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, new_AGEMA_signal_12991, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, new_AGEMA_signal_12331, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_36004, new_AGEMA_signal_36001, new_AGEMA_signal_35998, new_AGEMA_signal_35995}), .clk (clk), .r ({Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520], Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512]}), .c ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_36016, new_AGEMA_signal_36013, new_AGEMA_signal_36010, new_AGEMA_signal_36007}), .clk (clk), .r ({Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530], Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524]}), .c ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_33739, new_AGEMA_signal_33735, new_AGEMA_signal_33731, new_AGEMA_signal_33727}), .clk (clk), .r ({Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540], Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536]}), .c ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_36028, new_AGEMA_signal_36025, new_AGEMA_signal_36022, new_AGEMA_signal_36019}), .clk (clk), .r ({Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550], Fresh[7549], Fresh[7548]}), .c ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_36040, new_AGEMA_signal_36037, new_AGEMA_signal_36034, new_AGEMA_signal_36031}), .clk (clk), .r ({Fresh[7571], Fresh[7570], Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560]}), .c ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_36052, new_AGEMA_signal_36049, new_AGEMA_signal_36046, new_AGEMA_signal_36043}), .clk (clk), .r ({Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580], Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572]}), .c ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_36064, new_AGEMA_signal_36061, new_AGEMA_signal_36058, new_AGEMA_signal_36055}), .clk (clk), .r ({Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590], Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584]}), .c ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_36076, new_AGEMA_signal_36073, new_AGEMA_signal_36070, new_AGEMA_signal_36067}), .clk (clk), .r ({Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600], Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596]}), .c ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_36088, new_AGEMA_signal_36085, new_AGEMA_signal_36082, new_AGEMA_signal_36079}), .clk (clk), .r ({Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610], Fresh[7609], Fresh[7608]}), .c ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_36100, new_AGEMA_signal_36097, new_AGEMA_signal_36094, new_AGEMA_signal_36091}), .clk (clk), .r ({Fresh[7631], Fresh[7630], Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620]}), .c ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_36112, new_AGEMA_signal_36109, new_AGEMA_signal_36106, new_AGEMA_signal_36103}), .clk (clk), .r ({Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640], Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632]}), .c ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_36124, new_AGEMA_signal_36121, new_AGEMA_signal_36118, new_AGEMA_signal_36115}), .clk (clk), .r ({Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650], Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644]}), .c ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, new_AGEMA_signal_9784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_36136, new_AGEMA_signal_36133, new_AGEMA_signal_36130, new_AGEMA_signal_36127}), .clk (clk), .r ({Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660], Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656]}), .c ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_36148, new_AGEMA_signal_36145, new_AGEMA_signal_36142, new_AGEMA_signal_36139}), .clk (clk), .r ({Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670], Fresh[7669], Fresh[7668]}), .c ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_36160, new_AGEMA_signal_36157, new_AGEMA_signal_36154, new_AGEMA_signal_36151}), .clk (clk), .r ({Fresh[7691], Fresh[7690], Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680]}), .c ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, new_AGEMA_signal_9790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_36172, new_AGEMA_signal_36169, new_AGEMA_signal_36166, new_AGEMA_signal_36163}), .clk (clk), .r ({Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700], Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692]}), .c ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_36184, new_AGEMA_signal_36181, new_AGEMA_signal_36178, new_AGEMA_signal_36175}), .clk (clk), .r ({Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710], Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704]}), .c ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_36196, new_AGEMA_signal_36193, new_AGEMA_signal_36190, new_AGEMA_signal_36187}), .clk (clk), .r ({Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720], Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716]}), .c ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, new_AGEMA_signal_11206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, new_AGEMA_signal_11206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, new_AGEMA_signal_9790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, new_AGEMA_signal_10510, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, new_AGEMA_signal_12334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, new_AGEMA_signal_11209, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11214, new_AGEMA_signal_11213, new_AGEMA_signal_11212, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, new_AGEMA_signal_12337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, new_AGEMA_signal_9784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, new_AGEMA_signal_11218, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, new_AGEMA_signal_11806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_12342, new_AGEMA_signal_12341, new_AGEMA_signal_12340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, new_AGEMA_signal_12343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, new_AGEMA_signal_10510, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, new_AGEMA_signal_11218, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, new_AGEMA_signal_11812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_11214, new_AGEMA_signal_11213, new_AGEMA_signal_11212, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, new_AGEMA_signal_12346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, new_AGEMA_signal_12349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12354, new_AGEMA_signal_12353, new_AGEMA_signal_12352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, new_AGEMA_signal_12355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, new_AGEMA_signal_11209, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, new_AGEMA_signal_12358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, new_AGEMA_signal_12361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, new_AGEMA_signal_12346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_12996, new_AGEMA_signal_12995, new_AGEMA_signal_12994, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, new_AGEMA_signal_12337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_12354, new_AGEMA_signal_12353, new_AGEMA_signal_12352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, new_AGEMA_signal_12997, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, new_AGEMA_signal_11806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, new_AGEMA_signal_12358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_13002, new_AGEMA_signal_13001, new_AGEMA_signal_13000, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, new_AGEMA_signal_12343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, new_AGEMA_signal_13003, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_12342, new_AGEMA_signal_12341, new_AGEMA_signal_12340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_13008, new_AGEMA_signal_13007, new_AGEMA_signal_13006, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, new_AGEMA_signal_12349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, new_AGEMA_signal_12361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, new_AGEMA_signal_13009, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, new_AGEMA_signal_12334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, new_AGEMA_signal_12355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_13014, new_AGEMA_signal_13013, new_AGEMA_signal_13012, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, new_AGEMA_signal_11812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_12366, new_AGEMA_signal_12365, new_AGEMA_signal_12364, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_36208, new_AGEMA_signal_36205, new_AGEMA_signal_36202, new_AGEMA_signal_36199}), .clk (clk), .r ({Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730], Fresh[7729], Fresh[7728]}), .c ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_36220, new_AGEMA_signal_36217, new_AGEMA_signal_36214, new_AGEMA_signal_36211}), .clk (clk), .r ({Fresh[7751], Fresh[7750], Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740]}), .c ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, new_AGEMA_signal_9805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_35707, new_AGEMA_signal_35703, new_AGEMA_signal_35699, new_AGEMA_signal_35695}), .clk (clk), .r ({Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760], Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752]}), .c ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_36232, new_AGEMA_signal_36229, new_AGEMA_signal_36226, new_AGEMA_signal_36223}), .clk (clk), .r ({Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770], Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764]}), .c ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_36244, new_AGEMA_signal_36241, new_AGEMA_signal_36238, new_AGEMA_signal_36235}), .clk (clk), .r ({Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780], Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776]}), .c ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_36256, new_AGEMA_signal_36253, new_AGEMA_signal_36250, new_AGEMA_signal_36247}), .clk (clk), .r ({Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790], Fresh[7789], Fresh[7788]}), .c ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_36268, new_AGEMA_signal_36265, new_AGEMA_signal_36262, new_AGEMA_signal_36259}), .clk (clk), .r ({Fresh[7811], Fresh[7810], Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800]}), .c ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_36280, new_AGEMA_signal_36277, new_AGEMA_signal_36274, new_AGEMA_signal_36271}), .clk (clk), .r ({Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820], Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812]}), .c ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_36292, new_AGEMA_signal_36289, new_AGEMA_signal_36286, new_AGEMA_signal_36283}), .clk (clk), .r ({Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830], Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824]}), .c ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, new_AGEMA_signal_10525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_36304, new_AGEMA_signal_36301, new_AGEMA_signal_36298, new_AGEMA_signal_36295}), .clk (clk), .r ({Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840], Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836]}), .c ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_36316, new_AGEMA_signal_36313, new_AGEMA_signal_36310, new_AGEMA_signal_36307}), .clk (clk), .r ({Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850], Fresh[7849], Fresh[7848]}), .c ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_36328, new_AGEMA_signal_36325, new_AGEMA_signal_36322, new_AGEMA_signal_36319}), .clk (clk), .r ({Fresh[7871], Fresh[7870], Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860]}), .c ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, new_AGEMA_signal_9820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_36340, new_AGEMA_signal_36337, new_AGEMA_signal_36334, new_AGEMA_signal_36331}), .clk (clk), .r ({Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880], Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872]}), .c ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_36352, new_AGEMA_signal_36349, new_AGEMA_signal_36346, new_AGEMA_signal_36343}), .clk (clk), .r ({Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890], Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884]}), .c ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, new_AGEMA_signal_9823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_36364, new_AGEMA_signal_36361, new_AGEMA_signal_36358, new_AGEMA_signal_36355}), .clk (clk), .r ({Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900], Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896]}), .c ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, new_AGEMA_signal_9826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_36376, new_AGEMA_signal_36373, new_AGEMA_signal_36370, new_AGEMA_signal_36367}), .clk (clk), .r ({Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910], Fresh[7909], Fresh[7908]}), .c ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_36388, new_AGEMA_signal_36385, new_AGEMA_signal_36382, new_AGEMA_signal_36379}), .clk (clk), .r ({Fresh[7931], Fresh[7930], Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920]}), .c ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_36400, new_AGEMA_signal_36397, new_AGEMA_signal_36394, new_AGEMA_signal_36391}), .clk (clk), .r ({Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940], Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932]}), .c ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, new_AGEMA_signal_10537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, new_AGEMA_signal_9805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, new_AGEMA_signal_10525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11238, new_AGEMA_signal_11237, new_AGEMA_signal_11236, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_11238, new_AGEMA_signal_11237, new_AGEMA_signal_11236, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, new_AGEMA_signal_9823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, new_AGEMA_signal_9826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, new_AGEMA_signal_10546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, new_AGEMA_signal_12367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, new_AGEMA_signal_11242, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, new_AGEMA_signal_12370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, new_AGEMA_signal_9820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, new_AGEMA_signal_11245, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_11250, new_AGEMA_signal_11249, new_AGEMA_signal_11248, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, new_AGEMA_signal_10537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, new_AGEMA_signal_11833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, new_AGEMA_signal_12373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_12378, new_AGEMA_signal_12377, new_AGEMA_signal_12376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, new_AGEMA_signal_10546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, new_AGEMA_signal_11836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_11250, new_AGEMA_signal_11249, new_AGEMA_signal_11248, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, new_AGEMA_signal_11839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, new_AGEMA_signal_11242, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, new_AGEMA_signal_12379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, new_AGEMA_signal_12382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, new_AGEMA_signal_12385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12390, new_AGEMA_signal_12389, new_AGEMA_signal_12388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, new_AGEMA_signal_12391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, new_AGEMA_signal_11245, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, new_AGEMA_signal_12394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, new_AGEMA_signal_12379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, new_AGEMA_signal_13015, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, new_AGEMA_signal_12370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, new_AGEMA_signal_12385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_13020, new_AGEMA_signal_13019, new_AGEMA_signal_13018, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, new_AGEMA_signal_11833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, new_AGEMA_signal_12391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, new_AGEMA_signal_13021, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12378, new_AGEMA_signal_12377, new_AGEMA_signal_12376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_13026, new_AGEMA_signal_13025, new_AGEMA_signal_13024, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, new_AGEMA_signal_12373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, new_AGEMA_signal_11836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, new_AGEMA_signal_13027, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, new_AGEMA_signal_12382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, new_AGEMA_signal_12394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_13032, new_AGEMA_signal_13031, new_AGEMA_signal_13030, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, new_AGEMA_signal_12367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_12390, new_AGEMA_signal_12389, new_AGEMA_signal_12388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, new_AGEMA_signal_13033, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, new_AGEMA_signal_11839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, new_AGEMA_signal_12397, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_36412, new_AGEMA_signal_36409, new_AGEMA_signal_36406, new_AGEMA_signal_36403}), .clk (clk), .r ({Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950], Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944]}), .c ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_36424, new_AGEMA_signal_36421, new_AGEMA_signal_36418, new_AGEMA_signal_36415}), .clk (clk), .r ({Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960], Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956]}), .c ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, new_AGEMA_signal_9841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_34475, new_AGEMA_signal_34471, new_AGEMA_signal_34467, new_AGEMA_signal_34463}), .clk (clk), .r ({Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970], Fresh[7969], Fresh[7968]}), .c ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_36436, new_AGEMA_signal_36433, new_AGEMA_signal_36430, new_AGEMA_signal_36427}), .clk (clk), .r ({Fresh[7991], Fresh[7990], Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980]}), .c ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, new_AGEMA_signal_10555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_36448, new_AGEMA_signal_36445, new_AGEMA_signal_36442, new_AGEMA_signal_36439}), .clk (clk), .r ({Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000], Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992]}), .c ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_36460, new_AGEMA_signal_36457, new_AGEMA_signal_36454, new_AGEMA_signal_36451}), .clk (clk), .r ({Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010], Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004]}), .c ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_36472, new_AGEMA_signal_36469, new_AGEMA_signal_36466, new_AGEMA_signal_36463}), .clk (clk), .r ({Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020], Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016]}), .c ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_36484, new_AGEMA_signal_36481, new_AGEMA_signal_36478, new_AGEMA_signal_36475}), .clk (clk), .r ({Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030], Fresh[8029], Fresh[8028]}), .c ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_36496, new_AGEMA_signal_36493, new_AGEMA_signal_36490, new_AGEMA_signal_36487}), .clk (clk), .r ({Fresh[8051], Fresh[8050], Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040]}), .c ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, new_AGEMA_signal_10561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_36508, new_AGEMA_signal_36505, new_AGEMA_signal_36502, new_AGEMA_signal_36499}), .clk (clk), .r ({Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060], Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052]}), .c ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_36520, new_AGEMA_signal_36517, new_AGEMA_signal_36514, new_AGEMA_signal_36511}), .clk (clk), .r ({Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070], Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064]}), .c ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_36532, new_AGEMA_signal_36529, new_AGEMA_signal_36526, new_AGEMA_signal_36523}), .clk (clk), .r ({Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080], Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076]}), .c ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, new_AGEMA_signal_9856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_36544, new_AGEMA_signal_36541, new_AGEMA_signal_36538, new_AGEMA_signal_36535}), .clk (clk), .r ({Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090], Fresh[8089], Fresh[8088]}), .c ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_36556, new_AGEMA_signal_36553, new_AGEMA_signal_36550, new_AGEMA_signal_36547}), .clk (clk), .r ({Fresh[8111], Fresh[8110], Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100]}), .c ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, new_AGEMA_signal_9859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_36568, new_AGEMA_signal_36565, new_AGEMA_signal_36562, new_AGEMA_signal_36559}), .clk (clk), .r ({Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120], Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112]}), .c ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, new_AGEMA_signal_9862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_36580, new_AGEMA_signal_36577, new_AGEMA_signal_36574, new_AGEMA_signal_36571}), .clk (clk), .r ({Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130], Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124]}), .c ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_36592, new_AGEMA_signal_36589, new_AGEMA_signal_36586, new_AGEMA_signal_36583}), .clk (clk), .r ({Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140], Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136]}), .c ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_36604, new_AGEMA_signal_36601, new_AGEMA_signal_36598, new_AGEMA_signal_36595}), .clk (clk), .r ({Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150], Fresh[8149], Fresh[8148]}), .c ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, new_AGEMA_signal_10573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, new_AGEMA_signal_9841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, new_AGEMA_signal_10561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, new_AGEMA_signal_10555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, new_AGEMA_signal_11266, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, new_AGEMA_signal_11266, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, new_AGEMA_signal_9859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, new_AGEMA_signal_9862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, new_AGEMA_signal_10582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12402, new_AGEMA_signal_12401, new_AGEMA_signal_12400, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, new_AGEMA_signal_11269, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11274, new_AGEMA_signal_11273, new_AGEMA_signal_11272, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, new_AGEMA_signal_12403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, new_AGEMA_signal_9856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, new_AGEMA_signal_11278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, new_AGEMA_signal_10573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, new_AGEMA_signal_11860, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, new_AGEMA_signal_12406, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, new_AGEMA_signal_12409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, new_AGEMA_signal_10582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, new_AGEMA_signal_11863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, new_AGEMA_signal_11278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, new_AGEMA_signal_11866, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_11274, new_AGEMA_signal_11273, new_AGEMA_signal_11272, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12414, new_AGEMA_signal_12413, new_AGEMA_signal_12412, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, new_AGEMA_signal_12415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, new_AGEMA_signal_12418, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, new_AGEMA_signal_12421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, new_AGEMA_signal_11269, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_12426, new_AGEMA_signal_12425, new_AGEMA_signal_12424, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, new_AGEMA_signal_12427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12414, new_AGEMA_signal_12413, new_AGEMA_signal_12412, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_13038, new_AGEMA_signal_13037, new_AGEMA_signal_13036, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, new_AGEMA_signal_12403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, new_AGEMA_signal_12418, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, new_AGEMA_signal_13039, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, new_AGEMA_signal_11860, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_12426, new_AGEMA_signal_12425, new_AGEMA_signal_12424, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_13044, new_AGEMA_signal_13043, new_AGEMA_signal_13042, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, new_AGEMA_signal_12409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, new_AGEMA_signal_13045, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, new_AGEMA_signal_12406, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, new_AGEMA_signal_11863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_13050, new_AGEMA_signal_13049, new_AGEMA_signal_13048, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, new_AGEMA_signal_12415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, new_AGEMA_signal_12427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, new_AGEMA_signal_13051, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_12402, new_AGEMA_signal_12401, new_AGEMA_signal_12400, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, new_AGEMA_signal_12421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_13056, new_AGEMA_signal_13055, new_AGEMA_signal_13054, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, new_AGEMA_signal_11866, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, new_AGEMA_signal_12430, KeyExpansionIns_tmp[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_26127), .Q (new_AGEMA_signal_26128) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_26131), .Q (new_AGEMA_signal_26132) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_26135), .Q (new_AGEMA_signal_26136) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_26139), .Q (new_AGEMA_signal_26140) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_26143), .Q (new_AGEMA_signal_26144) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_26147), .Q (new_AGEMA_signal_26148) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_26151), .Q (new_AGEMA_signal_26152) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_26155), .Q (new_AGEMA_signal_26156) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_26159), .Q (new_AGEMA_signal_26160) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_26163), .Q (new_AGEMA_signal_26164) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_26167), .Q (new_AGEMA_signal_26168) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_26171), .Q (new_AGEMA_signal_26172) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_26175), .Q (new_AGEMA_signal_26176) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_26179), .Q (new_AGEMA_signal_26180) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_26183), .Q (new_AGEMA_signal_26184) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_26187), .Q (new_AGEMA_signal_26188) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_26191), .Q (new_AGEMA_signal_26192) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_26195), .Q (new_AGEMA_signal_26196) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_26199), .Q (new_AGEMA_signal_26200) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_26203), .Q (new_AGEMA_signal_26204) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_26207), .Q (new_AGEMA_signal_26208) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_26211), .Q (new_AGEMA_signal_26212) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_26215), .Q (new_AGEMA_signal_26216) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_26219), .Q (new_AGEMA_signal_26220) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_26223), .Q (new_AGEMA_signal_26224) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_26227), .Q (new_AGEMA_signal_26228) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_26231), .Q (new_AGEMA_signal_26232) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_26235), .Q (new_AGEMA_signal_26236) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_26239), .Q (new_AGEMA_signal_26240) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_26243), .Q (new_AGEMA_signal_26244) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_26247), .Q (new_AGEMA_signal_26248) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_26251), .Q (new_AGEMA_signal_26252) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_26255), .Q (new_AGEMA_signal_26256) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_26259), .Q (new_AGEMA_signal_26260) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_26263), .Q (new_AGEMA_signal_26264) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_26267), .Q (new_AGEMA_signal_26268) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_26271), .Q (new_AGEMA_signal_26272) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_26275), .Q (new_AGEMA_signal_26276) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_26279), .Q (new_AGEMA_signal_26280) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_26283), .Q (new_AGEMA_signal_26284) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_26287), .Q (new_AGEMA_signal_26288) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_26291), .Q (new_AGEMA_signal_26292) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_26295), .Q (new_AGEMA_signal_26296) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_26299), .Q (new_AGEMA_signal_26300) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_26303), .Q (new_AGEMA_signal_26304) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_26307), .Q (new_AGEMA_signal_26308) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_26311), .Q (new_AGEMA_signal_26312) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_26315), .Q (new_AGEMA_signal_26316) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_26319), .Q (new_AGEMA_signal_26320) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_26323), .Q (new_AGEMA_signal_26324) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_26327), .Q (new_AGEMA_signal_26328) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_26331), .Q (new_AGEMA_signal_26332) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_26335), .Q (new_AGEMA_signal_26336) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_26339), .Q (new_AGEMA_signal_26340) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_26343), .Q (new_AGEMA_signal_26344) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_26347), .Q (new_AGEMA_signal_26348) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_26351), .Q (new_AGEMA_signal_26352) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_26355), .Q (new_AGEMA_signal_26356) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_26359), .Q (new_AGEMA_signal_26360) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_26363), .Q (new_AGEMA_signal_26364) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_26367), .Q (new_AGEMA_signal_26368) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_26371), .Q (new_AGEMA_signal_26372) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_26375), .Q (new_AGEMA_signal_26376) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_26379), .Q (new_AGEMA_signal_26380) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_26383), .Q (new_AGEMA_signal_26384) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_26387), .Q (new_AGEMA_signal_26388) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_26391), .Q (new_AGEMA_signal_26392) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_26395), .Q (new_AGEMA_signal_26396) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_26399), .Q (new_AGEMA_signal_26400) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_26403), .Q (new_AGEMA_signal_26404) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_26407), .Q (new_AGEMA_signal_26408) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_26411), .Q (new_AGEMA_signal_26412) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_26415), .Q (new_AGEMA_signal_26416) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_26419), .Q (new_AGEMA_signal_26420) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_26423), .Q (new_AGEMA_signal_26424) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_26427), .Q (new_AGEMA_signal_26428) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_26431), .Q (new_AGEMA_signal_26432) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_26435), .Q (new_AGEMA_signal_26436) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_26439), .Q (new_AGEMA_signal_26440) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_26443), .Q (new_AGEMA_signal_26444) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_26447), .Q (new_AGEMA_signal_26448) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_26451), .Q (new_AGEMA_signal_26452) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_26455), .Q (new_AGEMA_signal_26456) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_26459), .Q (new_AGEMA_signal_26460) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_26463), .Q (new_AGEMA_signal_26464) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_26467), .Q (new_AGEMA_signal_26468) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_26471), .Q (new_AGEMA_signal_26472) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_26475), .Q (new_AGEMA_signal_26476) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_26479), .Q (new_AGEMA_signal_26480) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_26483), .Q (new_AGEMA_signal_26484) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_26487), .Q (new_AGEMA_signal_26488) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_26491), .Q (new_AGEMA_signal_26492) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_26495), .Q (new_AGEMA_signal_26496) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_26499), .Q (new_AGEMA_signal_26500) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_26503), .Q (new_AGEMA_signal_26504) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_26507), .Q (new_AGEMA_signal_26508) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_26511), .Q (new_AGEMA_signal_26512) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_26515), .Q (new_AGEMA_signal_26516) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_26519), .Q (new_AGEMA_signal_26520) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_26523), .Q (new_AGEMA_signal_26524) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_26527), .Q (new_AGEMA_signal_26528) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_26531), .Q (new_AGEMA_signal_26532) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_26535), .Q (new_AGEMA_signal_26536) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_26539), .Q (new_AGEMA_signal_26540) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_26543), .Q (new_AGEMA_signal_26544) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_26547), .Q (new_AGEMA_signal_26548) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_26551), .Q (new_AGEMA_signal_26552) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_26555), .Q (new_AGEMA_signal_26556) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_26559), .Q (new_AGEMA_signal_26560) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_26563), .Q (new_AGEMA_signal_26564) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_26567), .Q (new_AGEMA_signal_26568) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_26571), .Q (new_AGEMA_signal_26572) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_26575), .Q (new_AGEMA_signal_26576) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_26579), .Q (new_AGEMA_signal_26580) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_26583), .Q (new_AGEMA_signal_26584) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_26587), .Q (new_AGEMA_signal_26588) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_26591), .Q (new_AGEMA_signal_26592) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_26595), .Q (new_AGEMA_signal_26596) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_26599), .Q (new_AGEMA_signal_26600) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_26603), .Q (new_AGEMA_signal_26604) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_26607), .Q (new_AGEMA_signal_26608) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_26611), .Q (new_AGEMA_signal_26612) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_26615), .Q (new_AGEMA_signal_26616) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_26619), .Q (new_AGEMA_signal_26620) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_26623), .Q (new_AGEMA_signal_26624) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_26627), .Q (new_AGEMA_signal_26628) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_26631), .Q (new_AGEMA_signal_26632) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_26635), .Q (new_AGEMA_signal_26636) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_26639), .Q (new_AGEMA_signal_26640) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_26643), .Q (new_AGEMA_signal_26644) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_26647), .Q (new_AGEMA_signal_26648) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_26651), .Q (new_AGEMA_signal_26652) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_26655), .Q (new_AGEMA_signal_26656) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_26659), .Q (new_AGEMA_signal_26660) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_26663), .Q (new_AGEMA_signal_26664) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_26667), .Q (new_AGEMA_signal_26668) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_26671), .Q (new_AGEMA_signal_26672) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_26675), .Q (new_AGEMA_signal_26676) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_26679), .Q (new_AGEMA_signal_26680) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_26683), .Q (new_AGEMA_signal_26684) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_26687), .Q (new_AGEMA_signal_26688) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_26691), .Q (new_AGEMA_signal_26692) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_26695), .Q (new_AGEMA_signal_26696) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_26699), .Q (new_AGEMA_signal_26700) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_26703), .Q (new_AGEMA_signal_26704) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_26707), .Q (new_AGEMA_signal_26708) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_26711), .Q (new_AGEMA_signal_26712) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_26715), .Q (new_AGEMA_signal_26716) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_26719), .Q (new_AGEMA_signal_26720) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_26723), .Q (new_AGEMA_signal_26724) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_26727), .Q (new_AGEMA_signal_26728) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_26731), .Q (new_AGEMA_signal_26732) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_26735), .Q (new_AGEMA_signal_26736) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_26739), .Q (new_AGEMA_signal_26740) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_26743), .Q (new_AGEMA_signal_26744) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_26747), .Q (new_AGEMA_signal_26748) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_26751), .Q (new_AGEMA_signal_26752) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_26755), .Q (new_AGEMA_signal_26756) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_26759), .Q (new_AGEMA_signal_26760) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_26763), .Q (new_AGEMA_signal_26764) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_26767), .Q (new_AGEMA_signal_26768) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_26771), .Q (new_AGEMA_signal_26772) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_26775), .Q (new_AGEMA_signal_26776) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_26779), .Q (new_AGEMA_signal_26780) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_26783), .Q (new_AGEMA_signal_26784) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_26787), .Q (new_AGEMA_signal_26788) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_26791), .Q (new_AGEMA_signal_26792) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_26795), .Q (new_AGEMA_signal_26796) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_26799), .Q (new_AGEMA_signal_26800) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_26803), .Q (new_AGEMA_signal_26804) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_26807), .Q (new_AGEMA_signal_26808) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_26811), .Q (new_AGEMA_signal_26812) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_26815), .Q (new_AGEMA_signal_26816) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_26819), .Q (new_AGEMA_signal_26820) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_26823), .Q (new_AGEMA_signal_26824) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_26827), .Q (new_AGEMA_signal_26828) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_26831), .Q (new_AGEMA_signal_26832) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_26835), .Q (new_AGEMA_signal_26836) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_26839), .Q (new_AGEMA_signal_26840) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_26843), .Q (new_AGEMA_signal_26844) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_26847), .Q (new_AGEMA_signal_26848) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_26851), .Q (new_AGEMA_signal_26852) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_26855), .Q (new_AGEMA_signal_26856) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_26859), .Q (new_AGEMA_signal_26860) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_26863), .Q (new_AGEMA_signal_26864) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_26867), .Q (new_AGEMA_signal_26868) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_26871), .Q (new_AGEMA_signal_26872) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_26875), .Q (new_AGEMA_signal_26876) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_26879), .Q (new_AGEMA_signal_26880) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_26883), .Q (new_AGEMA_signal_26884) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_26887), .Q (new_AGEMA_signal_26888) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_26891), .Q (new_AGEMA_signal_26892) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_26895), .Q (new_AGEMA_signal_26896) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_26899), .Q (new_AGEMA_signal_26900) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_26903), .Q (new_AGEMA_signal_26904) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_26907), .Q (new_AGEMA_signal_26908) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_26911), .Q (new_AGEMA_signal_26912) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_26915), .Q (new_AGEMA_signal_26916) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_26919), .Q (new_AGEMA_signal_26920) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_26923), .Q (new_AGEMA_signal_26924) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_26927), .Q (new_AGEMA_signal_26928) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_26931), .Q (new_AGEMA_signal_26932) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_26935), .Q (new_AGEMA_signal_26936) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_26939), .Q (new_AGEMA_signal_26940) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_26943), .Q (new_AGEMA_signal_26944) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_26947), .Q (new_AGEMA_signal_26948) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_26951), .Q (new_AGEMA_signal_26952) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_26955), .Q (new_AGEMA_signal_26956) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_26959), .Q (new_AGEMA_signal_26960) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_26963), .Q (new_AGEMA_signal_26964) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_26967), .Q (new_AGEMA_signal_26968) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_26971), .Q (new_AGEMA_signal_26972) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_26975), .Q (new_AGEMA_signal_26976) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_26979), .Q (new_AGEMA_signal_26980) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_26983), .Q (new_AGEMA_signal_26984) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_26987), .Q (new_AGEMA_signal_26988) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_26991), .Q (new_AGEMA_signal_26992) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_26995), .Q (new_AGEMA_signal_26996) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_26999), .Q (new_AGEMA_signal_27000) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_27003), .Q (new_AGEMA_signal_27004) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_27007), .Q (new_AGEMA_signal_27008) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_27011), .Q (new_AGEMA_signal_27012) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_27015), .Q (new_AGEMA_signal_27016) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_27019), .Q (new_AGEMA_signal_27020) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_27023), .Q (new_AGEMA_signal_27024) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_27027), .Q (new_AGEMA_signal_27028) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_27031), .Q (new_AGEMA_signal_27032) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_27035), .Q (new_AGEMA_signal_27036) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C (clk), .D (new_AGEMA_signal_27039), .Q (new_AGEMA_signal_27040) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_27043), .Q (new_AGEMA_signal_27044) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_27047), .Q (new_AGEMA_signal_27048) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_27051), .Q (new_AGEMA_signal_27052) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_27055), .Q (new_AGEMA_signal_27056) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_27059), .Q (new_AGEMA_signal_27060) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_27063), .Q (new_AGEMA_signal_27064) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_27067), .Q (new_AGEMA_signal_27068) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_27071), .Q (new_AGEMA_signal_27072) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_27075), .Q (new_AGEMA_signal_27076) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_27079), .Q (new_AGEMA_signal_27080) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_27083), .Q (new_AGEMA_signal_27084) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_27087), .Q (new_AGEMA_signal_27088) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_27091), .Q (new_AGEMA_signal_27092) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_27095), .Q (new_AGEMA_signal_27096) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_27099), .Q (new_AGEMA_signal_27100) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_27103), .Q (new_AGEMA_signal_27104) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_27107), .Q (new_AGEMA_signal_27108) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_27111), .Q (new_AGEMA_signal_27112) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_27115), .Q (new_AGEMA_signal_27116) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_27119), .Q (new_AGEMA_signal_27120) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_27123), .Q (new_AGEMA_signal_27124) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_27127), .Q (new_AGEMA_signal_27128) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_27131), .Q (new_AGEMA_signal_27132) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_27135), .Q (new_AGEMA_signal_27136) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_27139), .Q (new_AGEMA_signal_27140) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_27143), .Q (new_AGEMA_signal_27144) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C (clk), .D (new_AGEMA_signal_27147), .Q (new_AGEMA_signal_27148) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_27151), .Q (new_AGEMA_signal_27152) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_27155), .Q (new_AGEMA_signal_27156) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_27159), .Q (new_AGEMA_signal_27160) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_27163), .Q (new_AGEMA_signal_27164) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_27167), .Q (new_AGEMA_signal_27168) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_27171), .Q (new_AGEMA_signal_27172) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_27175), .Q (new_AGEMA_signal_27176) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_27179), .Q (new_AGEMA_signal_27180) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_27183), .Q (new_AGEMA_signal_27184) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_27187), .Q (new_AGEMA_signal_27188) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_27191), .Q (new_AGEMA_signal_27192) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_27195), .Q (new_AGEMA_signal_27196) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_27199), .Q (new_AGEMA_signal_27200) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_27203), .Q (new_AGEMA_signal_27204) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_27207), .Q (new_AGEMA_signal_27208) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_27211), .Q (new_AGEMA_signal_27212) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_27215), .Q (new_AGEMA_signal_27216) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_27219), .Q (new_AGEMA_signal_27220) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_27223), .Q (new_AGEMA_signal_27224) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_27227), .Q (new_AGEMA_signal_27228) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_27231), .Q (new_AGEMA_signal_27232) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_27235), .Q (new_AGEMA_signal_27236) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_27239), .Q (new_AGEMA_signal_27240) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_27243), .Q (new_AGEMA_signal_27244) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_27247), .Q (new_AGEMA_signal_27248) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_27251), .Q (new_AGEMA_signal_27252) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C (clk), .D (new_AGEMA_signal_27255), .Q (new_AGEMA_signal_27256) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_27259), .Q (new_AGEMA_signal_27260) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_27263), .Q (new_AGEMA_signal_27264) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_27267), .Q (new_AGEMA_signal_27268) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_27271), .Q (new_AGEMA_signal_27272) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_27275), .Q (new_AGEMA_signal_27276) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_27279), .Q (new_AGEMA_signal_27280) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_27283), .Q (new_AGEMA_signal_27284) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_27287), .Q (new_AGEMA_signal_27288) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_27291), .Q (new_AGEMA_signal_27292) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_27295), .Q (new_AGEMA_signal_27296) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_27299), .Q (new_AGEMA_signal_27300) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_27303), .Q (new_AGEMA_signal_27304) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_27307), .Q (new_AGEMA_signal_27308) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_27311), .Q (new_AGEMA_signal_27312) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_27315), .Q (new_AGEMA_signal_27316) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_27319), .Q (new_AGEMA_signal_27320) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_27323), .Q (new_AGEMA_signal_27324) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_27327), .Q (new_AGEMA_signal_27328) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_27331), .Q (new_AGEMA_signal_27332) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_27335), .Q (new_AGEMA_signal_27336) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_27339), .Q (new_AGEMA_signal_27340) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_27343), .Q (new_AGEMA_signal_27344) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_27347), .Q (new_AGEMA_signal_27348) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_27351), .Q (new_AGEMA_signal_27352) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_27355), .Q (new_AGEMA_signal_27356) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_27359), .Q (new_AGEMA_signal_27360) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C (clk), .D (new_AGEMA_signal_27363), .Q (new_AGEMA_signal_27364) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_27367), .Q (new_AGEMA_signal_27368) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_27371), .Q (new_AGEMA_signal_27372) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_27375), .Q (new_AGEMA_signal_27376) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_27379), .Q (new_AGEMA_signal_27380) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_27383), .Q (new_AGEMA_signal_27384) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_27387), .Q (new_AGEMA_signal_27388) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_27391), .Q (new_AGEMA_signal_27392) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_27395), .Q (new_AGEMA_signal_27396) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_27399), .Q (new_AGEMA_signal_27400) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_27403), .Q (new_AGEMA_signal_27404) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_27407), .Q (new_AGEMA_signal_27408) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_27411), .Q (new_AGEMA_signal_27412) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_27415), .Q (new_AGEMA_signal_27416) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_27419), .Q (new_AGEMA_signal_27420) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_27423), .Q (new_AGEMA_signal_27424) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_27427), .Q (new_AGEMA_signal_27428) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_27431), .Q (new_AGEMA_signal_27432) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_27435), .Q (new_AGEMA_signal_27436) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_27439), .Q (new_AGEMA_signal_27440) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_27443), .Q (new_AGEMA_signal_27444) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_27447), .Q (new_AGEMA_signal_27448) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_27451), .Q (new_AGEMA_signal_27452) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_27455), .Q (new_AGEMA_signal_27456) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_27459), .Q (new_AGEMA_signal_27460) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_27463), .Q (new_AGEMA_signal_27464) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_27467), .Q (new_AGEMA_signal_27468) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C (clk), .D (new_AGEMA_signal_27471), .Q (new_AGEMA_signal_27472) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_27475), .Q (new_AGEMA_signal_27476) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C (clk), .D (new_AGEMA_signal_27479), .Q (new_AGEMA_signal_27480) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_27483), .Q (new_AGEMA_signal_27484) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_27487), .Q (new_AGEMA_signal_27488) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_27491), .Q (new_AGEMA_signal_27492) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_27495), .Q (new_AGEMA_signal_27496) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_27499), .Q (new_AGEMA_signal_27500) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_27503), .Q (new_AGEMA_signal_27504) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_27507), .Q (new_AGEMA_signal_27508) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_27511), .Q (new_AGEMA_signal_27512) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C (clk), .D (new_AGEMA_signal_27515), .Q (new_AGEMA_signal_27516) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_27519), .Q (new_AGEMA_signal_27520) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_27523), .Q (new_AGEMA_signal_27524) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_27527), .Q (new_AGEMA_signal_27528) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_27531), .Q (new_AGEMA_signal_27532) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_27535), .Q (new_AGEMA_signal_27536) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_27539), .Q (new_AGEMA_signal_27540) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_27543), .Q (new_AGEMA_signal_27544) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_27547), .Q (new_AGEMA_signal_27548) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C (clk), .D (new_AGEMA_signal_27551), .Q (new_AGEMA_signal_27552) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_27555), .Q (new_AGEMA_signal_27556) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_27559), .Q (new_AGEMA_signal_27560) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_27563), .Q (new_AGEMA_signal_27564) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_27567), .Q (new_AGEMA_signal_27568) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_27571), .Q (new_AGEMA_signal_27572) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_27575), .Q (new_AGEMA_signal_27576) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C (clk), .D (new_AGEMA_signal_27579), .Q (new_AGEMA_signal_27580) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_27583), .Q (new_AGEMA_signal_27584) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C (clk), .D (new_AGEMA_signal_27587), .Q (new_AGEMA_signal_27588) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_27591), .Q (new_AGEMA_signal_27592) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_27595), .Q (new_AGEMA_signal_27596) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_27599), .Q (new_AGEMA_signal_27600) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_27603), .Q (new_AGEMA_signal_27604) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_27607), .Q (new_AGEMA_signal_27608) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_27611), .Q (new_AGEMA_signal_27612) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_27615), .Q (new_AGEMA_signal_27616) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_27619), .Q (new_AGEMA_signal_27620) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C (clk), .D (new_AGEMA_signal_27623), .Q (new_AGEMA_signal_27624) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_27627), .Q (new_AGEMA_signal_27628) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_27631), .Q (new_AGEMA_signal_27632) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C (clk), .D (new_AGEMA_signal_27635), .Q (new_AGEMA_signal_27636) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_27639), .Q (new_AGEMA_signal_27640) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C (clk), .D (new_AGEMA_signal_27643), .Q (new_AGEMA_signal_27644) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C (clk), .D (new_AGEMA_signal_27647), .Q (new_AGEMA_signal_27648) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C (clk), .D (new_AGEMA_signal_27651), .Q (new_AGEMA_signal_27652) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C (clk), .D (new_AGEMA_signal_27655), .Q (new_AGEMA_signal_27656) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C (clk), .D (new_AGEMA_signal_27659), .Q (new_AGEMA_signal_27660) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C (clk), .D (new_AGEMA_signal_27663), .Q (new_AGEMA_signal_27664) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C (clk), .D (new_AGEMA_signal_27667), .Q (new_AGEMA_signal_27668) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C (clk), .D (new_AGEMA_signal_27671), .Q (new_AGEMA_signal_27672) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C (clk), .D (new_AGEMA_signal_27675), .Q (new_AGEMA_signal_27676) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C (clk), .D (new_AGEMA_signal_27679), .Q (new_AGEMA_signal_27680) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C (clk), .D (new_AGEMA_signal_27683), .Q (new_AGEMA_signal_27684) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C (clk), .D (new_AGEMA_signal_27687), .Q (new_AGEMA_signal_27688) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C (clk), .D (new_AGEMA_signal_27691), .Q (new_AGEMA_signal_27692) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C (clk), .D (new_AGEMA_signal_27695), .Q (new_AGEMA_signal_27696) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C (clk), .D (new_AGEMA_signal_27699), .Q (new_AGEMA_signal_27700) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C (clk), .D (new_AGEMA_signal_27703), .Q (new_AGEMA_signal_27704) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C (clk), .D (new_AGEMA_signal_27707), .Q (new_AGEMA_signal_27708) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C (clk), .D (new_AGEMA_signal_27711), .Q (new_AGEMA_signal_27712) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C (clk), .D (new_AGEMA_signal_27715), .Q (new_AGEMA_signal_27716) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C (clk), .D (new_AGEMA_signal_27719), .Q (new_AGEMA_signal_27720) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C (clk), .D (new_AGEMA_signal_27723), .Q (new_AGEMA_signal_27724) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C (clk), .D (new_AGEMA_signal_27727), .Q (new_AGEMA_signal_27728) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C (clk), .D (new_AGEMA_signal_27731), .Q (new_AGEMA_signal_27732) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C (clk), .D (new_AGEMA_signal_27735), .Q (new_AGEMA_signal_27736) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C (clk), .D (new_AGEMA_signal_27739), .Q (new_AGEMA_signal_27740) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C (clk), .D (new_AGEMA_signal_27743), .Q (new_AGEMA_signal_27744) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C (clk), .D (new_AGEMA_signal_27747), .Q (new_AGEMA_signal_27748) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C (clk), .D (new_AGEMA_signal_27751), .Q (new_AGEMA_signal_27752) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C (clk), .D (new_AGEMA_signal_27755), .Q (new_AGEMA_signal_27756) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C (clk), .D (new_AGEMA_signal_27759), .Q (new_AGEMA_signal_27760) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C (clk), .D (new_AGEMA_signal_27763), .Q (new_AGEMA_signal_27764) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C (clk), .D (new_AGEMA_signal_27767), .Q (new_AGEMA_signal_27768) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C (clk), .D (new_AGEMA_signal_27771), .Q (new_AGEMA_signal_27772) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C (clk), .D (new_AGEMA_signal_27775), .Q (new_AGEMA_signal_27776) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C (clk), .D (new_AGEMA_signal_27779), .Q (new_AGEMA_signal_27780) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C (clk), .D (new_AGEMA_signal_27783), .Q (new_AGEMA_signal_27784) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C (clk), .D (new_AGEMA_signal_27787), .Q (new_AGEMA_signal_27788) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C (clk), .D (new_AGEMA_signal_27791), .Q (new_AGEMA_signal_27792) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C (clk), .D (new_AGEMA_signal_27795), .Q (new_AGEMA_signal_27796) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C (clk), .D (new_AGEMA_signal_27799), .Q (new_AGEMA_signal_27800) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C (clk), .D (new_AGEMA_signal_27803), .Q (new_AGEMA_signal_27804) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C (clk), .D (new_AGEMA_signal_27807), .Q (new_AGEMA_signal_27808) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C (clk), .D (new_AGEMA_signal_27811), .Q (new_AGEMA_signal_27812) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C (clk), .D (new_AGEMA_signal_27815), .Q (new_AGEMA_signal_27816) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C (clk), .D (new_AGEMA_signal_27819), .Q (new_AGEMA_signal_27820) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C (clk), .D (new_AGEMA_signal_27823), .Q (new_AGEMA_signal_27824) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C (clk), .D (new_AGEMA_signal_27827), .Q (new_AGEMA_signal_27828) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C (clk), .D (new_AGEMA_signal_27831), .Q (new_AGEMA_signal_27832) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C (clk), .D (new_AGEMA_signal_27835), .Q (new_AGEMA_signal_27836) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C (clk), .D (new_AGEMA_signal_27839), .Q (new_AGEMA_signal_27840) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C (clk), .D (new_AGEMA_signal_27843), .Q (new_AGEMA_signal_27844) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C (clk), .D (new_AGEMA_signal_27847), .Q (new_AGEMA_signal_27848) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C (clk), .D (new_AGEMA_signal_27851), .Q (new_AGEMA_signal_27852) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C (clk), .D (new_AGEMA_signal_27855), .Q (new_AGEMA_signal_27856) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C (clk), .D (new_AGEMA_signal_27859), .Q (new_AGEMA_signal_27860) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C (clk), .D (new_AGEMA_signal_27863), .Q (new_AGEMA_signal_27864) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C (clk), .D (new_AGEMA_signal_27867), .Q (new_AGEMA_signal_27868) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C (clk), .D (new_AGEMA_signal_27871), .Q (new_AGEMA_signal_27872) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C (clk), .D (new_AGEMA_signal_27875), .Q (new_AGEMA_signal_27876) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C (clk), .D (new_AGEMA_signal_27879), .Q (new_AGEMA_signal_27880) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C (clk), .D (new_AGEMA_signal_27883), .Q (new_AGEMA_signal_27884) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C (clk), .D (new_AGEMA_signal_27887), .Q (new_AGEMA_signal_27888) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C (clk), .D (new_AGEMA_signal_27891), .Q (new_AGEMA_signal_27892) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C (clk), .D (new_AGEMA_signal_27895), .Q (new_AGEMA_signal_27896) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C (clk), .D (new_AGEMA_signal_27899), .Q (new_AGEMA_signal_27900) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C (clk), .D (new_AGEMA_signal_27903), .Q (new_AGEMA_signal_27904) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C (clk), .D (new_AGEMA_signal_27907), .Q (new_AGEMA_signal_27908) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C (clk), .D (new_AGEMA_signal_27911), .Q (new_AGEMA_signal_27912) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C (clk), .D (new_AGEMA_signal_27915), .Q (new_AGEMA_signal_27916) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C (clk), .D (new_AGEMA_signal_27919), .Q (new_AGEMA_signal_27920) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C (clk), .D (new_AGEMA_signal_27923), .Q (new_AGEMA_signal_27924) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C (clk), .D (new_AGEMA_signal_27927), .Q (new_AGEMA_signal_27928) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C (clk), .D (new_AGEMA_signal_27931), .Q (new_AGEMA_signal_27932) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C (clk), .D (new_AGEMA_signal_27935), .Q (new_AGEMA_signal_27936) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C (clk), .D (new_AGEMA_signal_27939), .Q (new_AGEMA_signal_27940) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C (clk), .D (new_AGEMA_signal_27943), .Q (new_AGEMA_signal_27944) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C (clk), .D (new_AGEMA_signal_27947), .Q (new_AGEMA_signal_27948) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C (clk), .D (new_AGEMA_signal_27951), .Q (new_AGEMA_signal_27952) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C (clk), .D (new_AGEMA_signal_27955), .Q (new_AGEMA_signal_27956) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C (clk), .D (new_AGEMA_signal_27959), .Q (new_AGEMA_signal_27960) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C (clk), .D (new_AGEMA_signal_27963), .Q (new_AGEMA_signal_27964) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C (clk), .D (new_AGEMA_signal_27967), .Q (new_AGEMA_signal_27968) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C (clk), .D (new_AGEMA_signal_27971), .Q (new_AGEMA_signal_27972) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C (clk), .D (new_AGEMA_signal_27975), .Q (new_AGEMA_signal_27976) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C (clk), .D (new_AGEMA_signal_27979), .Q (new_AGEMA_signal_27980) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C (clk), .D (new_AGEMA_signal_27983), .Q (new_AGEMA_signal_27984) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C (clk), .D (new_AGEMA_signal_27987), .Q (new_AGEMA_signal_27988) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C (clk), .D (new_AGEMA_signal_27991), .Q (new_AGEMA_signal_27992) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C (clk), .D (new_AGEMA_signal_27995), .Q (new_AGEMA_signal_27996) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C (clk), .D (new_AGEMA_signal_27999), .Q (new_AGEMA_signal_28000) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C (clk), .D (new_AGEMA_signal_28003), .Q (new_AGEMA_signal_28004) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C (clk), .D (new_AGEMA_signal_28007), .Q (new_AGEMA_signal_28008) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C (clk), .D (new_AGEMA_signal_28011), .Q (new_AGEMA_signal_28012) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C (clk), .D (new_AGEMA_signal_28015), .Q (new_AGEMA_signal_28016) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C (clk), .D (new_AGEMA_signal_28019), .Q (new_AGEMA_signal_28020) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C (clk), .D (new_AGEMA_signal_28023), .Q (new_AGEMA_signal_28024) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C (clk), .D (new_AGEMA_signal_28027), .Q (new_AGEMA_signal_28028) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C (clk), .D (new_AGEMA_signal_28031), .Q (new_AGEMA_signal_28032) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C (clk), .D (new_AGEMA_signal_28035), .Q (new_AGEMA_signal_28036) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C (clk), .D (new_AGEMA_signal_28039), .Q (new_AGEMA_signal_28040) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C (clk), .D (new_AGEMA_signal_28043), .Q (new_AGEMA_signal_28044) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C (clk), .D (new_AGEMA_signal_28047), .Q (new_AGEMA_signal_28048) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C (clk), .D (new_AGEMA_signal_28051), .Q (new_AGEMA_signal_28052) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C (clk), .D (new_AGEMA_signal_28055), .Q (new_AGEMA_signal_28056) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C (clk), .D (new_AGEMA_signal_28059), .Q (new_AGEMA_signal_28060) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C (clk), .D (new_AGEMA_signal_28063), .Q (new_AGEMA_signal_28064) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C (clk), .D (new_AGEMA_signal_28067), .Q (new_AGEMA_signal_28068) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C (clk), .D (new_AGEMA_signal_28071), .Q (new_AGEMA_signal_28072) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C (clk), .D (new_AGEMA_signal_28075), .Q (new_AGEMA_signal_28076) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C (clk), .D (new_AGEMA_signal_28079), .Q (new_AGEMA_signal_28080) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C (clk), .D (new_AGEMA_signal_28083), .Q (new_AGEMA_signal_28084) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C (clk), .D (new_AGEMA_signal_28087), .Q (new_AGEMA_signal_28088) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C (clk), .D (new_AGEMA_signal_28091), .Q (new_AGEMA_signal_28092) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C (clk), .D (new_AGEMA_signal_28095), .Q (new_AGEMA_signal_28096) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C (clk), .D (new_AGEMA_signal_28099), .Q (new_AGEMA_signal_28100) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C (clk), .D (new_AGEMA_signal_28103), .Q (new_AGEMA_signal_28104) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C (clk), .D (new_AGEMA_signal_28107), .Q (new_AGEMA_signal_28108) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C (clk), .D (new_AGEMA_signal_28111), .Q (new_AGEMA_signal_28112) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C (clk), .D (new_AGEMA_signal_28115), .Q (new_AGEMA_signal_28116) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C (clk), .D (new_AGEMA_signal_28119), .Q (new_AGEMA_signal_28120) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C (clk), .D (new_AGEMA_signal_28123), .Q (new_AGEMA_signal_28124) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C (clk), .D (new_AGEMA_signal_28127), .Q (new_AGEMA_signal_28128) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C (clk), .D (new_AGEMA_signal_28131), .Q (new_AGEMA_signal_28132) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C (clk), .D (new_AGEMA_signal_28135), .Q (new_AGEMA_signal_28136) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C (clk), .D (new_AGEMA_signal_28139), .Q (new_AGEMA_signal_28140) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C (clk), .D (new_AGEMA_signal_28143), .Q (new_AGEMA_signal_28144) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C (clk), .D (new_AGEMA_signal_28147), .Q (new_AGEMA_signal_28148) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C (clk), .D (new_AGEMA_signal_28151), .Q (new_AGEMA_signal_28152) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C (clk), .D (new_AGEMA_signal_28155), .Q (new_AGEMA_signal_28156) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C (clk), .D (new_AGEMA_signal_28159), .Q (new_AGEMA_signal_28160) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C (clk), .D (new_AGEMA_signal_28163), .Q (new_AGEMA_signal_28164) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C (clk), .D (new_AGEMA_signal_28167), .Q (new_AGEMA_signal_28168) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C (clk), .D (new_AGEMA_signal_28171), .Q (new_AGEMA_signal_28172) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C (clk), .D (new_AGEMA_signal_28175), .Q (new_AGEMA_signal_28176) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C (clk), .D (new_AGEMA_signal_28179), .Q (new_AGEMA_signal_28180) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C (clk), .D (new_AGEMA_signal_28183), .Q (new_AGEMA_signal_28184) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C (clk), .D (new_AGEMA_signal_28187), .Q (new_AGEMA_signal_28188) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C (clk), .D (new_AGEMA_signal_28191), .Q (new_AGEMA_signal_28192) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C (clk), .D (new_AGEMA_signal_28195), .Q (new_AGEMA_signal_28196) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C (clk), .D (new_AGEMA_signal_28199), .Q (new_AGEMA_signal_28200) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C (clk), .D (new_AGEMA_signal_28203), .Q (new_AGEMA_signal_28204) ) ;
    buf_clk new_AGEMA_reg_buffer_10708 ( .C (clk), .D (new_AGEMA_signal_31663), .Q (new_AGEMA_signal_31664) ) ;
    buf_clk new_AGEMA_reg_buffer_10712 ( .C (clk), .D (new_AGEMA_signal_31667), .Q (new_AGEMA_signal_31668) ) ;
    buf_clk new_AGEMA_reg_buffer_10716 ( .C (clk), .D (new_AGEMA_signal_31671), .Q (new_AGEMA_signal_31672) ) ;
    buf_clk new_AGEMA_reg_buffer_10720 ( .C (clk), .D (new_AGEMA_signal_31675), .Q (new_AGEMA_signal_31676) ) ;
    buf_clk new_AGEMA_reg_buffer_10724 ( .C (clk), .D (new_AGEMA_signal_31679), .Q (new_AGEMA_signal_31680) ) ;
    buf_clk new_AGEMA_reg_buffer_10728 ( .C (clk), .D (new_AGEMA_signal_31683), .Q (new_AGEMA_signal_31684) ) ;
    buf_clk new_AGEMA_reg_buffer_10732 ( .C (clk), .D (new_AGEMA_signal_31687), .Q (new_AGEMA_signal_31688) ) ;
    buf_clk new_AGEMA_reg_buffer_10736 ( .C (clk), .D (new_AGEMA_signal_31691), .Q (new_AGEMA_signal_31692) ) ;
    buf_clk new_AGEMA_reg_buffer_10740 ( .C (clk), .D (new_AGEMA_signal_31695), .Q (new_AGEMA_signal_31696) ) ;
    buf_clk new_AGEMA_reg_buffer_10744 ( .C (clk), .D (new_AGEMA_signal_31699), .Q (new_AGEMA_signal_31700) ) ;
    buf_clk new_AGEMA_reg_buffer_10748 ( .C (clk), .D (new_AGEMA_signal_31703), .Q (new_AGEMA_signal_31704) ) ;
    buf_clk new_AGEMA_reg_buffer_10752 ( .C (clk), .D (new_AGEMA_signal_31707), .Q (new_AGEMA_signal_31708) ) ;
    buf_clk new_AGEMA_reg_buffer_10756 ( .C (clk), .D (new_AGEMA_signal_31711), .Q (new_AGEMA_signal_31712) ) ;
    buf_clk new_AGEMA_reg_buffer_10760 ( .C (clk), .D (new_AGEMA_signal_31715), .Q (new_AGEMA_signal_31716) ) ;
    buf_clk new_AGEMA_reg_buffer_10764 ( .C (clk), .D (new_AGEMA_signal_31719), .Q (new_AGEMA_signal_31720) ) ;
    buf_clk new_AGEMA_reg_buffer_10768 ( .C (clk), .D (new_AGEMA_signal_31723), .Q (new_AGEMA_signal_31724) ) ;
    buf_clk new_AGEMA_reg_buffer_10772 ( .C (clk), .D (new_AGEMA_signal_31727), .Q (new_AGEMA_signal_31728) ) ;
    buf_clk new_AGEMA_reg_buffer_10776 ( .C (clk), .D (new_AGEMA_signal_31731), .Q (new_AGEMA_signal_31732) ) ;
    buf_clk new_AGEMA_reg_buffer_10780 ( .C (clk), .D (new_AGEMA_signal_31735), .Q (new_AGEMA_signal_31736) ) ;
    buf_clk new_AGEMA_reg_buffer_10784 ( .C (clk), .D (new_AGEMA_signal_31739), .Q (new_AGEMA_signal_31740) ) ;
    buf_clk new_AGEMA_reg_buffer_10788 ( .C (clk), .D (new_AGEMA_signal_31743), .Q (new_AGEMA_signal_31744) ) ;
    buf_clk new_AGEMA_reg_buffer_10792 ( .C (clk), .D (new_AGEMA_signal_31747), .Q (new_AGEMA_signal_31748) ) ;
    buf_clk new_AGEMA_reg_buffer_10796 ( .C (clk), .D (new_AGEMA_signal_31751), .Q (new_AGEMA_signal_31752) ) ;
    buf_clk new_AGEMA_reg_buffer_10800 ( .C (clk), .D (new_AGEMA_signal_31755), .Q (new_AGEMA_signal_31756) ) ;
    buf_clk new_AGEMA_reg_buffer_10804 ( .C (clk), .D (new_AGEMA_signal_31759), .Q (new_AGEMA_signal_31760) ) ;
    buf_clk new_AGEMA_reg_buffer_10808 ( .C (clk), .D (new_AGEMA_signal_31763), .Q (new_AGEMA_signal_31764) ) ;
    buf_clk new_AGEMA_reg_buffer_10812 ( .C (clk), .D (new_AGEMA_signal_31767), .Q (new_AGEMA_signal_31768) ) ;
    buf_clk new_AGEMA_reg_buffer_10816 ( .C (clk), .D (new_AGEMA_signal_31771), .Q (new_AGEMA_signal_31772) ) ;
    buf_clk new_AGEMA_reg_buffer_10820 ( .C (clk), .D (new_AGEMA_signal_31775), .Q (new_AGEMA_signal_31776) ) ;
    buf_clk new_AGEMA_reg_buffer_10824 ( .C (clk), .D (new_AGEMA_signal_31779), .Q (new_AGEMA_signal_31780) ) ;
    buf_clk new_AGEMA_reg_buffer_10828 ( .C (clk), .D (new_AGEMA_signal_31783), .Q (new_AGEMA_signal_31784) ) ;
    buf_clk new_AGEMA_reg_buffer_10832 ( .C (clk), .D (new_AGEMA_signal_31787), .Q (new_AGEMA_signal_31788) ) ;
    buf_clk new_AGEMA_reg_buffer_10836 ( .C (clk), .D (new_AGEMA_signal_31791), .Q (new_AGEMA_signal_31792) ) ;
    buf_clk new_AGEMA_reg_buffer_10840 ( .C (clk), .D (new_AGEMA_signal_31795), .Q (new_AGEMA_signal_31796) ) ;
    buf_clk new_AGEMA_reg_buffer_10844 ( .C (clk), .D (new_AGEMA_signal_31799), .Q (new_AGEMA_signal_31800) ) ;
    buf_clk new_AGEMA_reg_buffer_10848 ( .C (clk), .D (new_AGEMA_signal_31803), .Q (new_AGEMA_signal_31804) ) ;
    buf_clk new_AGEMA_reg_buffer_10852 ( .C (clk), .D (new_AGEMA_signal_31807), .Q (new_AGEMA_signal_31808) ) ;
    buf_clk new_AGEMA_reg_buffer_10856 ( .C (clk), .D (new_AGEMA_signal_31811), .Q (new_AGEMA_signal_31812) ) ;
    buf_clk new_AGEMA_reg_buffer_10860 ( .C (clk), .D (new_AGEMA_signal_31815), .Q (new_AGEMA_signal_31816) ) ;
    buf_clk new_AGEMA_reg_buffer_10864 ( .C (clk), .D (new_AGEMA_signal_31819), .Q (new_AGEMA_signal_31820) ) ;
    buf_clk new_AGEMA_reg_buffer_10868 ( .C (clk), .D (new_AGEMA_signal_31823), .Q (new_AGEMA_signal_31824) ) ;
    buf_clk new_AGEMA_reg_buffer_10872 ( .C (clk), .D (new_AGEMA_signal_31827), .Q (new_AGEMA_signal_31828) ) ;
    buf_clk new_AGEMA_reg_buffer_10876 ( .C (clk), .D (new_AGEMA_signal_31831), .Q (new_AGEMA_signal_31832) ) ;
    buf_clk new_AGEMA_reg_buffer_10880 ( .C (clk), .D (new_AGEMA_signal_31835), .Q (new_AGEMA_signal_31836) ) ;
    buf_clk new_AGEMA_reg_buffer_10884 ( .C (clk), .D (new_AGEMA_signal_31839), .Q (new_AGEMA_signal_31840) ) ;
    buf_clk new_AGEMA_reg_buffer_10888 ( .C (clk), .D (new_AGEMA_signal_31843), .Q (new_AGEMA_signal_31844) ) ;
    buf_clk new_AGEMA_reg_buffer_10892 ( .C (clk), .D (new_AGEMA_signal_31847), .Q (new_AGEMA_signal_31848) ) ;
    buf_clk new_AGEMA_reg_buffer_10896 ( .C (clk), .D (new_AGEMA_signal_31851), .Q (new_AGEMA_signal_31852) ) ;
    buf_clk new_AGEMA_reg_buffer_10900 ( .C (clk), .D (new_AGEMA_signal_31855), .Q (new_AGEMA_signal_31856) ) ;
    buf_clk new_AGEMA_reg_buffer_10904 ( .C (clk), .D (new_AGEMA_signal_31859), .Q (new_AGEMA_signal_31860) ) ;
    buf_clk new_AGEMA_reg_buffer_10908 ( .C (clk), .D (new_AGEMA_signal_31863), .Q (new_AGEMA_signal_31864) ) ;
    buf_clk new_AGEMA_reg_buffer_10912 ( .C (clk), .D (new_AGEMA_signal_31867), .Q (new_AGEMA_signal_31868) ) ;
    buf_clk new_AGEMA_reg_buffer_10916 ( .C (clk), .D (new_AGEMA_signal_31871), .Q (new_AGEMA_signal_31872) ) ;
    buf_clk new_AGEMA_reg_buffer_10920 ( .C (clk), .D (new_AGEMA_signal_31875), .Q (new_AGEMA_signal_31876) ) ;
    buf_clk new_AGEMA_reg_buffer_10924 ( .C (clk), .D (new_AGEMA_signal_31879), .Q (new_AGEMA_signal_31880) ) ;
    buf_clk new_AGEMA_reg_buffer_10928 ( .C (clk), .D (new_AGEMA_signal_31883), .Q (new_AGEMA_signal_31884) ) ;
    buf_clk new_AGEMA_reg_buffer_10932 ( .C (clk), .D (new_AGEMA_signal_31887), .Q (new_AGEMA_signal_31888) ) ;
    buf_clk new_AGEMA_reg_buffer_10936 ( .C (clk), .D (new_AGEMA_signal_31891), .Q (new_AGEMA_signal_31892) ) ;
    buf_clk new_AGEMA_reg_buffer_10940 ( .C (clk), .D (new_AGEMA_signal_31895), .Q (new_AGEMA_signal_31896) ) ;
    buf_clk new_AGEMA_reg_buffer_10944 ( .C (clk), .D (new_AGEMA_signal_31899), .Q (new_AGEMA_signal_31900) ) ;
    buf_clk new_AGEMA_reg_buffer_10948 ( .C (clk), .D (new_AGEMA_signal_31903), .Q (new_AGEMA_signal_31904) ) ;
    buf_clk new_AGEMA_reg_buffer_10952 ( .C (clk), .D (new_AGEMA_signal_31907), .Q (new_AGEMA_signal_31908) ) ;
    buf_clk new_AGEMA_reg_buffer_10956 ( .C (clk), .D (new_AGEMA_signal_31911), .Q (new_AGEMA_signal_31912) ) ;
    buf_clk new_AGEMA_reg_buffer_10960 ( .C (clk), .D (new_AGEMA_signal_31915), .Q (new_AGEMA_signal_31916) ) ;
    buf_clk new_AGEMA_reg_buffer_10964 ( .C (clk), .D (new_AGEMA_signal_31919), .Q (new_AGEMA_signal_31920) ) ;
    buf_clk new_AGEMA_reg_buffer_10968 ( .C (clk), .D (new_AGEMA_signal_31923), .Q (new_AGEMA_signal_31924) ) ;
    buf_clk new_AGEMA_reg_buffer_10972 ( .C (clk), .D (new_AGEMA_signal_31927), .Q (new_AGEMA_signal_31928) ) ;
    buf_clk new_AGEMA_reg_buffer_10976 ( .C (clk), .D (new_AGEMA_signal_31931), .Q (new_AGEMA_signal_31932) ) ;
    buf_clk new_AGEMA_reg_buffer_10980 ( .C (clk), .D (new_AGEMA_signal_31935), .Q (new_AGEMA_signal_31936) ) ;
    buf_clk new_AGEMA_reg_buffer_10984 ( .C (clk), .D (new_AGEMA_signal_31939), .Q (new_AGEMA_signal_31940) ) ;
    buf_clk new_AGEMA_reg_buffer_10988 ( .C (clk), .D (new_AGEMA_signal_31943), .Q (new_AGEMA_signal_31944) ) ;
    buf_clk new_AGEMA_reg_buffer_10992 ( .C (clk), .D (new_AGEMA_signal_31947), .Q (new_AGEMA_signal_31948) ) ;
    buf_clk new_AGEMA_reg_buffer_10996 ( .C (clk), .D (new_AGEMA_signal_31951), .Q (new_AGEMA_signal_31952) ) ;
    buf_clk new_AGEMA_reg_buffer_11000 ( .C (clk), .D (new_AGEMA_signal_31955), .Q (new_AGEMA_signal_31956) ) ;
    buf_clk new_AGEMA_reg_buffer_11004 ( .C (clk), .D (new_AGEMA_signal_31959), .Q (new_AGEMA_signal_31960) ) ;
    buf_clk new_AGEMA_reg_buffer_11008 ( .C (clk), .D (new_AGEMA_signal_31963), .Q (new_AGEMA_signal_31964) ) ;
    buf_clk new_AGEMA_reg_buffer_11012 ( .C (clk), .D (new_AGEMA_signal_31967), .Q (new_AGEMA_signal_31968) ) ;
    buf_clk new_AGEMA_reg_buffer_11016 ( .C (clk), .D (new_AGEMA_signal_31971), .Q (new_AGEMA_signal_31972) ) ;
    buf_clk new_AGEMA_reg_buffer_11020 ( .C (clk), .D (new_AGEMA_signal_31975), .Q (new_AGEMA_signal_31976) ) ;
    buf_clk new_AGEMA_reg_buffer_11024 ( .C (clk), .D (new_AGEMA_signal_31979), .Q (new_AGEMA_signal_31980) ) ;
    buf_clk new_AGEMA_reg_buffer_11028 ( .C (clk), .D (new_AGEMA_signal_31983), .Q (new_AGEMA_signal_31984) ) ;
    buf_clk new_AGEMA_reg_buffer_11032 ( .C (clk), .D (new_AGEMA_signal_31987), .Q (new_AGEMA_signal_31988) ) ;
    buf_clk new_AGEMA_reg_buffer_11036 ( .C (clk), .D (new_AGEMA_signal_31991), .Q (new_AGEMA_signal_31992) ) ;
    buf_clk new_AGEMA_reg_buffer_11040 ( .C (clk), .D (new_AGEMA_signal_31995), .Q (new_AGEMA_signal_31996) ) ;
    buf_clk new_AGEMA_reg_buffer_11044 ( .C (clk), .D (new_AGEMA_signal_31999), .Q (new_AGEMA_signal_32000) ) ;
    buf_clk new_AGEMA_reg_buffer_11048 ( .C (clk), .D (new_AGEMA_signal_32003), .Q (new_AGEMA_signal_32004) ) ;
    buf_clk new_AGEMA_reg_buffer_11052 ( .C (clk), .D (new_AGEMA_signal_32007), .Q (new_AGEMA_signal_32008) ) ;
    buf_clk new_AGEMA_reg_buffer_11056 ( .C (clk), .D (new_AGEMA_signal_32011), .Q (new_AGEMA_signal_32012) ) ;
    buf_clk new_AGEMA_reg_buffer_11060 ( .C (clk), .D (new_AGEMA_signal_32015), .Q (new_AGEMA_signal_32016) ) ;
    buf_clk new_AGEMA_reg_buffer_11064 ( .C (clk), .D (new_AGEMA_signal_32019), .Q (new_AGEMA_signal_32020) ) ;
    buf_clk new_AGEMA_reg_buffer_11068 ( .C (clk), .D (new_AGEMA_signal_32023), .Q (new_AGEMA_signal_32024) ) ;
    buf_clk new_AGEMA_reg_buffer_11072 ( .C (clk), .D (new_AGEMA_signal_32027), .Q (new_AGEMA_signal_32028) ) ;
    buf_clk new_AGEMA_reg_buffer_11076 ( .C (clk), .D (new_AGEMA_signal_32031), .Q (new_AGEMA_signal_32032) ) ;
    buf_clk new_AGEMA_reg_buffer_11080 ( .C (clk), .D (new_AGEMA_signal_32035), .Q (new_AGEMA_signal_32036) ) ;
    buf_clk new_AGEMA_reg_buffer_11084 ( .C (clk), .D (new_AGEMA_signal_32039), .Q (new_AGEMA_signal_32040) ) ;
    buf_clk new_AGEMA_reg_buffer_11088 ( .C (clk), .D (new_AGEMA_signal_32043), .Q (new_AGEMA_signal_32044) ) ;
    buf_clk new_AGEMA_reg_buffer_11092 ( .C (clk), .D (new_AGEMA_signal_32047), .Q (new_AGEMA_signal_32048) ) ;
    buf_clk new_AGEMA_reg_buffer_11096 ( .C (clk), .D (new_AGEMA_signal_32051), .Q (new_AGEMA_signal_32052) ) ;
    buf_clk new_AGEMA_reg_buffer_11100 ( .C (clk), .D (new_AGEMA_signal_32055), .Q (new_AGEMA_signal_32056) ) ;
    buf_clk new_AGEMA_reg_buffer_11104 ( .C (clk), .D (new_AGEMA_signal_32059), .Q (new_AGEMA_signal_32060) ) ;
    buf_clk new_AGEMA_reg_buffer_11108 ( .C (clk), .D (new_AGEMA_signal_32063), .Q (new_AGEMA_signal_32064) ) ;
    buf_clk new_AGEMA_reg_buffer_11112 ( .C (clk), .D (new_AGEMA_signal_32067), .Q (new_AGEMA_signal_32068) ) ;
    buf_clk new_AGEMA_reg_buffer_11116 ( .C (clk), .D (new_AGEMA_signal_32071), .Q (new_AGEMA_signal_32072) ) ;
    buf_clk new_AGEMA_reg_buffer_11120 ( .C (clk), .D (new_AGEMA_signal_32075), .Q (new_AGEMA_signal_32076) ) ;
    buf_clk new_AGEMA_reg_buffer_11124 ( .C (clk), .D (new_AGEMA_signal_32079), .Q (new_AGEMA_signal_32080) ) ;
    buf_clk new_AGEMA_reg_buffer_11128 ( .C (clk), .D (new_AGEMA_signal_32083), .Q (new_AGEMA_signal_32084) ) ;
    buf_clk new_AGEMA_reg_buffer_11132 ( .C (clk), .D (new_AGEMA_signal_32087), .Q (new_AGEMA_signal_32088) ) ;
    buf_clk new_AGEMA_reg_buffer_11136 ( .C (clk), .D (new_AGEMA_signal_32091), .Q (new_AGEMA_signal_32092) ) ;
    buf_clk new_AGEMA_reg_buffer_11140 ( .C (clk), .D (new_AGEMA_signal_32095), .Q (new_AGEMA_signal_32096) ) ;
    buf_clk new_AGEMA_reg_buffer_11144 ( .C (clk), .D (new_AGEMA_signal_32099), .Q (new_AGEMA_signal_32100) ) ;
    buf_clk new_AGEMA_reg_buffer_11148 ( .C (clk), .D (new_AGEMA_signal_32103), .Q (new_AGEMA_signal_32104) ) ;
    buf_clk new_AGEMA_reg_buffer_11152 ( .C (clk), .D (new_AGEMA_signal_32107), .Q (new_AGEMA_signal_32108) ) ;
    buf_clk new_AGEMA_reg_buffer_11156 ( .C (clk), .D (new_AGEMA_signal_32111), .Q (new_AGEMA_signal_32112) ) ;
    buf_clk new_AGEMA_reg_buffer_11160 ( .C (clk), .D (new_AGEMA_signal_32115), .Q (new_AGEMA_signal_32116) ) ;
    buf_clk new_AGEMA_reg_buffer_11164 ( .C (clk), .D (new_AGEMA_signal_32119), .Q (new_AGEMA_signal_32120) ) ;
    buf_clk new_AGEMA_reg_buffer_11168 ( .C (clk), .D (new_AGEMA_signal_32123), .Q (new_AGEMA_signal_32124) ) ;
    buf_clk new_AGEMA_reg_buffer_11172 ( .C (clk), .D (new_AGEMA_signal_32127), .Q (new_AGEMA_signal_32128) ) ;
    buf_clk new_AGEMA_reg_buffer_11176 ( .C (clk), .D (new_AGEMA_signal_32131), .Q (new_AGEMA_signal_32132) ) ;
    buf_clk new_AGEMA_reg_buffer_11180 ( .C (clk), .D (new_AGEMA_signal_32135), .Q (new_AGEMA_signal_32136) ) ;
    buf_clk new_AGEMA_reg_buffer_11184 ( .C (clk), .D (new_AGEMA_signal_32139), .Q (new_AGEMA_signal_32140) ) ;
    buf_clk new_AGEMA_reg_buffer_11188 ( .C (clk), .D (new_AGEMA_signal_32143), .Q (new_AGEMA_signal_32144) ) ;
    buf_clk new_AGEMA_reg_buffer_11192 ( .C (clk), .D (new_AGEMA_signal_32147), .Q (new_AGEMA_signal_32148) ) ;
    buf_clk new_AGEMA_reg_buffer_11196 ( .C (clk), .D (new_AGEMA_signal_32151), .Q (new_AGEMA_signal_32152) ) ;
    buf_clk new_AGEMA_reg_buffer_11200 ( .C (clk), .D (new_AGEMA_signal_32155), .Q (new_AGEMA_signal_32156) ) ;
    buf_clk new_AGEMA_reg_buffer_11204 ( .C (clk), .D (new_AGEMA_signal_32159), .Q (new_AGEMA_signal_32160) ) ;
    buf_clk new_AGEMA_reg_buffer_11208 ( .C (clk), .D (new_AGEMA_signal_32163), .Q (new_AGEMA_signal_32164) ) ;
    buf_clk new_AGEMA_reg_buffer_11212 ( .C (clk), .D (new_AGEMA_signal_32167), .Q (new_AGEMA_signal_32168) ) ;
    buf_clk new_AGEMA_reg_buffer_11216 ( .C (clk), .D (new_AGEMA_signal_32171), .Q (new_AGEMA_signal_32172) ) ;
    buf_clk new_AGEMA_reg_buffer_11220 ( .C (clk), .D (new_AGEMA_signal_32175), .Q (new_AGEMA_signal_32176) ) ;
    buf_clk new_AGEMA_reg_buffer_11224 ( .C (clk), .D (new_AGEMA_signal_32179), .Q (new_AGEMA_signal_32180) ) ;
    buf_clk new_AGEMA_reg_buffer_11228 ( .C (clk), .D (new_AGEMA_signal_32183), .Q (new_AGEMA_signal_32184) ) ;
    buf_clk new_AGEMA_reg_buffer_11232 ( .C (clk), .D (new_AGEMA_signal_32187), .Q (new_AGEMA_signal_32188) ) ;
    buf_clk new_AGEMA_reg_buffer_11236 ( .C (clk), .D (new_AGEMA_signal_32191), .Q (new_AGEMA_signal_32192) ) ;
    buf_clk new_AGEMA_reg_buffer_11240 ( .C (clk), .D (new_AGEMA_signal_32195), .Q (new_AGEMA_signal_32196) ) ;
    buf_clk new_AGEMA_reg_buffer_11244 ( .C (clk), .D (new_AGEMA_signal_32199), .Q (new_AGEMA_signal_32200) ) ;
    buf_clk new_AGEMA_reg_buffer_11248 ( .C (clk), .D (new_AGEMA_signal_32203), .Q (new_AGEMA_signal_32204) ) ;
    buf_clk new_AGEMA_reg_buffer_11252 ( .C (clk), .D (new_AGEMA_signal_32207), .Q (new_AGEMA_signal_32208) ) ;
    buf_clk new_AGEMA_reg_buffer_11256 ( .C (clk), .D (new_AGEMA_signal_32211), .Q (new_AGEMA_signal_32212) ) ;
    buf_clk new_AGEMA_reg_buffer_11260 ( .C (clk), .D (new_AGEMA_signal_32215), .Q (new_AGEMA_signal_32216) ) ;
    buf_clk new_AGEMA_reg_buffer_11264 ( .C (clk), .D (new_AGEMA_signal_32219), .Q (new_AGEMA_signal_32220) ) ;
    buf_clk new_AGEMA_reg_buffer_11268 ( .C (clk), .D (new_AGEMA_signal_32223), .Q (new_AGEMA_signal_32224) ) ;
    buf_clk new_AGEMA_reg_buffer_11272 ( .C (clk), .D (new_AGEMA_signal_32227), .Q (new_AGEMA_signal_32228) ) ;
    buf_clk new_AGEMA_reg_buffer_11276 ( .C (clk), .D (new_AGEMA_signal_32231), .Q (new_AGEMA_signal_32232) ) ;
    buf_clk new_AGEMA_reg_buffer_11280 ( .C (clk), .D (new_AGEMA_signal_32235), .Q (new_AGEMA_signal_32236) ) ;
    buf_clk new_AGEMA_reg_buffer_11284 ( .C (clk), .D (new_AGEMA_signal_32239), .Q (new_AGEMA_signal_32240) ) ;
    buf_clk new_AGEMA_reg_buffer_11288 ( .C (clk), .D (new_AGEMA_signal_32243), .Q (new_AGEMA_signal_32244) ) ;
    buf_clk new_AGEMA_reg_buffer_11292 ( .C (clk), .D (new_AGEMA_signal_32247), .Q (new_AGEMA_signal_32248) ) ;
    buf_clk new_AGEMA_reg_buffer_11296 ( .C (clk), .D (new_AGEMA_signal_32251), .Q (new_AGEMA_signal_32252) ) ;
    buf_clk new_AGEMA_reg_buffer_11300 ( .C (clk), .D (new_AGEMA_signal_32255), .Q (new_AGEMA_signal_32256) ) ;
    buf_clk new_AGEMA_reg_buffer_11304 ( .C (clk), .D (new_AGEMA_signal_32259), .Q (new_AGEMA_signal_32260) ) ;
    buf_clk new_AGEMA_reg_buffer_11308 ( .C (clk), .D (new_AGEMA_signal_32263), .Q (new_AGEMA_signal_32264) ) ;
    buf_clk new_AGEMA_reg_buffer_11312 ( .C (clk), .D (new_AGEMA_signal_32267), .Q (new_AGEMA_signal_32268) ) ;
    buf_clk new_AGEMA_reg_buffer_11316 ( .C (clk), .D (new_AGEMA_signal_32271), .Q (new_AGEMA_signal_32272) ) ;
    buf_clk new_AGEMA_reg_buffer_11320 ( .C (clk), .D (new_AGEMA_signal_32275), .Q (new_AGEMA_signal_32276) ) ;
    buf_clk new_AGEMA_reg_buffer_11324 ( .C (clk), .D (new_AGEMA_signal_32279), .Q (new_AGEMA_signal_32280) ) ;
    buf_clk new_AGEMA_reg_buffer_11328 ( .C (clk), .D (new_AGEMA_signal_32283), .Q (new_AGEMA_signal_32284) ) ;
    buf_clk new_AGEMA_reg_buffer_11332 ( .C (clk), .D (new_AGEMA_signal_32287), .Q (new_AGEMA_signal_32288) ) ;
    buf_clk new_AGEMA_reg_buffer_11336 ( .C (clk), .D (new_AGEMA_signal_32291), .Q (new_AGEMA_signal_32292) ) ;
    buf_clk new_AGEMA_reg_buffer_11340 ( .C (clk), .D (new_AGEMA_signal_32295), .Q (new_AGEMA_signal_32296) ) ;
    buf_clk new_AGEMA_reg_buffer_11344 ( .C (clk), .D (new_AGEMA_signal_32299), .Q (new_AGEMA_signal_32300) ) ;
    buf_clk new_AGEMA_reg_buffer_11348 ( .C (clk), .D (new_AGEMA_signal_32303), .Q (new_AGEMA_signal_32304) ) ;
    buf_clk new_AGEMA_reg_buffer_11352 ( .C (clk), .D (new_AGEMA_signal_32307), .Q (new_AGEMA_signal_32308) ) ;
    buf_clk new_AGEMA_reg_buffer_11356 ( .C (clk), .D (new_AGEMA_signal_32311), .Q (new_AGEMA_signal_32312) ) ;
    buf_clk new_AGEMA_reg_buffer_11360 ( .C (clk), .D (new_AGEMA_signal_32315), .Q (new_AGEMA_signal_32316) ) ;
    buf_clk new_AGEMA_reg_buffer_11364 ( .C (clk), .D (new_AGEMA_signal_32319), .Q (new_AGEMA_signal_32320) ) ;
    buf_clk new_AGEMA_reg_buffer_11368 ( .C (clk), .D (new_AGEMA_signal_32323), .Q (new_AGEMA_signal_32324) ) ;
    buf_clk new_AGEMA_reg_buffer_11372 ( .C (clk), .D (new_AGEMA_signal_32327), .Q (new_AGEMA_signal_32328) ) ;
    buf_clk new_AGEMA_reg_buffer_11376 ( .C (clk), .D (new_AGEMA_signal_32331), .Q (new_AGEMA_signal_32332) ) ;
    buf_clk new_AGEMA_reg_buffer_11380 ( .C (clk), .D (new_AGEMA_signal_32335), .Q (new_AGEMA_signal_32336) ) ;
    buf_clk new_AGEMA_reg_buffer_11384 ( .C (clk), .D (new_AGEMA_signal_32339), .Q (new_AGEMA_signal_32340) ) ;
    buf_clk new_AGEMA_reg_buffer_11388 ( .C (clk), .D (new_AGEMA_signal_32343), .Q (new_AGEMA_signal_32344) ) ;
    buf_clk new_AGEMA_reg_buffer_11392 ( .C (clk), .D (new_AGEMA_signal_32347), .Q (new_AGEMA_signal_32348) ) ;
    buf_clk new_AGEMA_reg_buffer_11396 ( .C (clk), .D (new_AGEMA_signal_32351), .Q (new_AGEMA_signal_32352) ) ;
    buf_clk new_AGEMA_reg_buffer_11400 ( .C (clk), .D (new_AGEMA_signal_32355), .Q (new_AGEMA_signal_32356) ) ;
    buf_clk new_AGEMA_reg_buffer_11404 ( .C (clk), .D (new_AGEMA_signal_32359), .Q (new_AGEMA_signal_32360) ) ;
    buf_clk new_AGEMA_reg_buffer_11408 ( .C (clk), .D (new_AGEMA_signal_32363), .Q (new_AGEMA_signal_32364) ) ;
    buf_clk new_AGEMA_reg_buffer_11412 ( .C (clk), .D (new_AGEMA_signal_32367), .Q (new_AGEMA_signal_32368) ) ;
    buf_clk new_AGEMA_reg_buffer_11416 ( .C (clk), .D (new_AGEMA_signal_32371), .Q (new_AGEMA_signal_32372) ) ;
    buf_clk new_AGEMA_reg_buffer_11420 ( .C (clk), .D (new_AGEMA_signal_32375), .Q (new_AGEMA_signal_32376) ) ;
    buf_clk new_AGEMA_reg_buffer_11424 ( .C (clk), .D (new_AGEMA_signal_32379), .Q (new_AGEMA_signal_32380) ) ;
    buf_clk new_AGEMA_reg_buffer_11428 ( .C (clk), .D (new_AGEMA_signal_32383), .Q (new_AGEMA_signal_32384) ) ;
    buf_clk new_AGEMA_reg_buffer_11432 ( .C (clk), .D (new_AGEMA_signal_32387), .Q (new_AGEMA_signal_32388) ) ;
    buf_clk new_AGEMA_reg_buffer_11436 ( .C (clk), .D (new_AGEMA_signal_32391), .Q (new_AGEMA_signal_32392) ) ;
    buf_clk new_AGEMA_reg_buffer_11440 ( .C (clk), .D (new_AGEMA_signal_32395), .Q (new_AGEMA_signal_32396) ) ;
    buf_clk new_AGEMA_reg_buffer_11444 ( .C (clk), .D (new_AGEMA_signal_32399), .Q (new_AGEMA_signal_32400) ) ;
    buf_clk new_AGEMA_reg_buffer_11448 ( .C (clk), .D (new_AGEMA_signal_32403), .Q (new_AGEMA_signal_32404) ) ;
    buf_clk new_AGEMA_reg_buffer_11452 ( .C (clk), .D (new_AGEMA_signal_32407), .Q (new_AGEMA_signal_32408) ) ;
    buf_clk new_AGEMA_reg_buffer_11456 ( .C (clk), .D (new_AGEMA_signal_32411), .Q (new_AGEMA_signal_32412) ) ;
    buf_clk new_AGEMA_reg_buffer_11460 ( .C (clk), .D (new_AGEMA_signal_32415), .Q (new_AGEMA_signal_32416) ) ;
    buf_clk new_AGEMA_reg_buffer_11464 ( .C (clk), .D (new_AGEMA_signal_32419), .Q (new_AGEMA_signal_32420) ) ;
    buf_clk new_AGEMA_reg_buffer_11468 ( .C (clk), .D (new_AGEMA_signal_32423), .Q (new_AGEMA_signal_32424) ) ;
    buf_clk new_AGEMA_reg_buffer_11472 ( .C (clk), .D (new_AGEMA_signal_32427), .Q (new_AGEMA_signal_32428) ) ;
    buf_clk new_AGEMA_reg_buffer_11476 ( .C (clk), .D (new_AGEMA_signal_32431), .Q (new_AGEMA_signal_32432) ) ;
    buf_clk new_AGEMA_reg_buffer_11480 ( .C (clk), .D (new_AGEMA_signal_32435), .Q (new_AGEMA_signal_32436) ) ;
    buf_clk new_AGEMA_reg_buffer_11484 ( .C (clk), .D (new_AGEMA_signal_32439), .Q (new_AGEMA_signal_32440) ) ;
    buf_clk new_AGEMA_reg_buffer_11488 ( .C (clk), .D (new_AGEMA_signal_32443), .Q (new_AGEMA_signal_32444) ) ;
    buf_clk new_AGEMA_reg_buffer_11492 ( .C (clk), .D (new_AGEMA_signal_32447), .Q (new_AGEMA_signal_32448) ) ;
    buf_clk new_AGEMA_reg_buffer_11496 ( .C (clk), .D (new_AGEMA_signal_32451), .Q (new_AGEMA_signal_32452) ) ;
    buf_clk new_AGEMA_reg_buffer_11500 ( .C (clk), .D (new_AGEMA_signal_32455), .Q (new_AGEMA_signal_32456) ) ;
    buf_clk new_AGEMA_reg_buffer_11504 ( .C (clk), .D (new_AGEMA_signal_32459), .Q (new_AGEMA_signal_32460) ) ;
    buf_clk new_AGEMA_reg_buffer_11508 ( .C (clk), .D (new_AGEMA_signal_32463), .Q (new_AGEMA_signal_32464) ) ;
    buf_clk new_AGEMA_reg_buffer_11512 ( .C (clk), .D (new_AGEMA_signal_32467), .Q (new_AGEMA_signal_32468) ) ;
    buf_clk new_AGEMA_reg_buffer_11516 ( .C (clk), .D (new_AGEMA_signal_32471), .Q (new_AGEMA_signal_32472) ) ;
    buf_clk new_AGEMA_reg_buffer_11520 ( .C (clk), .D (new_AGEMA_signal_32475), .Q (new_AGEMA_signal_32476) ) ;
    buf_clk new_AGEMA_reg_buffer_11524 ( .C (clk), .D (new_AGEMA_signal_32479), .Q (new_AGEMA_signal_32480) ) ;
    buf_clk new_AGEMA_reg_buffer_11528 ( .C (clk), .D (new_AGEMA_signal_32483), .Q (new_AGEMA_signal_32484) ) ;
    buf_clk new_AGEMA_reg_buffer_11532 ( .C (clk), .D (new_AGEMA_signal_32487), .Q (new_AGEMA_signal_32488) ) ;
    buf_clk new_AGEMA_reg_buffer_11536 ( .C (clk), .D (new_AGEMA_signal_32491), .Q (new_AGEMA_signal_32492) ) ;
    buf_clk new_AGEMA_reg_buffer_11540 ( .C (clk), .D (new_AGEMA_signal_32495), .Q (new_AGEMA_signal_32496) ) ;
    buf_clk new_AGEMA_reg_buffer_11544 ( .C (clk), .D (new_AGEMA_signal_32499), .Q (new_AGEMA_signal_32500) ) ;
    buf_clk new_AGEMA_reg_buffer_11548 ( .C (clk), .D (new_AGEMA_signal_32503), .Q (new_AGEMA_signal_32504) ) ;
    buf_clk new_AGEMA_reg_buffer_11552 ( .C (clk), .D (new_AGEMA_signal_32507), .Q (new_AGEMA_signal_32508) ) ;
    buf_clk new_AGEMA_reg_buffer_11556 ( .C (clk), .D (new_AGEMA_signal_32511), .Q (new_AGEMA_signal_32512) ) ;
    buf_clk new_AGEMA_reg_buffer_11560 ( .C (clk), .D (new_AGEMA_signal_32515), .Q (new_AGEMA_signal_32516) ) ;
    buf_clk new_AGEMA_reg_buffer_11564 ( .C (clk), .D (new_AGEMA_signal_32519), .Q (new_AGEMA_signal_32520) ) ;
    buf_clk new_AGEMA_reg_buffer_11568 ( .C (clk), .D (new_AGEMA_signal_32523), .Q (new_AGEMA_signal_32524) ) ;
    buf_clk new_AGEMA_reg_buffer_11572 ( .C (clk), .D (new_AGEMA_signal_32527), .Q (new_AGEMA_signal_32528) ) ;
    buf_clk new_AGEMA_reg_buffer_11576 ( .C (clk), .D (new_AGEMA_signal_32531), .Q (new_AGEMA_signal_32532) ) ;
    buf_clk new_AGEMA_reg_buffer_11580 ( .C (clk), .D (new_AGEMA_signal_32535), .Q (new_AGEMA_signal_32536) ) ;
    buf_clk new_AGEMA_reg_buffer_11584 ( .C (clk), .D (new_AGEMA_signal_32539), .Q (new_AGEMA_signal_32540) ) ;
    buf_clk new_AGEMA_reg_buffer_11588 ( .C (clk), .D (new_AGEMA_signal_32543), .Q (new_AGEMA_signal_32544) ) ;
    buf_clk new_AGEMA_reg_buffer_11592 ( .C (clk), .D (new_AGEMA_signal_32547), .Q (new_AGEMA_signal_32548) ) ;
    buf_clk new_AGEMA_reg_buffer_11596 ( .C (clk), .D (new_AGEMA_signal_32551), .Q (new_AGEMA_signal_32552) ) ;
    buf_clk new_AGEMA_reg_buffer_11600 ( .C (clk), .D (new_AGEMA_signal_32555), .Q (new_AGEMA_signal_32556) ) ;
    buf_clk new_AGEMA_reg_buffer_11604 ( .C (clk), .D (new_AGEMA_signal_32559), .Q (new_AGEMA_signal_32560) ) ;
    buf_clk new_AGEMA_reg_buffer_11608 ( .C (clk), .D (new_AGEMA_signal_32563), .Q (new_AGEMA_signal_32564) ) ;
    buf_clk new_AGEMA_reg_buffer_11612 ( .C (clk), .D (new_AGEMA_signal_32567), .Q (new_AGEMA_signal_32568) ) ;
    buf_clk new_AGEMA_reg_buffer_11616 ( .C (clk), .D (new_AGEMA_signal_32571), .Q (new_AGEMA_signal_32572) ) ;
    buf_clk new_AGEMA_reg_buffer_11620 ( .C (clk), .D (new_AGEMA_signal_32575), .Q (new_AGEMA_signal_32576) ) ;
    buf_clk new_AGEMA_reg_buffer_11624 ( .C (clk), .D (new_AGEMA_signal_32579), .Q (new_AGEMA_signal_32580) ) ;
    buf_clk new_AGEMA_reg_buffer_11628 ( .C (clk), .D (new_AGEMA_signal_32583), .Q (new_AGEMA_signal_32584) ) ;
    buf_clk new_AGEMA_reg_buffer_11632 ( .C (clk), .D (new_AGEMA_signal_32587), .Q (new_AGEMA_signal_32588) ) ;
    buf_clk new_AGEMA_reg_buffer_11636 ( .C (clk), .D (new_AGEMA_signal_32591), .Q (new_AGEMA_signal_32592) ) ;
    buf_clk new_AGEMA_reg_buffer_11640 ( .C (clk), .D (new_AGEMA_signal_32595), .Q (new_AGEMA_signal_32596) ) ;
    buf_clk new_AGEMA_reg_buffer_11644 ( .C (clk), .D (new_AGEMA_signal_32599), .Q (new_AGEMA_signal_32600) ) ;
    buf_clk new_AGEMA_reg_buffer_11648 ( .C (clk), .D (new_AGEMA_signal_32603), .Q (new_AGEMA_signal_32604) ) ;
    buf_clk new_AGEMA_reg_buffer_11652 ( .C (clk), .D (new_AGEMA_signal_32607), .Q (new_AGEMA_signal_32608) ) ;
    buf_clk new_AGEMA_reg_buffer_11656 ( .C (clk), .D (new_AGEMA_signal_32611), .Q (new_AGEMA_signal_32612) ) ;
    buf_clk new_AGEMA_reg_buffer_11660 ( .C (clk), .D (new_AGEMA_signal_32615), .Q (new_AGEMA_signal_32616) ) ;
    buf_clk new_AGEMA_reg_buffer_11664 ( .C (clk), .D (new_AGEMA_signal_32619), .Q (new_AGEMA_signal_32620) ) ;
    buf_clk new_AGEMA_reg_buffer_11668 ( .C (clk), .D (new_AGEMA_signal_32623), .Q (new_AGEMA_signal_32624) ) ;
    buf_clk new_AGEMA_reg_buffer_11672 ( .C (clk), .D (new_AGEMA_signal_32627), .Q (new_AGEMA_signal_32628) ) ;
    buf_clk new_AGEMA_reg_buffer_11676 ( .C (clk), .D (new_AGEMA_signal_32631), .Q (new_AGEMA_signal_32632) ) ;
    buf_clk new_AGEMA_reg_buffer_11680 ( .C (clk), .D (new_AGEMA_signal_32635), .Q (new_AGEMA_signal_32636) ) ;
    buf_clk new_AGEMA_reg_buffer_11684 ( .C (clk), .D (new_AGEMA_signal_32639), .Q (new_AGEMA_signal_32640) ) ;
    buf_clk new_AGEMA_reg_buffer_11688 ( .C (clk), .D (new_AGEMA_signal_32643), .Q (new_AGEMA_signal_32644) ) ;
    buf_clk new_AGEMA_reg_buffer_11692 ( .C (clk), .D (new_AGEMA_signal_32647), .Q (new_AGEMA_signal_32648) ) ;
    buf_clk new_AGEMA_reg_buffer_11696 ( .C (clk), .D (new_AGEMA_signal_32651), .Q (new_AGEMA_signal_32652) ) ;
    buf_clk new_AGEMA_reg_buffer_11700 ( .C (clk), .D (new_AGEMA_signal_32655), .Q (new_AGEMA_signal_32656) ) ;
    buf_clk new_AGEMA_reg_buffer_11704 ( .C (clk), .D (new_AGEMA_signal_32659), .Q (new_AGEMA_signal_32660) ) ;
    buf_clk new_AGEMA_reg_buffer_11708 ( .C (clk), .D (new_AGEMA_signal_32663), .Q (new_AGEMA_signal_32664) ) ;
    buf_clk new_AGEMA_reg_buffer_11712 ( .C (clk), .D (new_AGEMA_signal_32667), .Q (new_AGEMA_signal_32668) ) ;
    buf_clk new_AGEMA_reg_buffer_11716 ( .C (clk), .D (new_AGEMA_signal_32671), .Q (new_AGEMA_signal_32672) ) ;
    buf_clk new_AGEMA_reg_buffer_11720 ( .C (clk), .D (new_AGEMA_signal_32675), .Q (new_AGEMA_signal_32676) ) ;
    buf_clk new_AGEMA_reg_buffer_11724 ( .C (clk), .D (new_AGEMA_signal_32679), .Q (new_AGEMA_signal_32680) ) ;
    buf_clk new_AGEMA_reg_buffer_11728 ( .C (clk), .D (new_AGEMA_signal_32683), .Q (new_AGEMA_signal_32684) ) ;
    buf_clk new_AGEMA_reg_buffer_11732 ( .C (clk), .D (new_AGEMA_signal_32687), .Q (new_AGEMA_signal_32688) ) ;
    buf_clk new_AGEMA_reg_buffer_11736 ( .C (clk), .D (new_AGEMA_signal_32691), .Q (new_AGEMA_signal_32692) ) ;
    buf_clk new_AGEMA_reg_buffer_11740 ( .C (clk), .D (new_AGEMA_signal_32695), .Q (new_AGEMA_signal_32696) ) ;
    buf_clk new_AGEMA_reg_buffer_11744 ( .C (clk), .D (new_AGEMA_signal_32699), .Q (new_AGEMA_signal_32700) ) ;
    buf_clk new_AGEMA_reg_buffer_11748 ( .C (clk), .D (new_AGEMA_signal_32703), .Q (new_AGEMA_signal_32704) ) ;
    buf_clk new_AGEMA_reg_buffer_11752 ( .C (clk), .D (new_AGEMA_signal_32707), .Q (new_AGEMA_signal_32708) ) ;
    buf_clk new_AGEMA_reg_buffer_11756 ( .C (clk), .D (new_AGEMA_signal_32711), .Q (new_AGEMA_signal_32712) ) ;
    buf_clk new_AGEMA_reg_buffer_11760 ( .C (clk), .D (new_AGEMA_signal_32715), .Q (new_AGEMA_signal_32716) ) ;
    buf_clk new_AGEMA_reg_buffer_11764 ( .C (clk), .D (new_AGEMA_signal_32719), .Q (new_AGEMA_signal_32720) ) ;
    buf_clk new_AGEMA_reg_buffer_11768 ( .C (clk), .D (new_AGEMA_signal_32723), .Q (new_AGEMA_signal_32724) ) ;
    buf_clk new_AGEMA_reg_buffer_11772 ( .C (clk), .D (new_AGEMA_signal_32727), .Q (new_AGEMA_signal_32728) ) ;
    buf_clk new_AGEMA_reg_buffer_11776 ( .C (clk), .D (new_AGEMA_signal_32731), .Q (new_AGEMA_signal_32732) ) ;
    buf_clk new_AGEMA_reg_buffer_11780 ( .C (clk), .D (new_AGEMA_signal_32735), .Q (new_AGEMA_signal_32736) ) ;
    buf_clk new_AGEMA_reg_buffer_11784 ( .C (clk), .D (new_AGEMA_signal_32739), .Q (new_AGEMA_signal_32740) ) ;
    buf_clk new_AGEMA_reg_buffer_11788 ( .C (clk), .D (new_AGEMA_signal_32743), .Q (new_AGEMA_signal_32744) ) ;
    buf_clk new_AGEMA_reg_buffer_11792 ( .C (clk), .D (new_AGEMA_signal_32747), .Q (new_AGEMA_signal_32748) ) ;
    buf_clk new_AGEMA_reg_buffer_11796 ( .C (clk), .D (new_AGEMA_signal_32751), .Q (new_AGEMA_signal_32752) ) ;
    buf_clk new_AGEMA_reg_buffer_11800 ( .C (clk), .D (new_AGEMA_signal_32755), .Q (new_AGEMA_signal_32756) ) ;
    buf_clk new_AGEMA_reg_buffer_11804 ( .C (clk), .D (new_AGEMA_signal_32759), .Q (new_AGEMA_signal_32760) ) ;
    buf_clk new_AGEMA_reg_buffer_11808 ( .C (clk), .D (new_AGEMA_signal_32763), .Q (new_AGEMA_signal_32764) ) ;
    buf_clk new_AGEMA_reg_buffer_11812 ( .C (clk), .D (new_AGEMA_signal_32767), .Q (new_AGEMA_signal_32768) ) ;
    buf_clk new_AGEMA_reg_buffer_11816 ( .C (clk), .D (new_AGEMA_signal_32771), .Q (new_AGEMA_signal_32772) ) ;
    buf_clk new_AGEMA_reg_buffer_11820 ( .C (clk), .D (new_AGEMA_signal_32775), .Q (new_AGEMA_signal_32776) ) ;
    buf_clk new_AGEMA_reg_buffer_11824 ( .C (clk), .D (new_AGEMA_signal_32779), .Q (new_AGEMA_signal_32780) ) ;
    buf_clk new_AGEMA_reg_buffer_11828 ( .C (clk), .D (new_AGEMA_signal_32783), .Q (new_AGEMA_signal_32784) ) ;
    buf_clk new_AGEMA_reg_buffer_11832 ( .C (clk), .D (new_AGEMA_signal_32787), .Q (new_AGEMA_signal_32788) ) ;
    buf_clk new_AGEMA_reg_buffer_11836 ( .C (clk), .D (new_AGEMA_signal_32791), .Q (new_AGEMA_signal_32792) ) ;
    buf_clk new_AGEMA_reg_buffer_11840 ( .C (clk), .D (new_AGEMA_signal_32795), .Q (new_AGEMA_signal_32796) ) ;
    buf_clk new_AGEMA_reg_buffer_11844 ( .C (clk), .D (new_AGEMA_signal_32799), .Q (new_AGEMA_signal_32800) ) ;
    buf_clk new_AGEMA_reg_buffer_11848 ( .C (clk), .D (new_AGEMA_signal_32803), .Q (new_AGEMA_signal_32804) ) ;
    buf_clk new_AGEMA_reg_buffer_11852 ( .C (clk), .D (new_AGEMA_signal_32807), .Q (new_AGEMA_signal_32808) ) ;
    buf_clk new_AGEMA_reg_buffer_11856 ( .C (clk), .D (new_AGEMA_signal_32811), .Q (new_AGEMA_signal_32812) ) ;
    buf_clk new_AGEMA_reg_buffer_11860 ( .C (clk), .D (new_AGEMA_signal_32815), .Q (new_AGEMA_signal_32816) ) ;
    buf_clk new_AGEMA_reg_buffer_11864 ( .C (clk), .D (new_AGEMA_signal_32819), .Q (new_AGEMA_signal_32820) ) ;
    buf_clk new_AGEMA_reg_buffer_11868 ( .C (clk), .D (new_AGEMA_signal_32823), .Q (new_AGEMA_signal_32824) ) ;
    buf_clk new_AGEMA_reg_buffer_11872 ( .C (clk), .D (new_AGEMA_signal_32827), .Q (new_AGEMA_signal_32828) ) ;
    buf_clk new_AGEMA_reg_buffer_11876 ( .C (clk), .D (new_AGEMA_signal_32831), .Q (new_AGEMA_signal_32832) ) ;
    buf_clk new_AGEMA_reg_buffer_11880 ( .C (clk), .D (new_AGEMA_signal_32835), .Q (new_AGEMA_signal_32836) ) ;
    buf_clk new_AGEMA_reg_buffer_11884 ( .C (clk), .D (new_AGEMA_signal_32839), .Q (new_AGEMA_signal_32840) ) ;
    buf_clk new_AGEMA_reg_buffer_11888 ( .C (clk), .D (new_AGEMA_signal_32843), .Q (new_AGEMA_signal_32844) ) ;
    buf_clk new_AGEMA_reg_buffer_11892 ( .C (clk), .D (new_AGEMA_signal_32847), .Q (new_AGEMA_signal_32848) ) ;
    buf_clk new_AGEMA_reg_buffer_11896 ( .C (clk), .D (new_AGEMA_signal_32851), .Q (new_AGEMA_signal_32852) ) ;
    buf_clk new_AGEMA_reg_buffer_11900 ( .C (clk), .D (new_AGEMA_signal_32855), .Q (new_AGEMA_signal_32856) ) ;
    buf_clk new_AGEMA_reg_buffer_11904 ( .C (clk), .D (new_AGEMA_signal_32859), .Q (new_AGEMA_signal_32860) ) ;
    buf_clk new_AGEMA_reg_buffer_11908 ( .C (clk), .D (new_AGEMA_signal_32863), .Q (new_AGEMA_signal_32864) ) ;
    buf_clk new_AGEMA_reg_buffer_11912 ( .C (clk), .D (new_AGEMA_signal_32867), .Q (new_AGEMA_signal_32868) ) ;
    buf_clk new_AGEMA_reg_buffer_11916 ( .C (clk), .D (new_AGEMA_signal_32871), .Q (new_AGEMA_signal_32872) ) ;
    buf_clk new_AGEMA_reg_buffer_11920 ( .C (clk), .D (new_AGEMA_signal_32875), .Q (new_AGEMA_signal_32876) ) ;
    buf_clk new_AGEMA_reg_buffer_11924 ( .C (clk), .D (new_AGEMA_signal_32879), .Q (new_AGEMA_signal_32880) ) ;
    buf_clk new_AGEMA_reg_buffer_11928 ( .C (clk), .D (new_AGEMA_signal_32883), .Q (new_AGEMA_signal_32884) ) ;
    buf_clk new_AGEMA_reg_buffer_11932 ( .C (clk), .D (new_AGEMA_signal_32887), .Q (new_AGEMA_signal_32888) ) ;
    buf_clk new_AGEMA_reg_buffer_11936 ( .C (clk), .D (new_AGEMA_signal_32891), .Q (new_AGEMA_signal_32892) ) ;
    buf_clk new_AGEMA_reg_buffer_11940 ( .C (clk), .D (new_AGEMA_signal_32895), .Q (new_AGEMA_signal_32896) ) ;
    buf_clk new_AGEMA_reg_buffer_11944 ( .C (clk), .D (new_AGEMA_signal_32899), .Q (new_AGEMA_signal_32900) ) ;
    buf_clk new_AGEMA_reg_buffer_11948 ( .C (clk), .D (new_AGEMA_signal_32903), .Q (new_AGEMA_signal_32904) ) ;
    buf_clk new_AGEMA_reg_buffer_11952 ( .C (clk), .D (new_AGEMA_signal_32907), .Q (new_AGEMA_signal_32908) ) ;
    buf_clk new_AGEMA_reg_buffer_11956 ( .C (clk), .D (new_AGEMA_signal_32911), .Q (new_AGEMA_signal_32912) ) ;
    buf_clk new_AGEMA_reg_buffer_11960 ( .C (clk), .D (new_AGEMA_signal_32915), .Q (new_AGEMA_signal_32916) ) ;
    buf_clk new_AGEMA_reg_buffer_11964 ( .C (clk), .D (new_AGEMA_signal_32919), .Q (new_AGEMA_signal_32920) ) ;
    buf_clk new_AGEMA_reg_buffer_11968 ( .C (clk), .D (new_AGEMA_signal_32923), .Q (new_AGEMA_signal_32924) ) ;
    buf_clk new_AGEMA_reg_buffer_11972 ( .C (clk), .D (new_AGEMA_signal_32927), .Q (new_AGEMA_signal_32928) ) ;
    buf_clk new_AGEMA_reg_buffer_11976 ( .C (clk), .D (new_AGEMA_signal_32931), .Q (new_AGEMA_signal_32932) ) ;
    buf_clk new_AGEMA_reg_buffer_11980 ( .C (clk), .D (new_AGEMA_signal_32935), .Q (new_AGEMA_signal_32936) ) ;
    buf_clk new_AGEMA_reg_buffer_11984 ( .C (clk), .D (new_AGEMA_signal_32939), .Q (new_AGEMA_signal_32940) ) ;
    buf_clk new_AGEMA_reg_buffer_11988 ( .C (clk), .D (new_AGEMA_signal_32943), .Q (new_AGEMA_signal_32944) ) ;
    buf_clk new_AGEMA_reg_buffer_11992 ( .C (clk), .D (new_AGEMA_signal_32947), .Q (new_AGEMA_signal_32948) ) ;
    buf_clk new_AGEMA_reg_buffer_11996 ( .C (clk), .D (new_AGEMA_signal_32951), .Q (new_AGEMA_signal_32952) ) ;
    buf_clk new_AGEMA_reg_buffer_12000 ( .C (clk), .D (new_AGEMA_signal_32955), .Q (new_AGEMA_signal_32956) ) ;
    buf_clk new_AGEMA_reg_buffer_12004 ( .C (clk), .D (new_AGEMA_signal_32959), .Q (new_AGEMA_signal_32960) ) ;
    buf_clk new_AGEMA_reg_buffer_12008 ( .C (clk), .D (new_AGEMA_signal_32963), .Q (new_AGEMA_signal_32964) ) ;
    buf_clk new_AGEMA_reg_buffer_12012 ( .C (clk), .D (new_AGEMA_signal_32967), .Q (new_AGEMA_signal_32968) ) ;
    buf_clk new_AGEMA_reg_buffer_12016 ( .C (clk), .D (new_AGEMA_signal_32971), .Q (new_AGEMA_signal_32972) ) ;
    buf_clk new_AGEMA_reg_buffer_12020 ( .C (clk), .D (new_AGEMA_signal_32975), .Q (new_AGEMA_signal_32976) ) ;
    buf_clk new_AGEMA_reg_buffer_12024 ( .C (clk), .D (new_AGEMA_signal_32979), .Q (new_AGEMA_signal_32980) ) ;
    buf_clk new_AGEMA_reg_buffer_12028 ( .C (clk), .D (new_AGEMA_signal_32983), .Q (new_AGEMA_signal_32984) ) ;
    buf_clk new_AGEMA_reg_buffer_12032 ( .C (clk), .D (new_AGEMA_signal_32987), .Q (new_AGEMA_signal_32988) ) ;
    buf_clk new_AGEMA_reg_buffer_12036 ( .C (clk), .D (new_AGEMA_signal_32991), .Q (new_AGEMA_signal_32992) ) ;
    buf_clk new_AGEMA_reg_buffer_12040 ( .C (clk), .D (new_AGEMA_signal_32995), .Q (new_AGEMA_signal_32996) ) ;
    buf_clk new_AGEMA_reg_buffer_12044 ( .C (clk), .D (new_AGEMA_signal_32999), .Q (new_AGEMA_signal_33000) ) ;
    buf_clk new_AGEMA_reg_buffer_12048 ( .C (clk), .D (new_AGEMA_signal_33003), .Q (new_AGEMA_signal_33004) ) ;
    buf_clk new_AGEMA_reg_buffer_12052 ( .C (clk), .D (new_AGEMA_signal_33007), .Q (new_AGEMA_signal_33008) ) ;
    buf_clk new_AGEMA_reg_buffer_12056 ( .C (clk), .D (new_AGEMA_signal_33011), .Q (new_AGEMA_signal_33012) ) ;
    buf_clk new_AGEMA_reg_buffer_12060 ( .C (clk), .D (new_AGEMA_signal_33015), .Q (new_AGEMA_signal_33016) ) ;
    buf_clk new_AGEMA_reg_buffer_12064 ( .C (clk), .D (new_AGEMA_signal_33019), .Q (new_AGEMA_signal_33020) ) ;
    buf_clk new_AGEMA_reg_buffer_12068 ( .C (clk), .D (new_AGEMA_signal_33023), .Q (new_AGEMA_signal_33024) ) ;
    buf_clk new_AGEMA_reg_buffer_12072 ( .C (clk), .D (new_AGEMA_signal_33027), .Q (new_AGEMA_signal_33028) ) ;
    buf_clk new_AGEMA_reg_buffer_12076 ( .C (clk), .D (new_AGEMA_signal_33031), .Q (new_AGEMA_signal_33032) ) ;
    buf_clk new_AGEMA_reg_buffer_12080 ( .C (clk), .D (new_AGEMA_signal_33035), .Q (new_AGEMA_signal_33036) ) ;
    buf_clk new_AGEMA_reg_buffer_12084 ( .C (clk), .D (new_AGEMA_signal_33039), .Q (new_AGEMA_signal_33040) ) ;
    buf_clk new_AGEMA_reg_buffer_12088 ( .C (clk), .D (new_AGEMA_signal_33043), .Q (new_AGEMA_signal_33044) ) ;
    buf_clk new_AGEMA_reg_buffer_12092 ( .C (clk), .D (new_AGEMA_signal_33047), .Q (new_AGEMA_signal_33048) ) ;
    buf_clk new_AGEMA_reg_buffer_12096 ( .C (clk), .D (new_AGEMA_signal_33051), .Q (new_AGEMA_signal_33052) ) ;
    buf_clk new_AGEMA_reg_buffer_12100 ( .C (clk), .D (new_AGEMA_signal_33055), .Q (new_AGEMA_signal_33056) ) ;
    buf_clk new_AGEMA_reg_buffer_12104 ( .C (clk), .D (new_AGEMA_signal_33059), .Q (new_AGEMA_signal_33060) ) ;
    buf_clk new_AGEMA_reg_buffer_12108 ( .C (clk), .D (new_AGEMA_signal_33063), .Q (new_AGEMA_signal_33064) ) ;
    buf_clk new_AGEMA_reg_buffer_12112 ( .C (clk), .D (new_AGEMA_signal_33067), .Q (new_AGEMA_signal_33068) ) ;
    buf_clk new_AGEMA_reg_buffer_12116 ( .C (clk), .D (new_AGEMA_signal_33071), .Q (new_AGEMA_signal_33072) ) ;
    buf_clk new_AGEMA_reg_buffer_12120 ( .C (clk), .D (new_AGEMA_signal_33075), .Q (new_AGEMA_signal_33076) ) ;
    buf_clk new_AGEMA_reg_buffer_12124 ( .C (clk), .D (new_AGEMA_signal_33079), .Q (new_AGEMA_signal_33080) ) ;
    buf_clk new_AGEMA_reg_buffer_12128 ( .C (clk), .D (new_AGEMA_signal_33083), .Q (new_AGEMA_signal_33084) ) ;
    buf_clk new_AGEMA_reg_buffer_12132 ( .C (clk), .D (new_AGEMA_signal_33087), .Q (new_AGEMA_signal_33088) ) ;
    buf_clk new_AGEMA_reg_buffer_12136 ( .C (clk), .D (new_AGEMA_signal_33091), .Q (new_AGEMA_signal_33092) ) ;
    buf_clk new_AGEMA_reg_buffer_12140 ( .C (clk), .D (new_AGEMA_signal_33095), .Q (new_AGEMA_signal_33096) ) ;
    buf_clk new_AGEMA_reg_buffer_12144 ( .C (clk), .D (new_AGEMA_signal_33099), .Q (new_AGEMA_signal_33100) ) ;
    buf_clk new_AGEMA_reg_buffer_12148 ( .C (clk), .D (new_AGEMA_signal_33103), .Q (new_AGEMA_signal_33104) ) ;
    buf_clk new_AGEMA_reg_buffer_12152 ( .C (clk), .D (new_AGEMA_signal_33107), .Q (new_AGEMA_signal_33108) ) ;
    buf_clk new_AGEMA_reg_buffer_12156 ( .C (clk), .D (new_AGEMA_signal_33111), .Q (new_AGEMA_signal_33112) ) ;
    buf_clk new_AGEMA_reg_buffer_12160 ( .C (clk), .D (new_AGEMA_signal_33115), .Q (new_AGEMA_signal_33116) ) ;
    buf_clk new_AGEMA_reg_buffer_12164 ( .C (clk), .D (new_AGEMA_signal_33119), .Q (new_AGEMA_signal_33120) ) ;
    buf_clk new_AGEMA_reg_buffer_12168 ( .C (clk), .D (new_AGEMA_signal_33123), .Q (new_AGEMA_signal_33124) ) ;
    buf_clk new_AGEMA_reg_buffer_12172 ( .C (clk), .D (new_AGEMA_signal_33127), .Q (new_AGEMA_signal_33128) ) ;
    buf_clk new_AGEMA_reg_buffer_12176 ( .C (clk), .D (new_AGEMA_signal_33131), .Q (new_AGEMA_signal_33132) ) ;
    buf_clk new_AGEMA_reg_buffer_12180 ( .C (clk), .D (new_AGEMA_signal_33135), .Q (new_AGEMA_signal_33136) ) ;
    buf_clk new_AGEMA_reg_buffer_12184 ( .C (clk), .D (new_AGEMA_signal_33139), .Q (new_AGEMA_signal_33140) ) ;
    buf_clk new_AGEMA_reg_buffer_12188 ( .C (clk), .D (new_AGEMA_signal_33143), .Q (new_AGEMA_signal_33144) ) ;
    buf_clk new_AGEMA_reg_buffer_12192 ( .C (clk), .D (new_AGEMA_signal_33147), .Q (new_AGEMA_signal_33148) ) ;
    buf_clk new_AGEMA_reg_buffer_12196 ( .C (clk), .D (new_AGEMA_signal_33151), .Q (new_AGEMA_signal_33152) ) ;
    buf_clk new_AGEMA_reg_buffer_12200 ( .C (clk), .D (new_AGEMA_signal_33155), .Q (new_AGEMA_signal_33156) ) ;
    buf_clk new_AGEMA_reg_buffer_12204 ( .C (clk), .D (new_AGEMA_signal_33159), .Q (new_AGEMA_signal_33160) ) ;
    buf_clk new_AGEMA_reg_buffer_12208 ( .C (clk), .D (new_AGEMA_signal_33163), .Q (new_AGEMA_signal_33164) ) ;
    buf_clk new_AGEMA_reg_buffer_12212 ( .C (clk), .D (new_AGEMA_signal_33167), .Q (new_AGEMA_signal_33168) ) ;
    buf_clk new_AGEMA_reg_buffer_12216 ( .C (clk), .D (new_AGEMA_signal_33171), .Q (new_AGEMA_signal_33172) ) ;
    buf_clk new_AGEMA_reg_buffer_12220 ( .C (clk), .D (new_AGEMA_signal_33175), .Q (new_AGEMA_signal_33176) ) ;
    buf_clk new_AGEMA_reg_buffer_12224 ( .C (clk), .D (new_AGEMA_signal_33179), .Q (new_AGEMA_signal_33180) ) ;
    buf_clk new_AGEMA_reg_buffer_12228 ( .C (clk), .D (new_AGEMA_signal_33183), .Q (new_AGEMA_signal_33184) ) ;
    buf_clk new_AGEMA_reg_buffer_12232 ( .C (clk), .D (new_AGEMA_signal_33187), .Q (new_AGEMA_signal_33188) ) ;
    buf_clk new_AGEMA_reg_buffer_12236 ( .C (clk), .D (new_AGEMA_signal_33191), .Q (new_AGEMA_signal_33192) ) ;
    buf_clk new_AGEMA_reg_buffer_12240 ( .C (clk), .D (new_AGEMA_signal_33195), .Q (new_AGEMA_signal_33196) ) ;
    buf_clk new_AGEMA_reg_buffer_12244 ( .C (clk), .D (new_AGEMA_signal_33199), .Q (new_AGEMA_signal_33200) ) ;
    buf_clk new_AGEMA_reg_buffer_12248 ( .C (clk), .D (new_AGEMA_signal_33203), .Q (new_AGEMA_signal_33204) ) ;
    buf_clk new_AGEMA_reg_buffer_12252 ( .C (clk), .D (new_AGEMA_signal_33207), .Q (new_AGEMA_signal_33208) ) ;
    buf_clk new_AGEMA_reg_buffer_12256 ( .C (clk), .D (new_AGEMA_signal_33211), .Q (new_AGEMA_signal_33212) ) ;
    buf_clk new_AGEMA_reg_buffer_12260 ( .C (clk), .D (new_AGEMA_signal_33215), .Q (new_AGEMA_signal_33216) ) ;
    buf_clk new_AGEMA_reg_buffer_12264 ( .C (clk), .D (new_AGEMA_signal_33219), .Q (new_AGEMA_signal_33220) ) ;
    buf_clk new_AGEMA_reg_buffer_12268 ( .C (clk), .D (new_AGEMA_signal_33223), .Q (new_AGEMA_signal_33224) ) ;
    buf_clk new_AGEMA_reg_buffer_12272 ( .C (clk), .D (new_AGEMA_signal_33227), .Q (new_AGEMA_signal_33228) ) ;
    buf_clk new_AGEMA_reg_buffer_12276 ( .C (clk), .D (new_AGEMA_signal_33231), .Q (new_AGEMA_signal_33232) ) ;
    buf_clk new_AGEMA_reg_buffer_12280 ( .C (clk), .D (new_AGEMA_signal_33235), .Q (new_AGEMA_signal_33236) ) ;
    buf_clk new_AGEMA_reg_buffer_12284 ( .C (clk), .D (new_AGEMA_signal_33239), .Q (new_AGEMA_signal_33240) ) ;
    buf_clk new_AGEMA_reg_buffer_12288 ( .C (clk), .D (new_AGEMA_signal_33243), .Q (new_AGEMA_signal_33244) ) ;
    buf_clk new_AGEMA_reg_buffer_12292 ( .C (clk), .D (new_AGEMA_signal_33247), .Q (new_AGEMA_signal_33248) ) ;
    buf_clk new_AGEMA_reg_buffer_12296 ( .C (clk), .D (new_AGEMA_signal_33251), .Q (new_AGEMA_signal_33252) ) ;
    buf_clk new_AGEMA_reg_buffer_12300 ( .C (clk), .D (new_AGEMA_signal_33255), .Q (new_AGEMA_signal_33256) ) ;
    buf_clk new_AGEMA_reg_buffer_12304 ( .C (clk), .D (new_AGEMA_signal_33259), .Q (new_AGEMA_signal_33260) ) ;
    buf_clk new_AGEMA_reg_buffer_12308 ( .C (clk), .D (new_AGEMA_signal_33263), .Q (new_AGEMA_signal_33264) ) ;
    buf_clk new_AGEMA_reg_buffer_12312 ( .C (clk), .D (new_AGEMA_signal_33267), .Q (new_AGEMA_signal_33268) ) ;
    buf_clk new_AGEMA_reg_buffer_12316 ( .C (clk), .D (new_AGEMA_signal_33271), .Q (new_AGEMA_signal_33272) ) ;
    buf_clk new_AGEMA_reg_buffer_12320 ( .C (clk), .D (new_AGEMA_signal_33275), .Q (new_AGEMA_signal_33276) ) ;
    buf_clk new_AGEMA_reg_buffer_12324 ( .C (clk), .D (new_AGEMA_signal_33279), .Q (new_AGEMA_signal_33280) ) ;
    buf_clk new_AGEMA_reg_buffer_12328 ( .C (clk), .D (new_AGEMA_signal_33283), .Q (new_AGEMA_signal_33284) ) ;
    buf_clk new_AGEMA_reg_buffer_12332 ( .C (clk), .D (new_AGEMA_signal_33287), .Q (new_AGEMA_signal_33288) ) ;
    buf_clk new_AGEMA_reg_buffer_12336 ( .C (clk), .D (new_AGEMA_signal_33291), .Q (new_AGEMA_signal_33292) ) ;
    buf_clk new_AGEMA_reg_buffer_12340 ( .C (clk), .D (new_AGEMA_signal_33295), .Q (new_AGEMA_signal_33296) ) ;
    buf_clk new_AGEMA_reg_buffer_12344 ( .C (clk), .D (new_AGEMA_signal_33299), .Q (new_AGEMA_signal_33300) ) ;
    buf_clk new_AGEMA_reg_buffer_12348 ( .C (clk), .D (new_AGEMA_signal_33303), .Q (new_AGEMA_signal_33304) ) ;
    buf_clk new_AGEMA_reg_buffer_12352 ( .C (clk), .D (new_AGEMA_signal_33307), .Q (new_AGEMA_signal_33308) ) ;
    buf_clk new_AGEMA_reg_buffer_12356 ( .C (clk), .D (new_AGEMA_signal_33311), .Q (new_AGEMA_signal_33312) ) ;
    buf_clk new_AGEMA_reg_buffer_12360 ( .C (clk), .D (new_AGEMA_signal_33315), .Q (new_AGEMA_signal_33316) ) ;
    buf_clk new_AGEMA_reg_buffer_12364 ( .C (clk), .D (new_AGEMA_signal_33319), .Q (new_AGEMA_signal_33320) ) ;
    buf_clk new_AGEMA_reg_buffer_12368 ( .C (clk), .D (new_AGEMA_signal_33323), .Q (new_AGEMA_signal_33324) ) ;
    buf_clk new_AGEMA_reg_buffer_12372 ( .C (clk), .D (new_AGEMA_signal_33327), .Q (new_AGEMA_signal_33328) ) ;
    buf_clk new_AGEMA_reg_buffer_12376 ( .C (clk), .D (new_AGEMA_signal_33331), .Q (new_AGEMA_signal_33332) ) ;
    buf_clk new_AGEMA_reg_buffer_12380 ( .C (clk), .D (new_AGEMA_signal_33335), .Q (new_AGEMA_signal_33336) ) ;
    buf_clk new_AGEMA_reg_buffer_12384 ( .C (clk), .D (new_AGEMA_signal_33339), .Q (new_AGEMA_signal_33340) ) ;
    buf_clk new_AGEMA_reg_buffer_12388 ( .C (clk), .D (new_AGEMA_signal_33343), .Q (new_AGEMA_signal_33344) ) ;
    buf_clk new_AGEMA_reg_buffer_12392 ( .C (clk), .D (new_AGEMA_signal_33347), .Q (new_AGEMA_signal_33348) ) ;
    buf_clk new_AGEMA_reg_buffer_12396 ( .C (clk), .D (new_AGEMA_signal_33351), .Q (new_AGEMA_signal_33352) ) ;
    buf_clk new_AGEMA_reg_buffer_12400 ( .C (clk), .D (new_AGEMA_signal_33355), .Q (new_AGEMA_signal_33356) ) ;
    buf_clk new_AGEMA_reg_buffer_12404 ( .C (clk), .D (new_AGEMA_signal_33359), .Q (new_AGEMA_signal_33360) ) ;
    buf_clk new_AGEMA_reg_buffer_12408 ( .C (clk), .D (new_AGEMA_signal_33363), .Q (new_AGEMA_signal_33364) ) ;
    buf_clk new_AGEMA_reg_buffer_12412 ( .C (clk), .D (new_AGEMA_signal_33367), .Q (new_AGEMA_signal_33368) ) ;
    buf_clk new_AGEMA_reg_buffer_12416 ( .C (clk), .D (new_AGEMA_signal_33371), .Q (new_AGEMA_signal_33372) ) ;
    buf_clk new_AGEMA_reg_buffer_12420 ( .C (clk), .D (new_AGEMA_signal_33375), .Q (new_AGEMA_signal_33376) ) ;
    buf_clk new_AGEMA_reg_buffer_12424 ( .C (clk), .D (new_AGEMA_signal_33379), .Q (new_AGEMA_signal_33380) ) ;
    buf_clk new_AGEMA_reg_buffer_12428 ( .C (clk), .D (new_AGEMA_signal_33383), .Q (new_AGEMA_signal_33384) ) ;
    buf_clk new_AGEMA_reg_buffer_12432 ( .C (clk), .D (new_AGEMA_signal_33387), .Q (new_AGEMA_signal_33388) ) ;
    buf_clk new_AGEMA_reg_buffer_12436 ( .C (clk), .D (new_AGEMA_signal_33391), .Q (new_AGEMA_signal_33392) ) ;
    buf_clk new_AGEMA_reg_buffer_12440 ( .C (clk), .D (new_AGEMA_signal_33395), .Q (new_AGEMA_signal_33396) ) ;
    buf_clk new_AGEMA_reg_buffer_12444 ( .C (clk), .D (new_AGEMA_signal_33399), .Q (new_AGEMA_signal_33400) ) ;
    buf_clk new_AGEMA_reg_buffer_12448 ( .C (clk), .D (new_AGEMA_signal_33403), .Q (new_AGEMA_signal_33404) ) ;
    buf_clk new_AGEMA_reg_buffer_12452 ( .C (clk), .D (new_AGEMA_signal_33407), .Q (new_AGEMA_signal_33408) ) ;
    buf_clk new_AGEMA_reg_buffer_12456 ( .C (clk), .D (new_AGEMA_signal_33411), .Q (new_AGEMA_signal_33412) ) ;
    buf_clk new_AGEMA_reg_buffer_12460 ( .C (clk), .D (new_AGEMA_signal_33415), .Q (new_AGEMA_signal_33416) ) ;
    buf_clk new_AGEMA_reg_buffer_12464 ( .C (clk), .D (new_AGEMA_signal_33419), .Q (new_AGEMA_signal_33420) ) ;
    buf_clk new_AGEMA_reg_buffer_12468 ( .C (clk), .D (new_AGEMA_signal_33423), .Q (new_AGEMA_signal_33424) ) ;
    buf_clk new_AGEMA_reg_buffer_12472 ( .C (clk), .D (new_AGEMA_signal_33427), .Q (new_AGEMA_signal_33428) ) ;
    buf_clk new_AGEMA_reg_buffer_12476 ( .C (clk), .D (new_AGEMA_signal_33431), .Q (new_AGEMA_signal_33432) ) ;
    buf_clk new_AGEMA_reg_buffer_12480 ( .C (clk), .D (new_AGEMA_signal_33435), .Q (new_AGEMA_signal_33436) ) ;
    buf_clk new_AGEMA_reg_buffer_12484 ( .C (clk), .D (new_AGEMA_signal_33439), .Q (new_AGEMA_signal_33440) ) ;
    buf_clk new_AGEMA_reg_buffer_12488 ( .C (clk), .D (new_AGEMA_signal_33443), .Q (new_AGEMA_signal_33444) ) ;
    buf_clk new_AGEMA_reg_buffer_12492 ( .C (clk), .D (new_AGEMA_signal_33447), .Q (new_AGEMA_signal_33448) ) ;
    buf_clk new_AGEMA_reg_buffer_12496 ( .C (clk), .D (new_AGEMA_signal_33451), .Q (new_AGEMA_signal_33452) ) ;
    buf_clk new_AGEMA_reg_buffer_12500 ( .C (clk), .D (new_AGEMA_signal_33455), .Q (new_AGEMA_signal_33456) ) ;
    buf_clk new_AGEMA_reg_buffer_12504 ( .C (clk), .D (new_AGEMA_signal_33459), .Q (new_AGEMA_signal_33460) ) ;
    buf_clk new_AGEMA_reg_buffer_12508 ( .C (clk), .D (new_AGEMA_signal_33463), .Q (new_AGEMA_signal_33464) ) ;
    buf_clk new_AGEMA_reg_buffer_12512 ( .C (clk), .D (new_AGEMA_signal_33467), .Q (new_AGEMA_signal_33468) ) ;
    buf_clk new_AGEMA_reg_buffer_12516 ( .C (clk), .D (new_AGEMA_signal_33471), .Q (new_AGEMA_signal_33472) ) ;
    buf_clk new_AGEMA_reg_buffer_12520 ( .C (clk), .D (new_AGEMA_signal_33475), .Q (new_AGEMA_signal_33476) ) ;
    buf_clk new_AGEMA_reg_buffer_12524 ( .C (clk), .D (new_AGEMA_signal_33479), .Q (new_AGEMA_signal_33480) ) ;
    buf_clk new_AGEMA_reg_buffer_12528 ( .C (clk), .D (new_AGEMA_signal_33483), .Q (new_AGEMA_signal_33484) ) ;
    buf_clk new_AGEMA_reg_buffer_12532 ( .C (clk), .D (new_AGEMA_signal_33487), .Q (new_AGEMA_signal_33488) ) ;
    buf_clk new_AGEMA_reg_buffer_12536 ( .C (clk), .D (new_AGEMA_signal_33491), .Q (new_AGEMA_signal_33492) ) ;
    buf_clk new_AGEMA_reg_buffer_12540 ( .C (clk), .D (new_AGEMA_signal_33495), .Q (new_AGEMA_signal_33496) ) ;
    buf_clk new_AGEMA_reg_buffer_12544 ( .C (clk), .D (new_AGEMA_signal_33499), .Q (new_AGEMA_signal_33500) ) ;
    buf_clk new_AGEMA_reg_buffer_12548 ( .C (clk), .D (new_AGEMA_signal_33503), .Q (new_AGEMA_signal_33504) ) ;
    buf_clk new_AGEMA_reg_buffer_12552 ( .C (clk), .D (new_AGEMA_signal_33507), .Q (new_AGEMA_signal_33508) ) ;
    buf_clk new_AGEMA_reg_buffer_12556 ( .C (clk), .D (new_AGEMA_signal_33511), .Q (new_AGEMA_signal_33512) ) ;
    buf_clk new_AGEMA_reg_buffer_12560 ( .C (clk), .D (new_AGEMA_signal_33515), .Q (new_AGEMA_signal_33516) ) ;
    buf_clk new_AGEMA_reg_buffer_12564 ( .C (clk), .D (new_AGEMA_signal_33519), .Q (new_AGEMA_signal_33520) ) ;
    buf_clk new_AGEMA_reg_buffer_12568 ( .C (clk), .D (new_AGEMA_signal_33523), .Q (new_AGEMA_signal_33524) ) ;
    buf_clk new_AGEMA_reg_buffer_12572 ( .C (clk), .D (new_AGEMA_signal_33527), .Q (new_AGEMA_signal_33528) ) ;
    buf_clk new_AGEMA_reg_buffer_12576 ( .C (clk), .D (new_AGEMA_signal_33531), .Q (new_AGEMA_signal_33532) ) ;
    buf_clk new_AGEMA_reg_buffer_12580 ( .C (clk), .D (new_AGEMA_signal_33535), .Q (new_AGEMA_signal_33536) ) ;
    buf_clk new_AGEMA_reg_buffer_12584 ( .C (clk), .D (new_AGEMA_signal_33539), .Q (new_AGEMA_signal_33540) ) ;
    buf_clk new_AGEMA_reg_buffer_12588 ( .C (clk), .D (new_AGEMA_signal_33543), .Q (new_AGEMA_signal_33544) ) ;
    buf_clk new_AGEMA_reg_buffer_12592 ( .C (clk), .D (new_AGEMA_signal_33547), .Q (new_AGEMA_signal_33548) ) ;
    buf_clk new_AGEMA_reg_buffer_12596 ( .C (clk), .D (new_AGEMA_signal_33551), .Q (new_AGEMA_signal_33552) ) ;
    buf_clk new_AGEMA_reg_buffer_12600 ( .C (clk), .D (new_AGEMA_signal_33555), .Q (new_AGEMA_signal_33556) ) ;
    buf_clk new_AGEMA_reg_buffer_12604 ( .C (clk), .D (new_AGEMA_signal_33559), .Q (new_AGEMA_signal_33560) ) ;
    buf_clk new_AGEMA_reg_buffer_12608 ( .C (clk), .D (new_AGEMA_signal_33563), .Q (new_AGEMA_signal_33564) ) ;
    buf_clk new_AGEMA_reg_buffer_12612 ( .C (clk), .D (new_AGEMA_signal_33567), .Q (new_AGEMA_signal_33568) ) ;
    buf_clk new_AGEMA_reg_buffer_12616 ( .C (clk), .D (new_AGEMA_signal_33571), .Q (new_AGEMA_signal_33572) ) ;
    buf_clk new_AGEMA_reg_buffer_12620 ( .C (clk), .D (new_AGEMA_signal_33575), .Q (new_AGEMA_signal_33576) ) ;
    buf_clk new_AGEMA_reg_buffer_12624 ( .C (clk), .D (new_AGEMA_signal_33579), .Q (new_AGEMA_signal_33580) ) ;
    buf_clk new_AGEMA_reg_buffer_12628 ( .C (clk), .D (new_AGEMA_signal_33583), .Q (new_AGEMA_signal_33584) ) ;
    buf_clk new_AGEMA_reg_buffer_12632 ( .C (clk), .D (new_AGEMA_signal_33587), .Q (new_AGEMA_signal_33588) ) ;
    buf_clk new_AGEMA_reg_buffer_12636 ( .C (clk), .D (new_AGEMA_signal_33591), .Q (new_AGEMA_signal_33592) ) ;
    buf_clk new_AGEMA_reg_buffer_12640 ( .C (clk), .D (new_AGEMA_signal_33595), .Q (new_AGEMA_signal_33596) ) ;
    buf_clk new_AGEMA_reg_buffer_12644 ( .C (clk), .D (new_AGEMA_signal_33599), .Q (new_AGEMA_signal_33600) ) ;
    buf_clk new_AGEMA_reg_buffer_12648 ( .C (clk), .D (new_AGEMA_signal_33603), .Q (new_AGEMA_signal_33604) ) ;
    buf_clk new_AGEMA_reg_buffer_12652 ( .C (clk), .D (new_AGEMA_signal_33607), .Q (new_AGEMA_signal_33608) ) ;
    buf_clk new_AGEMA_reg_buffer_12656 ( .C (clk), .D (new_AGEMA_signal_33611), .Q (new_AGEMA_signal_33612) ) ;
    buf_clk new_AGEMA_reg_buffer_12660 ( .C (clk), .D (new_AGEMA_signal_33615), .Q (new_AGEMA_signal_33616) ) ;
    buf_clk new_AGEMA_reg_buffer_12664 ( .C (clk), .D (new_AGEMA_signal_33619), .Q (new_AGEMA_signal_33620) ) ;
    buf_clk new_AGEMA_reg_buffer_12668 ( .C (clk), .D (new_AGEMA_signal_33623), .Q (new_AGEMA_signal_33624) ) ;
    buf_clk new_AGEMA_reg_buffer_12672 ( .C (clk), .D (new_AGEMA_signal_33627), .Q (new_AGEMA_signal_33628) ) ;
    buf_clk new_AGEMA_reg_buffer_12676 ( .C (clk), .D (new_AGEMA_signal_33631), .Q (new_AGEMA_signal_33632) ) ;
    buf_clk new_AGEMA_reg_buffer_12680 ( .C (clk), .D (new_AGEMA_signal_33635), .Q (new_AGEMA_signal_33636) ) ;
    buf_clk new_AGEMA_reg_buffer_12684 ( .C (clk), .D (new_AGEMA_signal_33639), .Q (new_AGEMA_signal_33640) ) ;
    buf_clk new_AGEMA_reg_buffer_12688 ( .C (clk), .D (new_AGEMA_signal_33643), .Q (new_AGEMA_signal_33644) ) ;
    buf_clk new_AGEMA_reg_buffer_12692 ( .C (clk), .D (new_AGEMA_signal_33647), .Q (new_AGEMA_signal_33648) ) ;
    buf_clk new_AGEMA_reg_buffer_12696 ( .C (clk), .D (new_AGEMA_signal_33651), .Q (new_AGEMA_signal_33652) ) ;
    buf_clk new_AGEMA_reg_buffer_12700 ( .C (clk), .D (new_AGEMA_signal_33655), .Q (new_AGEMA_signal_33656) ) ;
    buf_clk new_AGEMA_reg_buffer_12704 ( .C (clk), .D (new_AGEMA_signal_33659), .Q (new_AGEMA_signal_33660) ) ;
    buf_clk new_AGEMA_reg_buffer_12708 ( .C (clk), .D (new_AGEMA_signal_33663), .Q (new_AGEMA_signal_33664) ) ;
    buf_clk new_AGEMA_reg_buffer_12712 ( .C (clk), .D (new_AGEMA_signal_33667), .Q (new_AGEMA_signal_33668) ) ;
    buf_clk new_AGEMA_reg_buffer_12716 ( .C (clk), .D (new_AGEMA_signal_33671), .Q (new_AGEMA_signal_33672) ) ;
    buf_clk new_AGEMA_reg_buffer_12720 ( .C (clk), .D (new_AGEMA_signal_33675), .Q (new_AGEMA_signal_33676) ) ;
    buf_clk new_AGEMA_reg_buffer_12724 ( .C (clk), .D (new_AGEMA_signal_33679), .Q (new_AGEMA_signal_33680) ) ;
    buf_clk new_AGEMA_reg_buffer_12728 ( .C (clk), .D (new_AGEMA_signal_33683), .Q (new_AGEMA_signal_33684) ) ;
    buf_clk new_AGEMA_reg_buffer_12732 ( .C (clk), .D (new_AGEMA_signal_33687), .Q (new_AGEMA_signal_33688) ) ;
    buf_clk new_AGEMA_reg_buffer_12736 ( .C (clk), .D (new_AGEMA_signal_33691), .Q (new_AGEMA_signal_33692) ) ;
    buf_clk new_AGEMA_reg_buffer_12740 ( .C (clk), .D (new_AGEMA_signal_33695), .Q (new_AGEMA_signal_33696) ) ;
    buf_clk new_AGEMA_reg_buffer_12744 ( .C (clk), .D (new_AGEMA_signal_33699), .Q (new_AGEMA_signal_33700) ) ;
    buf_clk new_AGEMA_reg_buffer_12748 ( .C (clk), .D (new_AGEMA_signal_33703), .Q (new_AGEMA_signal_33704) ) ;
    buf_clk new_AGEMA_reg_buffer_12752 ( .C (clk), .D (new_AGEMA_signal_33707), .Q (new_AGEMA_signal_33708) ) ;
    buf_clk new_AGEMA_reg_buffer_12756 ( .C (clk), .D (new_AGEMA_signal_33711), .Q (new_AGEMA_signal_33712) ) ;
    buf_clk new_AGEMA_reg_buffer_12760 ( .C (clk), .D (new_AGEMA_signal_33715), .Q (new_AGEMA_signal_33716) ) ;
    buf_clk new_AGEMA_reg_buffer_12764 ( .C (clk), .D (new_AGEMA_signal_33719), .Q (new_AGEMA_signal_33720) ) ;
    buf_clk new_AGEMA_reg_buffer_12768 ( .C (clk), .D (new_AGEMA_signal_33723), .Q (new_AGEMA_signal_33724) ) ;
    buf_clk new_AGEMA_reg_buffer_12772 ( .C (clk), .D (new_AGEMA_signal_33727), .Q (new_AGEMA_signal_33728) ) ;
    buf_clk new_AGEMA_reg_buffer_12776 ( .C (clk), .D (new_AGEMA_signal_33731), .Q (new_AGEMA_signal_33732) ) ;
    buf_clk new_AGEMA_reg_buffer_12780 ( .C (clk), .D (new_AGEMA_signal_33735), .Q (new_AGEMA_signal_33736) ) ;
    buf_clk new_AGEMA_reg_buffer_12784 ( .C (clk), .D (new_AGEMA_signal_33739), .Q (new_AGEMA_signal_33740) ) ;
    buf_clk new_AGEMA_reg_buffer_12788 ( .C (clk), .D (new_AGEMA_signal_33743), .Q (new_AGEMA_signal_33744) ) ;
    buf_clk new_AGEMA_reg_buffer_12792 ( .C (clk), .D (new_AGEMA_signal_33747), .Q (new_AGEMA_signal_33748) ) ;
    buf_clk new_AGEMA_reg_buffer_12796 ( .C (clk), .D (new_AGEMA_signal_33751), .Q (new_AGEMA_signal_33752) ) ;
    buf_clk new_AGEMA_reg_buffer_12800 ( .C (clk), .D (new_AGEMA_signal_33755), .Q (new_AGEMA_signal_33756) ) ;
    buf_clk new_AGEMA_reg_buffer_12804 ( .C (clk), .D (new_AGEMA_signal_33759), .Q (new_AGEMA_signal_33760) ) ;
    buf_clk new_AGEMA_reg_buffer_12808 ( .C (clk), .D (new_AGEMA_signal_33763), .Q (new_AGEMA_signal_33764) ) ;
    buf_clk new_AGEMA_reg_buffer_12812 ( .C (clk), .D (new_AGEMA_signal_33767), .Q (new_AGEMA_signal_33768) ) ;
    buf_clk new_AGEMA_reg_buffer_12816 ( .C (clk), .D (new_AGEMA_signal_33771), .Q (new_AGEMA_signal_33772) ) ;
    buf_clk new_AGEMA_reg_buffer_12820 ( .C (clk), .D (new_AGEMA_signal_33775), .Q (new_AGEMA_signal_33776) ) ;
    buf_clk new_AGEMA_reg_buffer_12824 ( .C (clk), .D (new_AGEMA_signal_33779), .Q (new_AGEMA_signal_33780) ) ;
    buf_clk new_AGEMA_reg_buffer_12828 ( .C (clk), .D (new_AGEMA_signal_33783), .Q (new_AGEMA_signal_33784) ) ;
    buf_clk new_AGEMA_reg_buffer_12832 ( .C (clk), .D (new_AGEMA_signal_33787), .Q (new_AGEMA_signal_33788) ) ;
    buf_clk new_AGEMA_reg_buffer_12836 ( .C (clk), .D (new_AGEMA_signal_33791), .Q (new_AGEMA_signal_33792) ) ;
    buf_clk new_AGEMA_reg_buffer_12840 ( .C (clk), .D (new_AGEMA_signal_33795), .Q (new_AGEMA_signal_33796) ) ;
    buf_clk new_AGEMA_reg_buffer_12844 ( .C (clk), .D (new_AGEMA_signal_33799), .Q (new_AGEMA_signal_33800) ) ;
    buf_clk new_AGEMA_reg_buffer_12848 ( .C (clk), .D (new_AGEMA_signal_33803), .Q (new_AGEMA_signal_33804) ) ;
    buf_clk new_AGEMA_reg_buffer_12852 ( .C (clk), .D (new_AGEMA_signal_33807), .Q (new_AGEMA_signal_33808) ) ;
    buf_clk new_AGEMA_reg_buffer_12856 ( .C (clk), .D (new_AGEMA_signal_33811), .Q (new_AGEMA_signal_33812) ) ;
    buf_clk new_AGEMA_reg_buffer_12860 ( .C (clk), .D (new_AGEMA_signal_33815), .Q (new_AGEMA_signal_33816) ) ;
    buf_clk new_AGEMA_reg_buffer_12864 ( .C (clk), .D (new_AGEMA_signal_33819), .Q (new_AGEMA_signal_33820) ) ;
    buf_clk new_AGEMA_reg_buffer_12868 ( .C (clk), .D (new_AGEMA_signal_33823), .Q (new_AGEMA_signal_33824) ) ;
    buf_clk new_AGEMA_reg_buffer_12872 ( .C (clk), .D (new_AGEMA_signal_33827), .Q (new_AGEMA_signal_33828) ) ;
    buf_clk new_AGEMA_reg_buffer_12876 ( .C (clk), .D (new_AGEMA_signal_33831), .Q (new_AGEMA_signal_33832) ) ;
    buf_clk new_AGEMA_reg_buffer_12880 ( .C (clk), .D (new_AGEMA_signal_33835), .Q (new_AGEMA_signal_33836) ) ;
    buf_clk new_AGEMA_reg_buffer_12884 ( .C (clk), .D (new_AGEMA_signal_33839), .Q (new_AGEMA_signal_33840) ) ;
    buf_clk new_AGEMA_reg_buffer_12888 ( .C (clk), .D (new_AGEMA_signal_33843), .Q (new_AGEMA_signal_33844) ) ;
    buf_clk new_AGEMA_reg_buffer_12892 ( .C (clk), .D (new_AGEMA_signal_33847), .Q (new_AGEMA_signal_33848) ) ;
    buf_clk new_AGEMA_reg_buffer_12896 ( .C (clk), .D (new_AGEMA_signal_33851), .Q (new_AGEMA_signal_33852) ) ;
    buf_clk new_AGEMA_reg_buffer_12900 ( .C (clk), .D (new_AGEMA_signal_33855), .Q (new_AGEMA_signal_33856) ) ;
    buf_clk new_AGEMA_reg_buffer_12904 ( .C (clk), .D (new_AGEMA_signal_33859), .Q (new_AGEMA_signal_33860) ) ;
    buf_clk new_AGEMA_reg_buffer_12908 ( .C (clk), .D (new_AGEMA_signal_33863), .Q (new_AGEMA_signal_33864) ) ;
    buf_clk new_AGEMA_reg_buffer_12912 ( .C (clk), .D (new_AGEMA_signal_33867), .Q (new_AGEMA_signal_33868) ) ;
    buf_clk new_AGEMA_reg_buffer_12916 ( .C (clk), .D (new_AGEMA_signal_33871), .Q (new_AGEMA_signal_33872) ) ;
    buf_clk new_AGEMA_reg_buffer_12920 ( .C (clk), .D (new_AGEMA_signal_33875), .Q (new_AGEMA_signal_33876) ) ;
    buf_clk new_AGEMA_reg_buffer_12924 ( .C (clk), .D (new_AGEMA_signal_33879), .Q (new_AGEMA_signal_33880) ) ;
    buf_clk new_AGEMA_reg_buffer_12928 ( .C (clk), .D (new_AGEMA_signal_33883), .Q (new_AGEMA_signal_33884) ) ;
    buf_clk new_AGEMA_reg_buffer_12932 ( .C (clk), .D (new_AGEMA_signal_33887), .Q (new_AGEMA_signal_33888) ) ;
    buf_clk new_AGEMA_reg_buffer_12936 ( .C (clk), .D (new_AGEMA_signal_33891), .Q (new_AGEMA_signal_33892) ) ;
    buf_clk new_AGEMA_reg_buffer_12940 ( .C (clk), .D (new_AGEMA_signal_33895), .Q (new_AGEMA_signal_33896) ) ;
    buf_clk new_AGEMA_reg_buffer_12944 ( .C (clk), .D (new_AGEMA_signal_33899), .Q (new_AGEMA_signal_33900) ) ;
    buf_clk new_AGEMA_reg_buffer_12948 ( .C (clk), .D (new_AGEMA_signal_33903), .Q (new_AGEMA_signal_33904) ) ;
    buf_clk new_AGEMA_reg_buffer_12952 ( .C (clk), .D (new_AGEMA_signal_33907), .Q (new_AGEMA_signal_33908) ) ;
    buf_clk new_AGEMA_reg_buffer_12956 ( .C (clk), .D (new_AGEMA_signal_33911), .Q (new_AGEMA_signal_33912) ) ;
    buf_clk new_AGEMA_reg_buffer_12960 ( .C (clk), .D (new_AGEMA_signal_33915), .Q (new_AGEMA_signal_33916) ) ;
    buf_clk new_AGEMA_reg_buffer_12964 ( .C (clk), .D (new_AGEMA_signal_33919), .Q (new_AGEMA_signal_33920) ) ;
    buf_clk new_AGEMA_reg_buffer_12968 ( .C (clk), .D (new_AGEMA_signal_33923), .Q (new_AGEMA_signal_33924) ) ;
    buf_clk new_AGEMA_reg_buffer_12972 ( .C (clk), .D (new_AGEMA_signal_33927), .Q (new_AGEMA_signal_33928) ) ;
    buf_clk new_AGEMA_reg_buffer_12976 ( .C (clk), .D (new_AGEMA_signal_33931), .Q (new_AGEMA_signal_33932) ) ;
    buf_clk new_AGEMA_reg_buffer_12980 ( .C (clk), .D (new_AGEMA_signal_33935), .Q (new_AGEMA_signal_33936) ) ;
    buf_clk new_AGEMA_reg_buffer_12984 ( .C (clk), .D (new_AGEMA_signal_33939), .Q (new_AGEMA_signal_33940) ) ;
    buf_clk new_AGEMA_reg_buffer_12988 ( .C (clk), .D (new_AGEMA_signal_33943), .Q (new_AGEMA_signal_33944) ) ;
    buf_clk new_AGEMA_reg_buffer_12992 ( .C (clk), .D (new_AGEMA_signal_33947), .Q (new_AGEMA_signal_33948) ) ;
    buf_clk new_AGEMA_reg_buffer_12996 ( .C (clk), .D (new_AGEMA_signal_33951), .Q (new_AGEMA_signal_33952) ) ;
    buf_clk new_AGEMA_reg_buffer_13000 ( .C (clk), .D (new_AGEMA_signal_33955), .Q (new_AGEMA_signal_33956) ) ;
    buf_clk new_AGEMA_reg_buffer_13004 ( .C (clk), .D (new_AGEMA_signal_33959), .Q (new_AGEMA_signal_33960) ) ;
    buf_clk new_AGEMA_reg_buffer_13008 ( .C (clk), .D (new_AGEMA_signal_33963), .Q (new_AGEMA_signal_33964) ) ;
    buf_clk new_AGEMA_reg_buffer_13012 ( .C (clk), .D (new_AGEMA_signal_33967), .Q (new_AGEMA_signal_33968) ) ;
    buf_clk new_AGEMA_reg_buffer_13016 ( .C (clk), .D (new_AGEMA_signal_33971), .Q (new_AGEMA_signal_33972) ) ;
    buf_clk new_AGEMA_reg_buffer_13020 ( .C (clk), .D (new_AGEMA_signal_33975), .Q (new_AGEMA_signal_33976) ) ;
    buf_clk new_AGEMA_reg_buffer_13024 ( .C (clk), .D (new_AGEMA_signal_33979), .Q (new_AGEMA_signal_33980) ) ;
    buf_clk new_AGEMA_reg_buffer_13028 ( .C (clk), .D (new_AGEMA_signal_33983), .Q (new_AGEMA_signal_33984) ) ;
    buf_clk new_AGEMA_reg_buffer_13032 ( .C (clk), .D (new_AGEMA_signal_33987), .Q (new_AGEMA_signal_33988) ) ;
    buf_clk new_AGEMA_reg_buffer_13036 ( .C (clk), .D (new_AGEMA_signal_33991), .Q (new_AGEMA_signal_33992) ) ;
    buf_clk new_AGEMA_reg_buffer_13040 ( .C (clk), .D (new_AGEMA_signal_33995), .Q (new_AGEMA_signal_33996) ) ;
    buf_clk new_AGEMA_reg_buffer_13044 ( .C (clk), .D (new_AGEMA_signal_33999), .Q (new_AGEMA_signal_34000) ) ;
    buf_clk new_AGEMA_reg_buffer_13048 ( .C (clk), .D (new_AGEMA_signal_34003), .Q (new_AGEMA_signal_34004) ) ;
    buf_clk new_AGEMA_reg_buffer_13052 ( .C (clk), .D (new_AGEMA_signal_34007), .Q (new_AGEMA_signal_34008) ) ;
    buf_clk new_AGEMA_reg_buffer_13056 ( .C (clk), .D (new_AGEMA_signal_34011), .Q (new_AGEMA_signal_34012) ) ;
    buf_clk new_AGEMA_reg_buffer_13060 ( .C (clk), .D (new_AGEMA_signal_34015), .Q (new_AGEMA_signal_34016) ) ;
    buf_clk new_AGEMA_reg_buffer_13064 ( .C (clk), .D (new_AGEMA_signal_34019), .Q (new_AGEMA_signal_34020) ) ;
    buf_clk new_AGEMA_reg_buffer_13068 ( .C (clk), .D (new_AGEMA_signal_34023), .Q (new_AGEMA_signal_34024) ) ;
    buf_clk new_AGEMA_reg_buffer_13072 ( .C (clk), .D (new_AGEMA_signal_34027), .Q (new_AGEMA_signal_34028) ) ;
    buf_clk new_AGEMA_reg_buffer_13076 ( .C (clk), .D (new_AGEMA_signal_34031), .Q (new_AGEMA_signal_34032) ) ;
    buf_clk new_AGEMA_reg_buffer_13080 ( .C (clk), .D (new_AGEMA_signal_34035), .Q (new_AGEMA_signal_34036) ) ;
    buf_clk new_AGEMA_reg_buffer_13084 ( .C (clk), .D (new_AGEMA_signal_34039), .Q (new_AGEMA_signal_34040) ) ;
    buf_clk new_AGEMA_reg_buffer_13088 ( .C (clk), .D (new_AGEMA_signal_34043), .Q (new_AGEMA_signal_34044) ) ;
    buf_clk new_AGEMA_reg_buffer_13092 ( .C (clk), .D (new_AGEMA_signal_34047), .Q (new_AGEMA_signal_34048) ) ;
    buf_clk new_AGEMA_reg_buffer_13096 ( .C (clk), .D (new_AGEMA_signal_34051), .Q (new_AGEMA_signal_34052) ) ;
    buf_clk new_AGEMA_reg_buffer_13100 ( .C (clk), .D (new_AGEMA_signal_34055), .Q (new_AGEMA_signal_34056) ) ;
    buf_clk new_AGEMA_reg_buffer_13104 ( .C (clk), .D (new_AGEMA_signal_34059), .Q (new_AGEMA_signal_34060) ) ;
    buf_clk new_AGEMA_reg_buffer_13108 ( .C (clk), .D (new_AGEMA_signal_34063), .Q (new_AGEMA_signal_34064) ) ;
    buf_clk new_AGEMA_reg_buffer_13112 ( .C (clk), .D (new_AGEMA_signal_34067), .Q (new_AGEMA_signal_34068) ) ;
    buf_clk new_AGEMA_reg_buffer_13116 ( .C (clk), .D (new_AGEMA_signal_34071), .Q (new_AGEMA_signal_34072) ) ;
    buf_clk new_AGEMA_reg_buffer_13120 ( .C (clk), .D (new_AGEMA_signal_34075), .Q (new_AGEMA_signal_34076) ) ;
    buf_clk new_AGEMA_reg_buffer_13124 ( .C (clk), .D (new_AGEMA_signal_34079), .Q (new_AGEMA_signal_34080) ) ;
    buf_clk new_AGEMA_reg_buffer_13128 ( .C (clk), .D (new_AGEMA_signal_34083), .Q (new_AGEMA_signal_34084) ) ;
    buf_clk new_AGEMA_reg_buffer_13132 ( .C (clk), .D (new_AGEMA_signal_34087), .Q (new_AGEMA_signal_34088) ) ;
    buf_clk new_AGEMA_reg_buffer_13136 ( .C (clk), .D (new_AGEMA_signal_34091), .Q (new_AGEMA_signal_34092) ) ;
    buf_clk new_AGEMA_reg_buffer_13140 ( .C (clk), .D (new_AGEMA_signal_34095), .Q (new_AGEMA_signal_34096) ) ;
    buf_clk new_AGEMA_reg_buffer_13144 ( .C (clk), .D (new_AGEMA_signal_34099), .Q (new_AGEMA_signal_34100) ) ;
    buf_clk new_AGEMA_reg_buffer_13148 ( .C (clk), .D (new_AGEMA_signal_34103), .Q (new_AGEMA_signal_34104) ) ;
    buf_clk new_AGEMA_reg_buffer_13152 ( .C (clk), .D (new_AGEMA_signal_34107), .Q (new_AGEMA_signal_34108) ) ;
    buf_clk new_AGEMA_reg_buffer_13156 ( .C (clk), .D (new_AGEMA_signal_34111), .Q (new_AGEMA_signal_34112) ) ;
    buf_clk new_AGEMA_reg_buffer_13160 ( .C (clk), .D (new_AGEMA_signal_34115), .Q (new_AGEMA_signal_34116) ) ;
    buf_clk new_AGEMA_reg_buffer_13164 ( .C (clk), .D (new_AGEMA_signal_34119), .Q (new_AGEMA_signal_34120) ) ;
    buf_clk new_AGEMA_reg_buffer_13168 ( .C (clk), .D (new_AGEMA_signal_34123), .Q (new_AGEMA_signal_34124) ) ;
    buf_clk new_AGEMA_reg_buffer_13172 ( .C (clk), .D (new_AGEMA_signal_34127), .Q (new_AGEMA_signal_34128) ) ;
    buf_clk new_AGEMA_reg_buffer_13176 ( .C (clk), .D (new_AGEMA_signal_34131), .Q (new_AGEMA_signal_34132) ) ;
    buf_clk new_AGEMA_reg_buffer_13180 ( .C (clk), .D (new_AGEMA_signal_34135), .Q (new_AGEMA_signal_34136) ) ;
    buf_clk new_AGEMA_reg_buffer_13184 ( .C (clk), .D (new_AGEMA_signal_34139), .Q (new_AGEMA_signal_34140) ) ;
    buf_clk new_AGEMA_reg_buffer_13188 ( .C (clk), .D (new_AGEMA_signal_34143), .Q (new_AGEMA_signal_34144) ) ;
    buf_clk new_AGEMA_reg_buffer_13192 ( .C (clk), .D (new_AGEMA_signal_34147), .Q (new_AGEMA_signal_34148) ) ;
    buf_clk new_AGEMA_reg_buffer_13196 ( .C (clk), .D (new_AGEMA_signal_34151), .Q (new_AGEMA_signal_34152) ) ;
    buf_clk new_AGEMA_reg_buffer_13200 ( .C (clk), .D (new_AGEMA_signal_34155), .Q (new_AGEMA_signal_34156) ) ;
    buf_clk new_AGEMA_reg_buffer_13204 ( .C (clk), .D (new_AGEMA_signal_34159), .Q (new_AGEMA_signal_34160) ) ;
    buf_clk new_AGEMA_reg_buffer_13208 ( .C (clk), .D (new_AGEMA_signal_34163), .Q (new_AGEMA_signal_34164) ) ;
    buf_clk new_AGEMA_reg_buffer_13212 ( .C (clk), .D (new_AGEMA_signal_34167), .Q (new_AGEMA_signal_34168) ) ;
    buf_clk new_AGEMA_reg_buffer_13216 ( .C (clk), .D (new_AGEMA_signal_34171), .Q (new_AGEMA_signal_34172) ) ;
    buf_clk new_AGEMA_reg_buffer_13220 ( .C (clk), .D (new_AGEMA_signal_34175), .Q (new_AGEMA_signal_34176) ) ;
    buf_clk new_AGEMA_reg_buffer_13224 ( .C (clk), .D (new_AGEMA_signal_34179), .Q (new_AGEMA_signal_34180) ) ;
    buf_clk new_AGEMA_reg_buffer_13228 ( .C (clk), .D (new_AGEMA_signal_34183), .Q (new_AGEMA_signal_34184) ) ;
    buf_clk new_AGEMA_reg_buffer_13232 ( .C (clk), .D (new_AGEMA_signal_34187), .Q (new_AGEMA_signal_34188) ) ;
    buf_clk new_AGEMA_reg_buffer_13236 ( .C (clk), .D (new_AGEMA_signal_34191), .Q (new_AGEMA_signal_34192) ) ;
    buf_clk new_AGEMA_reg_buffer_13240 ( .C (clk), .D (new_AGEMA_signal_34195), .Q (new_AGEMA_signal_34196) ) ;
    buf_clk new_AGEMA_reg_buffer_13244 ( .C (clk), .D (new_AGEMA_signal_34199), .Q (new_AGEMA_signal_34200) ) ;
    buf_clk new_AGEMA_reg_buffer_13248 ( .C (clk), .D (new_AGEMA_signal_34203), .Q (new_AGEMA_signal_34204) ) ;
    buf_clk new_AGEMA_reg_buffer_13252 ( .C (clk), .D (new_AGEMA_signal_34207), .Q (new_AGEMA_signal_34208) ) ;
    buf_clk new_AGEMA_reg_buffer_13256 ( .C (clk), .D (new_AGEMA_signal_34211), .Q (new_AGEMA_signal_34212) ) ;
    buf_clk new_AGEMA_reg_buffer_13260 ( .C (clk), .D (new_AGEMA_signal_34215), .Q (new_AGEMA_signal_34216) ) ;
    buf_clk new_AGEMA_reg_buffer_13264 ( .C (clk), .D (new_AGEMA_signal_34219), .Q (new_AGEMA_signal_34220) ) ;
    buf_clk new_AGEMA_reg_buffer_13268 ( .C (clk), .D (new_AGEMA_signal_34223), .Q (new_AGEMA_signal_34224) ) ;
    buf_clk new_AGEMA_reg_buffer_13272 ( .C (clk), .D (new_AGEMA_signal_34227), .Q (new_AGEMA_signal_34228) ) ;
    buf_clk new_AGEMA_reg_buffer_13276 ( .C (clk), .D (new_AGEMA_signal_34231), .Q (new_AGEMA_signal_34232) ) ;
    buf_clk new_AGEMA_reg_buffer_13280 ( .C (clk), .D (new_AGEMA_signal_34235), .Q (new_AGEMA_signal_34236) ) ;
    buf_clk new_AGEMA_reg_buffer_13284 ( .C (clk), .D (new_AGEMA_signal_34239), .Q (new_AGEMA_signal_34240) ) ;
    buf_clk new_AGEMA_reg_buffer_13288 ( .C (clk), .D (new_AGEMA_signal_34243), .Q (new_AGEMA_signal_34244) ) ;
    buf_clk new_AGEMA_reg_buffer_13292 ( .C (clk), .D (new_AGEMA_signal_34247), .Q (new_AGEMA_signal_34248) ) ;
    buf_clk new_AGEMA_reg_buffer_13296 ( .C (clk), .D (new_AGEMA_signal_34251), .Q (new_AGEMA_signal_34252) ) ;
    buf_clk new_AGEMA_reg_buffer_13300 ( .C (clk), .D (new_AGEMA_signal_34255), .Q (new_AGEMA_signal_34256) ) ;
    buf_clk new_AGEMA_reg_buffer_13304 ( .C (clk), .D (new_AGEMA_signal_34259), .Q (new_AGEMA_signal_34260) ) ;
    buf_clk new_AGEMA_reg_buffer_13308 ( .C (clk), .D (new_AGEMA_signal_34263), .Q (new_AGEMA_signal_34264) ) ;
    buf_clk new_AGEMA_reg_buffer_13312 ( .C (clk), .D (new_AGEMA_signal_34267), .Q (new_AGEMA_signal_34268) ) ;
    buf_clk new_AGEMA_reg_buffer_13316 ( .C (clk), .D (new_AGEMA_signal_34271), .Q (new_AGEMA_signal_34272) ) ;
    buf_clk new_AGEMA_reg_buffer_13320 ( .C (clk), .D (new_AGEMA_signal_34275), .Q (new_AGEMA_signal_34276) ) ;
    buf_clk new_AGEMA_reg_buffer_13324 ( .C (clk), .D (new_AGEMA_signal_34279), .Q (new_AGEMA_signal_34280) ) ;
    buf_clk new_AGEMA_reg_buffer_13328 ( .C (clk), .D (new_AGEMA_signal_34283), .Q (new_AGEMA_signal_34284) ) ;
    buf_clk new_AGEMA_reg_buffer_13332 ( .C (clk), .D (new_AGEMA_signal_34287), .Q (new_AGEMA_signal_34288) ) ;
    buf_clk new_AGEMA_reg_buffer_13336 ( .C (clk), .D (new_AGEMA_signal_34291), .Q (new_AGEMA_signal_34292) ) ;
    buf_clk new_AGEMA_reg_buffer_13340 ( .C (clk), .D (new_AGEMA_signal_34295), .Q (new_AGEMA_signal_34296) ) ;
    buf_clk new_AGEMA_reg_buffer_13344 ( .C (clk), .D (new_AGEMA_signal_34299), .Q (new_AGEMA_signal_34300) ) ;
    buf_clk new_AGEMA_reg_buffer_13348 ( .C (clk), .D (new_AGEMA_signal_34303), .Q (new_AGEMA_signal_34304) ) ;
    buf_clk new_AGEMA_reg_buffer_13352 ( .C (clk), .D (new_AGEMA_signal_34307), .Q (new_AGEMA_signal_34308) ) ;
    buf_clk new_AGEMA_reg_buffer_13356 ( .C (clk), .D (new_AGEMA_signal_34311), .Q (new_AGEMA_signal_34312) ) ;
    buf_clk new_AGEMA_reg_buffer_13360 ( .C (clk), .D (new_AGEMA_signal_34315), .Q (new_AGEMA_signal_34316) ) ;
    buf_clk new_AGEMA_reg_buffer_13364 ( .C (clk), .D (new_AGEMA_signal_34319), .Q (new_AGEMA_signal_34320) ) ;
    buf_clk new_AGEMA_reg_buffer_13368 ( .C (clk), .D (new_AGEMA_signal_34323), .Q (new_AGEMA_signal_34324) ) ;
    buf_clk new_AGEMA_reg_buffer_13372 ( .C (clk), .D (new_AGEMA_signal_34327), .Q (new_AGEMA_signal_34328) ) ;
    buf_clk new_AGEMA_reg_buffer_13376 ( .C (clk), .D (new_AGEMA_signal_34331), .Q (new_AGEMA_signal_34332) ) ;
    buf_clk new_AGEMA_reg_buffer_13380 ( .C (clk), .D (new_AGEMA_signal_34335), .Q (new_AGEMA_signal_34336) ) ;
    buf_clk new_AGEMA_reg_buffer_13384 ( .C (clk), .D (new_AGEMA_signal_34339), .Q (new_AGEMA_signal_34340) ) ;
    buf_clk new_AGEMA_reg_buffer_13388 ( .C (clk), .D (new_AGEMA_signal_34343), .Q (new_AGEMA_signal_34344) ) ;
    buf_clk new_AGEMA_reg_buffer_13392 ( .C (clk), .D (new_AGEMA_signal_34347), .Q (new_AGEMA_signal_34348) ) ;
    buf_clk new_AGEMA_reg_buffer_13396 ( .C (clk), .D (new_AGEMA_signal_34351), .Q (new_AGEMA_signal_34352) ) ;
    buf_clk new_AGEMA_reg_buffer_13400 ( .C (clk), .D (new_AGEMA_signal_34355), .Q (new_AGEMA_signal_34356) ) ;
    buf_clk new_AGEMA_reg_buffer_13404 ( .C (clk), .D (new_AGEMA_signal_34359), .Q (new_AGEMA_signal_34360) ) ;
    buf_clk new_AGEMA_reg_buffer_13408 ( .C (clk), .D (new_AGEMA_signal_34363), .Q (new_AGEMA_signal_34364) ) ;
    buf_clk new_AGEMA_reg_buffer_13412 ( .C (clk), .D (new_AGEMA_signal_34367), .Q (new_AGEMA_signal_34368) ) ;
    buf_clk new_AGEMA_reg_buffer_13416 ( .C (clk), .D (new_AGEMA_signal_34371), .Q (new_AGEMA_signal_34372) ) ;
    buf_clk new_AGEMA_reg_buffer_13420 ( .C (clk), .D (new_AGEMA_signal_34375), .Q (new_AGEMA_signal_34376) ) ;
    buf_clk new_AGEMA_reg_buffer_13424 ( .C (clk), .D (new_AGEMA_signal_34379), .Q (new_AGEMA_signal_34380) ) ;
    buf_clk new_AGEMA_reg_buffer_13428 ( .C (clk), .D (new_AGEMA_signal_34383), .Q (new_AGEMA_signal_34384) ) ;
    buf_clk new_AGEMA_reg_buffer_13432 ( .C (clk), .D (new_AGEMA_signal_34387), .Q (new_AGEMA_signal_34388) ) ;
    buf_clk new_AGEMA_reg_buffer_13436 ( .C (clk), .D (new_AGEMA_signal_34391), .Q (new_AGEMA_signal_34392) ) ;
    buf_clk new_AGEMA_reg_buffer_13440 ( .C (clk), .D (new_AGEMA_signal_34395), .Q (new_AGEMA_signal_34396) ) ;
    buf_clk new_AGEMA_reg_buffer_13444 ( .C (clk), .D (new_AGEMA_signal_34399), .Q (new_AGEMA_signal_34400) ) ;
    buf_clk new_AGEMA_reg_buffer_13448 ( .C (clk), .D (new_AGEMA_signal_34403), .Q (new_AGEMA_signal_34404) ) ;
    buf_clk new_AGEMA_reg_buffer_13452 ( .C (clk), .D (new_AGEMA_signal_34407), .Q (new_AGEMA_signal_34408) ) ;
    buf_clk new_AGEMA_reg_buffer_13456 ( .C (clk), .D (new_AGEMA_signal_34411), .Q (new_AGEMA_signal_34412) ) ;
    buf_clk new_AGEMA_reg_buffer_13460 ( .C (clk), .D (new_AGEMA_signal_34415), .Q (new_AGEMA_signal_34416) ) ;
    buf_clk new_AGEMA_reg_buffer_13464 ( .C (clk), .D (new_AGEMA_signal_34419), .Q (new_AGEMA_signal_34420) ) ;
    buf_clk new_AGEMA_reg_buffer_13468 ( .C (clk), .D (new_AGEMA_signal_34423), .Q (new_AGEMA_signal_34424) ) ;
    buf_clk new_AGEMA_reg_buffer_13472 ( .C (clk), .D (new_AGEMA_signal_34427), .Q (new_AGEMA_signal_34428) ) ;
    buf_clk new_AGEMA_reg_buffer_13476 ( .C (clk), .D (new_AGEMA_signal_34431), .Q (new_AGEMA_signal_34432) ) ;
    buf_clk new_AGEMA_reg_buffer_13480 ( .C (clk), .D (new_AGEMA_signal_34435), .Q (new_AGEMA_signal_34436) ) ;
    buf_clk new_AGEMA_reg_buffer_13484 ( .C (clk), .D (new_AGEMA_signal_34439), .Q (new_AGEMA_signal_34440) ) ;
    buf_clk new_AGEMA_reg_buffer_13488 ( .C (clk), .D (new_AGEMA_signal_34443), .Q (new_AGEMA_signal_34444) ) ;
    buf_clk new_AGEMA_reg_buffer_13492 ( .C (clk), .D (new_AGEMA_signal_34447), .Q (new_AGEMA_signal_34448) ) ;
    buf_clk new_AGEMA_reg_buffer_13496 ( .C (clk), .D (new_AGEMA_signal_34451), .Q (new_AGEMA_signal_34452) ) ;
    buf_clk new_AGEMA_reg_buffer_13500 ( .C (clk), .D (new_AGEMA_signal_34455), .Q (new_AGEMA_signal_34456) ) ;
    buf_clk new_AGEMA_reg_buffer_13504 ( .C (clk), .D (new_AGEMA_signal_34459), .Q (new_AGEMA_signal_34460) ) ;
    buf_clk new_AGEMA_reg_buffer_13508 ( .C (clk), .D (new_AGEMA_signal_34463), .Q (new_AGEMA_signal_34464) ) ;
    buf_clk new_AGEMA_reg_buffer_13512 ( .C (clk), .D (new_AGEMA_signal_34467), .Q (new_AGEMA_signal_34468) ) ;
    buf_clk new_AGEMA_reg_buffer_13516 ( .C (clk), .D (new_AGEMA_signal_34471), .Q (new_AGEMA_signal_34472) ) ;
    buf_clk new_AGEMA_reg_buffer_13520 ( .C (clk), .D (new_AGEMA_signal_34475), .Q (new_AGEMA_signal_34476) ) ;
    buf_clk new_AGEMA_reg_buffer_13524 ( .C (clk), .D (new_AGEMA_signal_34479), .Q (new_AGEMA_signal_34480) ) ;
    buf_clk new_AGEMA_reg_buffer_13528 ( .C (clk), .D (new_AGEMA_signal_34483), .Q (new_AGEMA_signal_34484) ) ;
    buf_clk new_AGEMA_reg_buffer_13532 ( .C (clk), .D (new_AGEMA_signal_34487), .Q (new_AGEMA_signal_34488) ) ;
    buf_clk new_AGEMA_reg_buffer_13536 ( .C (clk), .D (new_AGEMA_signal_34491), .Q (new_AGEMA_signal_34492) ) ;
    buf_clk new_AGEMA_reg_buffer_13540 ( .C (clk), .D (new_AGEMA_signal_34495), .Q (new_AGEMA_signal_34496) ) ;
    buf_clk new_AGEMA_reg_buffer_13544 ( .C (clk), .D (new_AGEMA_signal_34499), .Q (new_AGEMA_signal_34500) ) ;
    buf_clk new_AGEMA_reg_buffer_13548 ( .C (clk), .D (new_AGEMA_signal_34503), .Q (new_AGEMA_signal_34504) ) ;
    buf_clk new_AGEMA_reg_buffer_13552 ( .C (clk), .D (new_AGEMA_signal_34507), .Q (new_AGEMA_signal_34508) ) ;
    buf_clk new_AGEMA_reg_buffer_13556 ( .C (clk), .D (new_AGEMA_signal_34511), .Q (new_AGEMA_signal_34512) ) ;
    buf_clk new_AGEMA_reg_buffer_13560 ( .C (clk), .D (new_AGEMA_signal_34515), .Q (new_AGEMA_signal_34516) ) ;
    buf_clk new_AGEMA_reg_buffer_13564 ( .C (clk), .D (new_AGEMA_signal_34519), .Q (new_AGEMA_signal_34520) ) ;
    buf_clk new_AGEMA_reg_buffer_13568 ( .C (clk), .D (new_AGEMA_signal_34523), .Q (new_AGEMA_signal_34524) ) ;
    buf_clk new_AGEMA_reg_buffer_13572 ( .C (clk), .D (new_AGEMA_signal_34527), .Q (new_AGEMA_signal_34528) ) ;
    buf_clk new_AGEMA_reg_buffer_13576 ( .C (clk), .D (new_AGEMA_signal_34531), .Q (new_AGEMA_signal_34532) ) ;
    buf_clk new_AGEMA_reg_buffer_13580 ( .C (clk), .D (new_AGEMA_signal_34535), .Q (new_AGEMA_signal_34536) ) ;
    buf_clk new_AGEMA_reg_buffer_13584 ( .C (clk), .D (new_AGEMA_signal_34539), .Q (new_AGEMA_signal_34540) ) ;
    buf_clk new_AGEMA_reg_buffer_13588 ( .C (clk), .D (new_AGEMA_signal_34543), .Q (new_AGEMA_signal_34544) ) ;
    buf_clk new_AGEMA_reg_buffer_13592 ( .C (clk), .D (new_AGEMA_signal_34547), .Q (new_AGEMA_signal_34548) ) ;
    buf_clk new_AGEMA_reg_buffer_13596 ( .C (clk), .D (new_AGEMA_signal_34551), .Q (new_AGEMA_signal_34552) ) ;
    buf_clk new_AGEMA_reg_buffer_13600 ( .C (clk), .D (new_AGEMA_signal_34555), .Q (new_AGEMA_signal_34556) ) ;
    buf_clk new_AGEMA_reg_buffer_13604 ( .C (clk), .D (new_AGEMA_signal_34559), .Q (new_AGEMA_signal_34560) ) ;
    buf_clk new_AGEMA_reg_buffer_13608 ( .C (clk), .D (new_AGEMA_signal_34563), .Q (new_AGEMA_signal_34564) ) ;
    buf_clk new_AGEMA_reg_buffer_13612 ( .C (clk), .D (new_AGEMA_signal_34567), .Q (new_AGEMA_signal_34568) ) ;
    buf_clk new_AGEMA_reg_buffer_13616 ( .C (clk), .D (new_AGEMA_signal_34571), .Q (new_AGEMA_signal_34572) ) ;
    buf_clk new_AGEMA_reg_buffer_13620 ( .C (clk), .D (new_AGEMA_signal_34575), .Q (new_AGEMA_signal_34576) ) ;
    buf_clk new_AGEMA_reg_buffer_13624 ( .C (clk), .D (new_AGEMA_signal_34579), .Q (new_AGEMA_signal_34580) ) ;
    buf_clk new_AGEMA_reg_buffer_13628 ( .C (clk), .D (new_AGEMA_signal_34583), .Q (new_AGEMA_signal_34584) ) ;
    buf_clk new_AGEMA_reg_buffer_13632 ( .C (clk), .D (new_AGEMA_signal_34587), .Q (new_AGEMA_signal_34588) ) ;
    buf_clk new_AGEMA_reg_buffer_13636 ( .C (clk), .D (new_AGEMA_signal_34591), .Q (new_AGEMA_signal_34592) ) ;
    buf_clk new_AGEMA_reg_buffer_13640 ( .C (clk), .D (new_AGEMA_signal_34595), .Q (new_AGEMA_signal_34596) ) ;
    buf_clk new_AGEMA_reg_buffer_13644 ( .C (clk), .D (new_AGEMA_signal_34599), .Q (new_AGEMA_signal_34600) ) ;
    buf_clk new_AGEMA_reg_buffer_13648 ( .C (clk), .D (new_AGEMA_signal_34603), .Q (new_AGEMA_signal_34604) ) ;
    buf_clk new_AGEMA_reg_buffer_13652 ( .C (clk), .D (new_AGEMA_signal_34607), .Q (new_AGEMA_signal_34608) ) ;
    buf_clk new_AGEMA_reg_buffer_13656 ( .C (clk), .D (new_AGEMA_signal_34611), .Q (new_AGEMA_signal_34612) ) ;
    buf_clk new_AGEMA_reg_buffer_13660 ( .C (clk), .D (new_AGEMA_signal_34615), .Q (new_AGEMA_signal_34616) ) ;
    buf_clk new_AGEMA_reg_buffer_13664 ( .C (clk), .D (new_AGEMA_signal_34619), .Q (new_AGEMA_signal_34620) ) ;
    buf_clk new_AGEMA_reg_buffer_13668 ( .C (clk), .D (new_AGEMA_signal_34623), .Q (new_AGEMA_signal_34624) ) ;
    buf_clk new_AGEMA_reg_buffer_13672 ( .C (clk), .D (new_AGEMA_signal_34627), .Q (new_AGEMA_signal_34628) ) ;
    buf_clk new_AGEMA_reg_buffer_13676 ( .C (clk), .D (new_AGEMA_signal_34631), .Q (new_AGEMA_signal_34632) ) ;
    buf_clk new_AGEMA_reg_buffer_13680 ( .C (clk), .D (new_AGEMA_signal_34635), .Q (new_AGEMA_signal_34636) ) ;
    buf_clk new_AGEMA_reg_buffer_13684 ( .C (clk), .D (new_AGEMA_signal_34639), .Q (new_AGEMA_signal_34640) ) ;
    buf_clk new_AGEMA_reg_buffer_13688 ( .C (clk), .D (new_AGEMA_signal_34643), .Q (new_AGEMA_signal_34644) ) ;
    buf_clk new_AGEMA_reg_buffer_13692 ( .C (clk), .D (new_AGEMA_signal_34647), .Q (new_AGEMA_signal_34648) ) ;
    buf_clk new_AGEMA_reg_buffer_13696 ( .C (clk), .D (new_AGEMA_signal_34651), .Q (new_AGEMA_signal_34652) ) ;
    buf_clk new_AGEMA_reg_buffer_13700 ( .C (clk), .D (new_AGEMA_signal_34655), .Q (new_AGEMA_signal_34656) ) ;
    buf_clk new_AGEMA_reg_buffer_13704 ( .C (clk), .D (new_AGEMA_signal_34659), .Q (new_AGEMA_signal_34660) ) ;
    buf_clk new_AGEMA_reg_buffer_13708 ( .C (clk), .D (new_AGEMA_signal_34663), .Q (new_AGEMA_signal_34664) ) ;
    buf_clk new_AGEMA_reg_buffer_13712 ( .C (clk), .D (new_AGEMA_signal_34667), .Q (new_AGEMA_signal_34668) ) ;
    buf_clk new_AGEMA_reg_buffer_13716 ( .C (clk), .D (new_AGEMA_signal_34671), .Q (new_AGEMA_signal_34672) ) ;
    buf_clk new_AGEMA_reg_buffer_13720 ( .C (clk), .D (new_AGEMA_signal_34675), .Q (new_AGEMA_signal_34676) ) ;
    buf_clk new_AGEMA_reg_buffer_13724 ( .C (clk), .D (new_AGEMA_signal_34679), .Q (new_AGEMA_signal_34680) ) ;
    buf_clk new_AGEMA_reg_buffer_13728 ( .C (clk), .D (new_AGEMA_signal_34683), .Q (new_AGEMA_signal_34684) ) ;
    buf_clk new_AGEMA_reg_buffer_13732 ( .C (clk), .D (new_AGEMA_signal_34687), .Q (new_AGEMA_signal_34688) ) ;
    buf_clk new_AGEMA_reg_buffer_13736 ( .C (clk), .D (new_AGEMA_signal_34691), .Q (new_AGEMA_signal_34692) ) ;
    buf_clk new_AGEMA_reg_buffer_13740 ( .C (clk), .D (new_AGEMA_signal_34695), .Q (new_AGEMA_signal_34696) ) ;
    buf_clk new_AGEMA_reg_buffer_13744 ( .C (clk), .D (new_AGEMA_signal_34699), .Q (new_AGEMA_signal_34700) ) ;
    buf_clk new_AGEMA_reg_buffer_13748 ( .C (clk), .D (new_AGEMA_signal_34703), .Q (new_AGEMA_signal_34704) ) ;
    buf_clk new_AGEMA_reg_buffer_13752 ( .C (clk), .D (new_AGEMA_signal_34707), .Q (new_AGEMA_signal_34708) ) ;
    buf_clk new_AGEMA_reg_buffer_13756 ( .C (clk), .D (new_AGEMA_signal_34711), .Q (new_AGEMA_signal_34712) ) ;
    buf_clk new_AGEMA_reg_buffer_13760 ( .C (clk), .D (new_AGEMA_signal_34715), .Q (new_AGEMA_signal_34716) ) ;
    buf_clk new_AGEMA_reg_buffer_13764 ( .C (clk), .D (new_AGEMA_signal_34719), .Q (new_AGEMA_signal_34720) ) ;
    buf_clk new_AGEMA_reg_buffer_13768 ( .C (clk), .D (new_AGEMA_signal_34723), .Q (new_AGEMA_signal_34724) ) ;
    buf_clk new_AGEMA_reg_buffer_13772 ( .C (clk), .D (new_AGEMA_signal_34727), .Q (new_AGEMA_signal_34728) ) ;
    buf_clk new_AGEMA_reg_buffer_13776 ( .C (clk), .D (new_AGEMA_signal_34731), .Q (new_AGEMA_signal_34732) ) ;
    buf_clk new_AGEMA_reg_buffer_13780 ( .C (clk), .D (new_AGEMA_signal_34735), .Q (new_AGEMA_signal_34736) ) ;
    buf_clk new_AGEMA_reg_buffer_13784 ( .C (clk), .D (new_AGEMA_signal_34739), .Q (new_AGEMA_signal_34740) ) ;
    buf_clk new_AGEMA_reg_buffer_13788 ( .C (clk), .D (new_AGEMA_signal_34743), .Q (new_AGEMA_signal_34744) ) ;
    buf_clk new_AGEMA_reg_buffer_13792 ( .C (clk), .D (new_AGEMA_signal_34747), .Q (new_AGEMA_signal_34748) ) ;
    buf_clk new_AGEMA_reg_buffer_13796 ( .C (clk), .D (new_AGEMA_signal_34751), .Q (new_AGEMA_signal_34752) ) ;
    buf_clk new_AGEMA_reg_buffer_13800 ( .C (clk), .D (new_AGEMA_signal_34755), .Q (new_AGEMA_signal_34756) ) ;
    buf_clk new_AGEMA_reg_buffer_13804 ( .C (clk), .D (new_AGEMA_signal_34759), .Q (new_AGEMA_signal_34760) ) ;
    buf_clk new_AGEMA_reg_buffer_13808 ( .C (clk), .D (new_AGEMA_signal_34763), .Q (new_AGEMA_signal_34764) ) ;
    buf_clk new_AGEMA_reg_buffer_13812 ( .C (clk), .D (new_AGEMA_signal_34767), .Q (new_AGEMA_signal_34768) ) ;
    buf_clk new_AGEMA_reg_buffer_13816 ( .C (clk), .D (new_AGEMA_signal_34771), .Q (new_AGEMA_signal_34772) ) ;
    buf_clk new_AGEMA_reg_buffer_13820 ( .C (clk), .D (new_AGEMA_signal_34775), .Q (new_AGEMA_signal_34776) ) ;
    buf_clk new_AGEMA_reg_buffer_13824 ( .C (clk), .D (new_AGEMA_signal_34779), .Q (new_AGEMA_signal_34780) ) ;
    buf_clk new_AGEMA_reg_buffer_13828 ( .C (clk), .D (new_AGEMA_signal_34783), .Q (new_AGEMA_signal_34784) ) ;
    buf_clk new_AGEMA_reg_buffer_13832 ( .C (clk), .D (new_AGEMA_signal_34787), .Q (new_AGEMA_signal_34788) ) ;
    buf_clk new_AGEMA_reg_buffer_13836 ( .C (clk), .D (new_AGEMA_signal_34791), .Q (new_AGEMA_signal_34792) ) ;
    buf_clk new_AGEMA_reg_buffer_13840 ( .C (clk), .D (new_AGEMA_signal_34795), .Q (new_AGEMA_signal_34796) ) ;
    buf_clk new_AGEMA_reg_buffer_13844 ( .C (clk), .D (new_AGEMA_signal_34799), .Q (new_AGEMA_signal_34800) ) ;
    buf_clk new_AGEMA_reg_buffer_13848 ( .C (clk), .D (new_AGEMA_signal_34803), .Q (new_AGEMA_signal_34804) ) ;
    buf_clk new_AGEMA_reg_buffer_13852 ( .C (clk), .D (new_AGEMA_signal_34807), .Q (new_AGEMA_signal_34808) ) ;
    buf_clk new_AGEMA_reg_buffer_13856 ( .C (clk), .D (new_AGEMA_signal_34811), .Q (new_AGEMA_signal_34812) ) ;
    buf_clk new_AGEMA_reg_buffer_13860 ( .C (clk), .D (new_AGEMA_signal_34815), .Q (new_AGEMA_signal_34816) ) ;
    buf_clk new_AGEMA_reg_buffer_13864 ( .C (clk), .D (new_AGEMA_signal_34819), .Q (new_AGEMA_signal_34820) ) ;
    buf_clk new_AGEMA_reg_buffer_13868 ( .C (clk), .D (new_AGEMA_signal_34823), .Q (new_AGEMA_signal_34824) ) ;
    buf_clk new_AGEMA_reg_buffer_13872 ( .C (clk), .D (new_AGEMA_signal_34827), .Q (new_AGEMA_signal_34828) ) ;
    buf_clk new_AGEMA_reg_buffer_13876 ( .C (clk), .D (new_AGEMA_signal_34831), .Q (new_AGEMA_signal_34832) ) ;
    buf_clk new_AGEMA_reg_buffer_13880 ( .C (clk), .D (new_AGEMA_signal_34835), .Q (new_AGEMA_signal_34836) ) ;
    buf_clk new_AGEMA_reg_buffer_13884 ( .C (clk), .D (new_AGEMA_signal_34839), .Q (new_AGEMA_signal_34840) ) ;
    buf_clk new_AGEMA_reg_buffer_13888 ( .C (clk), .D (new_AGEMA_signal_34843), .Q (new_AGEMA_signal_34844) ) ;
    buf_clk new_AGEMA_reg_buffer_13892 ( .C (clk), .D (new_AGEMA_signal_34847), .Q (new_AGEMA_signal_34848) ) ;
    buf_clk new_AGEMA_reg_buffer_13896 ( .C (clk), .D (new_AGEMA_signal_34851), .Q (new_AGEMA_signal_34852) ) ;
    buf_clk new_AGEMA_reg_buffer_13900 ( .C (clk), .D (new_AGEMA_signal_34855), .Q (new_AGEMA_signal_34856) ) ;
    buf_clk new_AGEMA_reg_buffer_13904 ( .C (clk), .D (new_AGEMA_signal_34859), .Q (new_AGEMA_signal_34860) ) ;
    buf_clk new_AGEMA_reg_buffer_13908 ( .C (clk), .D (new_AGEMA_signal_34863), .Q (new_AGEMA_signal_34864) ) ;
    buf_clk new_AGEMA_reg_buffer_13912 ( .C (clk), .D (new_AGEMA_signal_34867), .Q (new_AGEMA_signal_34868) ) ;
    buf_clk new_AGEMA_reg_buffer_13916 ( .C (clk), .D (new_AGEMA_signal_34871), .Q (new_AGEMA_signal_34872) ) ;
    buf_clk new_AGEMA_reg_buffer_13920 ( .C (clk), .D (new_AGEMA_signal_34875), .Q (new_AGEMA_signal_34876) ) ;
    buf_clk new_AGEMA_reg_buffer_13924 ( .C (clk), .D (new_AGEMA_signal_34879), .Q (new_AGEMA_signal_34880) ) ;
    buf_clk new_AGEMA_reg_buffer_13928 ( .C (clk), .D (new_AGEMA_signal_34883), .Q (new_AGEMA_signal_34884) ) ;
    buf_clk new_AGEMA_reg_buffer_13932 ( .C (clk), .D (new_AGEMA_signal_34887), .Q (new_AGEMA_signal_34888) ) ;
    buf_clk new_AGEMA_reg_buffer_13936 ( .C (clk), .D (new_AGEMA_signal_34891), .Q (new_AGEMA_signal_34892) ) ;
    buf_clk new_AGEMA_reg_buffer_13940 ( .C (clk), .D (new_AGEMA_signal_34895), .Q (new_AGEMA_signal_34896) ) ;
    buf_clk new_AGEMA_reg_buffer_13944 ( .C (clk), .D (new_AGEMA_signal_34899), .Q (new_AGEMA_signal_34900) ) ;
    buf_clk new_AGEMA_reg_buffer_13948 ( .C (clk), .D (new_AGEMA_signal_34903), .Q (new_AGEMA_signal_34904) ) ;
    buf_clk new_AGEMA_reg_buffer_13952 ( .C (clk), .D (new_AGEMA_signal_34907), .Q (new_AGEMA_signal_34908) ) ;
    buf_clk new_AGEMA_reg_buffer_13956 ( .C (clk), .D (new_AGEMA_signal_34911), .Q (new_AGEMA_signal_34912) ) ;
    buf_clk new_AGEMA_reg_buffer_13960 ( .C (clk), .D (new_AGEMA_signal_34915), .Q (new_AGEMA_signal_34916) ) ;
    buf_clk new_AGEMA_reg_buffer_13964 ( .C (clk), .D (new_AGEMA_signal_34919), .Q (new_AGEMA_signal_34920) ) ;
    buf_clk new_AGEMA_reg_buffer_13968 ( .C (clk), .D (new_AGEMA_signal_34923), .Q (new_AGEMA_signal_34924) ) ;
    buf_clk new_AGEMA_reg_buffer_13972 ( .C (clk), .D (new_AGEMA_signal_34927), .Q (new_AGEMA_signal_34928) ) ;
    buf_clk new_AGEMA_reg_buffer_13976 ( .C (clk), .D (new_AGEMA_signal_34931), .Q (new_AGEMA_signal_34932) ) ;
    buf_clk new_AGEMA_reg_buffer_13980 ( .C (clk), .D (new_AGEMA_signal_34935), .Q (new_AGEMA_signal_34936) ) ;
    buf_clk new_AGEMA_reg_buffer_13984 ( .C (clk), .D (new_AGEMA_signal_34939), .Q (new_AGEMA_signal_34940) ) ;
    buf_clk new_AGEMA_reg_buffer_13988 ( .C (clk), .D (new_AGEMA_signal_34943), .Q (new_AGEMA_signal_34944) ) ;
    buf_clk new_AGEMA_reg_buffer_13992 ( .C (clk), .D (new_AGEMA_signal_34947), .Q (new_AGEMA_signal_34948) ) ;
    buf_clk new_AGEMA_reg_buffer_13996 ( .C (clk), .D (new_AGEMA_signal_34951), .Q (new_AGEMA_signal_34952) ) ;
    buf_clk new_AGEMA_reg_buffer_14000 ( .C (clk), .D (new_AGEMA_signal_34955), .Q (new_AGEMA_signal_34956) ) ;
    buf_clk new_AGEMA_reg_buffer_14004 ( .C (clk), .D (new_AGEMA_signal_34959), .Q (new_AGEMA_signal_34960) ) ;
    buf_clk new_AGEMA_reg_buffer_14008 ( .C (clk), .D (new_AGEMA_signal_34963), .Q (new_AGEMA_signal_34964) ) ;
    buf_clk new_AGEMA_reg_buffer_14012 ( .C (clk), .D (new_AGEMA_signal_34967), .Q (new_AGEMA_signal_34968) ) ;
    buf_clk new_AGEMA_reg_buffer_14016 ( .C (clk), .D (new_AGEMA_signal_34971), .Q (new_AGEMA_signal_34972) ) ;
    buf_clk new_AGEMA_reg_buffer_14020 ( .C (clk), .D (new_AGEMA_signal_34975), .Q (new_AGEMA_signal_34976) ) ;
    buf_clk new_AGEMA_reg_buffer_14024 ( .C (clk), .D (new_AGEMA_signal_34979), .Q (new_AGEMA_signal_34980) ) ;
    buf_clk new_AGEMA_reg_buffer_14028 ( .C (clk), .D (new_AGEMA_signal_34983), .Q (new_AGEMA_signal_34984) ) ;
    buf_clk new_AGEMA_reg_buffer_14032 ( .C (clk), .D (new_AGEMA_signal_34987), .Q (new_AGEMA_signal_34988) ) ;
    buf_clk new_AGEMA_reg_buffer_14036 ( .C (clk), .D (new_AGEMA_signal_34991), .Q (new_AGEMA_signal_34992) ) ;
    buf_clk new_AGEMA_reg_buffer_14040 ( .C (clk), .D (new_AGEMA_signal_34995), .Q (new_AGEMA_signal_34996) ) ;
    buf_clk new_AGEMA_reg_buffer_14044 ( .C (clk), .D (new_AGEMA_signal_34999), .Q (new_AGEMA_signal_35000) ) ;
    buf_clk new_AGEMA_reg_buffer_14048 ( .C (clk), .D (new_AGEMA_signal_35003), .Q (new_AGEMA_signal_35004) ) ;
    buf_clk new_AGEMA_reg_buffer_14052 ( .C (clk), .D (new_AGEMA_signal_35007), .Q (new_AGEMA_signal_35008) ) ;
    buf_clk new_AGEMA_reg_buffer_14056 ( .C (clk), .D (new_AGEMA_signal_35011), .Q (new_AGEMA_signal_35012) ) ;
    buf_clk new_AGEMA_reg_buffer_14060 ( .C (clk), .D (new_AGEMA_signal_35015), .Q (new_AGEMA_signal_35016) ) ;
    buf_clk new_AGEMA_reg_buffer_14064 ( .C (clk), .D (new_AGEMA_signal_35019), .Q (new_AGEMA_signal_35020) ) ;
    buf_clk new_AGEMA_reg_buffer_14068 ( .C (clk), .D (new_AGEMA_signal_35023), .Q (new_AGEMA_signal_35024) ) ;
    buf_clk new_AGEMA_reg_buffer_14072 ( .C (clk), .D (new_AGEMA_signal_35027), .Q (new_AGEMA_signal_35028) ) ;
    buf_clk new_AGEMA_reg_buffer_14076 ( .C (clk), .D (new_AGEMA_signal_35031), .Q (new_AGEMA_signal_35032) ) ;
    buf_clk new_AGEMA_reg_buffer_14080 ( .C (clk), .D (new_AGEMA_signal_35035), .Q (new_AGEMA_signal_35036) ) ;
    buf_clk new_AGEMA_reg_buffer_14084 ( .C (clk), .D (new_AGEMA_signal_35039), .Q (new_AGEMA_signal_35040) ) ;
    buf_clk new_AGEMA_reg_buffer_14088 ( .C (clk), .D (new_AGEMA_signal_35043), .Q (new_AGEMA_signal_35044) ) ;
    buf_clk new_AGEMA_reg_buffer_14092 ( .C (clk), .D (new_AGEMA_signal_35047), .Q (new_AGEMA_signal_35048) ) ;
    buf_clk new_AGEMA_reg_buffer_14096 ( .C (clk), .D (new_AGEMA_signal_35051), .Q (new_AGEMA_signal_35052) ) ;
    buf_clk new_AGEMA_reg_buffer_14100 ( .C (clk), .D (new_AGEMA_signal_35055), .Q (new_AGEMA_signal_35056) ) ;
    buf_clk new_AGEMA_reg_buffer_14104 ( .C (clk), .D (new_AGEMA_signal_35059), .Q (new_AGEMA_signal_35060) ) ;
    buf_clk new_AGEMA_reg_buffer_14108 ( .C (clk), .D (new_AGEMA_signal_35063), .Q (new_AGEMA_signal_35064) ) ;
    buf_clk new_AGEMA_reg_buffer_14112 ( .C (clk), .D (new_AGEMA_signal_35067), .Q (new_AGEMA_signal_35068) ) ;
    buf_clk new_AGEMA_reg_buffer_14116 ( .C (clk), .D (new_AGEMA_signal_35071), .Q (new_AGEMA_signal_35072) ) ;
    buf_clk new_AGEMA_reg_buffer_14120 ( .C (clk), .D (new_AGEMA_signal_35075), .Q (new_AGEMA_signal_35076) ) ;
    buf_clk new_AGEMA_reg_buffer_14124 ( .C (clk), .D (new_AGEMA_signal_35079), .Q (new_AGEMA_signal_35080) ) ;
    buf_clk new_AGEMA_reg_buffer_14128 ( .C (clk), .D (new_AGEMA_signal_35083), .Q (new_AGEMA_signal_35084) ) ;
    buf_clk new_AGEMA_reg_buffer_14132 ( .C (clk), .D (new_AGEMA_signal_35087), .Q (new_AGEMA_signal_35088) ) ;
    buf_clk new_AGEMA_reg_buffer_14136 ( .C (clk), .D (new_AGEMA_signal_35091), .Q (new_AGEMA_signal_35092) ) ;
    buf_clk new_AGEMA_reg_buffer_14140 ( .C (clk), .D (new_AGEMA_signal_35095), .Q (new_AGEMA_signal_35096) ) ;
    buf_clk new_AGEMA_reg_buffer_14144 ( .C (clk), .D (new_AGEMA_signal_35099), .Q (new_AGEMA_signal_35100) ) ;
    buf_clk new_AGEMA_reg_buffer_14148 ( .C (clk), .D (new_AGEMA_signal_35103), .Q (new_AGEMA_signal_35104) ) ;
    buf_clk new_AGEMA_reg_buffer_14152 ( .C (clk), .D (new_AGEMA_signal_35107), .Q (new_AGEMA_signal_35108) ) ;
    buf_clk new_AGEMA_reg_buffer_14156 ( .C (clk), .D (new_AGEMA_signal_35111), .Q (new_AGEMA_signal_35112) ) ;
    buf_clk new_AGEMA_reg_buffer_14160 ( .C (clk), .D (new_AGEMA_signal_35115), .Q (new_AGEMA_signal_35116) ) ;
    buf_clk new_AGEMA_reg_buffer_14164 ( .C (clk), .D (new_AGEMA_signal_35119), .Q (new_AGEMA_signal_35120) ) ;
    buf_clk new_AGEMA_reg_buffer_14168 ( .C (clk), .D (new_AGEMA_signal_35123), .Q (new_AGEMA_signal_35124) ) ;
    buf_clk new_AGEMA_reg_buffer_14172 ( .C (clk), .D (new_AGEMA_signal_35127), .Q (new_AGEMA_signal_35128) ) ;
    buf_clk new_AGEMA_reg_buffer_14176 ( .C (clk), .D (new_AGEMA_signal_35131), .Q (new_AGEMA_signal_35132) ) ;
    buf_clk new_AGEMA_reg_buffer_14180 ( .C (clk), .D (new_AGEMA_signal_35135), .Q (new_AGEMA_signal_35136) ) ;
    buf_clk new_AGEMA_reg_buffer_14184 ( .C (clk), .D (new_AGEMA_signal_35139), .Q (new_AGEMA_signal_35140) ) ;
    buf_clk new_AGEMA_reg_buffer_14188 ( .C (clk), .D (new_AGEMA_signal_35143), .Q (new_AGEMA_signal_35144) ) ;
    buf_clk new_AGEMA_reg_buffer_14192 ( .C (clk), .D (new_AGEMA_signal_35147), .Q (new_AGEMA_signal_35148) ) ;
    buf_clk new_AGEMA_reg_buffer_14196 ( .C (clk), .D (new_AGEMA_signal_35151), .Q (new_AGEMA_signal_35152) ) ;
    buf_clk new_AGEMA_reg_buffer_14200 ( .C (clk), .D (new_AGEMA_signal_35155), .Q (new_AGEMA_signal_35156) ) ;
    buf_clk new_AGEMA_reg_buffer_14204 ( .C (clk), .D (new_AGEMA_signal_35159), .Q (new_AGEMA_signal_35160) ) ;
    buf_clk new_AGEMA_reg_buffer_14208 ( .C (clk), .D (new_AGEMA_signal_35163), .Q (new_AGEMA_signal_35164) ) ;
    buf_clk new_AGEMA_reg_buffer_14212 ( .C (clk), .D (new_AGEMA_signal_35167), .Q (new_AGEMA_signal_35168) ) ;
    buf_clk new_AGEMA_reg_buffer_14216 ( .C (clk), .D (new_AGEMA_signal_35171), .Q (new_AGEMA_signal_35172) ) ;
    buf_clk new_AGEMA_reg_buffer_14220 ( .C (clk), .D (new_AGEMA_signal_35175), .Q (new_AGEMA_signal_35176) ) ;
    buf_clk new_AGEMA_reg_buffer_14224 ( .C (clk), .D (new_AGEMA_signal_35179), .Q (new_AGEMA_signal_35180) ) ;
    buf_clk new_AGEMA_reg_buffer_14228 ( .C (clk), .D (new_AGEMA_signal_35183), .Q (new_AGEMA_signal_35184) ) ;
    buf_clk new_AGEMA_reg_buffer_14232 ( .C (clk), .D (new_AGEMA_signal_35187), .Q (new_AGEMA_signal_35188) ) ;
    buf_clk new_AGEMA_reg_buffer_14236 ( .C (clk), .D (new_AGEMA_signal_35191), .Q (new_AGEMA_signal_35192) ) ;
    buf_clk new_AGEMA_reg_buffer_14240 ( .C (clk), .D (new_AGEMA_signal_35195), .Q (new_AGEMA_signal_35196) ) ;
    buf_clk new_AGEMA_reg_buffer_14244 ( .C (clk), .D (new_AGEMA_signal_35199), .Q (new_AGEMA_signal_35200) ) ;
    buf_clk new_AGEMA_reg_buffer_14248 ( .C (clk), .D (new_AGEMA_signal_35203), .Q (new_AGEMA_signal_35204) ) ;
    buf_clk new_AGEMA_reg_buffer_14252 ( .C (clk), .D (new_AGEMA_signal_35207), .Q (new_AGEMA_signal_35208) ) ;
    buf_clk new_AGEMA_reg_buffer_14256 ( .C (clk), .D (new_AGEMA_signal_35211), .Q (new_AGEMA_signal_35212) ) ;
    buf_clk new_AGEMA_reg_buffer_14260 ( .C (clk), .D (new_AGEMA_signal_35215), .Q (new_AGEMA_signal_35216) ) ;
    buf_clk new_AGEMA_reg_buffer_14264 ( .C (clk), .D (new_AGEMA_signal_35219), .Q (new_AGEMA_signal_35220) ) ;
    buf_clk new_AGEMA_reg_buffer_14268 ( .C (clk), .D (new_AGEMA_signal_35223), .Q (new_AGEMA_signal_35224) ) ;
    buf_clk new_AGEMA_reg_buffer_14272 ( .C (clk), .D (new_AGEMA_signal_35227), .Q (new_AGEMA_signal_35228) ) ;
    buf_clk new_AGEMA_reg_buffer_14276 ( .C (clk), .D (new_AGEMA_signal_35231), .Q (new_AGEMA_signal_35232) ) ;
    buf_clk new_AGEMA_reg_buffer_14280 ( .C (clk), .D (new_AGEMA_signal_35235), .Q (new_AGEMA_signal_35236) ) ;
    buf_clk new_AGEMA_reg_buffer_14284 ( .C (clk), .D (new_AGEMA_signal_35239), .Q (new_AGEMA_signal_35240) ) ;
    buf_clk new_AGEMA_reg_buffer_14288 ( .C (clk), .D (new_AGEMA_signal_35243), .Q (new_AGEMA_signal_35244) ) ;
    buf_clk new_AGEMA_reg_buffer_14292 ( .C (clk), .D (new_AGEMA_signal_35247), .Q (new_AGEMA_signal_35248) ) ;
    buf_clk new_AGEMA_reg_buffer_14296 ( .C (clk), .D (new_AGEMA_signal_35251), .Q (new_AGEMA_signal_35252) ) ;
    buf_clk new_AGEMA_reg_buffer_14300 ( .C (clk), .D (new_AGEMA_signal_35255), .Q (new_AGEMA_signal_35256) ) ;
    buf_clk new_AGEMA_reg_buffer_14304 ( .C (clk), .D (new_AGEMA_signal_35259), .Q (new_AGEMA_signal_35260) ) ;
    buf_clk new_AGEMA_reg_buffer_14308 ( .C (clk), .D (new_AGEMA_signal_35263), .Q (new_AGEMA_signal_35264) ) ;
    buf_clk new_AGEMA_reg_buffer_14312 ( .C (clk), .D (new_AGEMA_signal_35267), .Q (new_AGEMA_signal_35268) ) ;
    buf_clk new_AGEMA_reg_buffer_14316 ( .C (clk), .D (new_AGEMA_signal_35271), .Q (new_AGEMA_signal_35272) ) ;
    buf_clk new_AGEMA_reg_buffer_14320 ( .C (clk), .D (new_AGEMA_signal_35275), .Q (new_AGEMA_signal_35276) ) ;
    buf_clk new_AGEMA_reg_buffer_14324 ( .C (clk), .D (new_AGEMA_signal_35279), .Q (new_AGEMA_signal_35280) ) ;
    buf_clk new_AGEMA_reg_buffer_14328 ( .C (clk), .D (new_AGEMA_signal_35283), .Q (new_AGEMA_signal_35284) ) ;
    buf_clk new_AGEMA_reg_buffer_14332 ( .C (clk), .D (new_AGEMA_signal_35287), .Q (new_AGEMA_signal_35288) ) ;
    buf_clk new_AGEMA_reg_buffer_14336 ( .C (clk), .D (new_AGEMA_signal_35291), .Q (new_AGEMA_signal_35292) ) ;
    buf_clk new_AGEMA_reg_buffer_14340 ( .C (clk), .D (new_AGEMA_signal_35295), .Q (new_AGEMA_signal_35296) ) ;
    buf_clk new_AGEMA_reg_buffer_14344 ( .C (clk), .D (new_AGEMA_signal_35299), .Q (new_AGEMA_signal_35300) ) ;
    buf_clk new_AGEMA_reg_buffer_14348 ( .C (clk), .D (new_AGEMA_signal_35303), .Q (new_AGEMA_signal_35304) ) ;
    buf_clk new_AGEMA_reg_buffer_14352 ( .C (clk), .D (new_AGEMA_signal_35307), .Q (new_AGEMA_signal_35308) ) ;
    buf_clk new_AGEMA_reg_buffer_14356 ( .C (clk), .D (new_AGEMA_signal_35311), .Q (new_AGEMA_signal_35312) ) ;
    buf_clk new_AGEMA_reg_buffer_14360 ( .C (clk), .D (new_AGEMA_signal_35315), .Q (new_AGEMA_signal_35316) ) ;
    buf_clk new_AGEMA_reg_buffer_14364 ( .C (clk), .D (new_AGEMA_signal_35319), .Q (new_AGEMA_signal_35320) ) ;
    buf_clk new_AGEMA_reg_buffer_14368 ( .C (clk), .D (new_AGEMA_signal_35323), .Q (new_AGEMA_signal_35324) ) ;
    buf_clk new_AGEMA_reg_buffer_14372 ( .C (clk), .D (new_AGEMA_signal_35327), .Q (new_AGEMA_signal_35328) ) ;
    buf_clk new_AGEMA_reg_buffer_14376 ( .C (clk), .D (new_AGEMA_signal_35331), .Q (new_AGEMA_signal_35332) ) ;
    buf_clk new_AGEMA_reg_buffer_14380 ( .C (clk), .D (new_AGEMA_signal_35335), .Q (new_AGEMA_signal_35336) ) ;
    buf_clk new_AGEMA_reg_buffer_14384 ( .C (clk), .D (new_AGEMA_signal_35339), .Q (new_AGEMA_signal_35340) ) ;
    buf_clk new_AGEMA_reg_buffer_14388 ( .C (clk), .D (new_AGEMA_signal_35343), .Q (new_AGEMA_signal_35344) ) ;
    buf_clk new_AGEMA_reg_buffer_14392 ( .C (clk), .D (new_AGEMA_signal_35347), .Q (new_AGEMA_signal_35348) ) ;
    buf_clk new_AGEMA_reg_buffer_14396 ( .C (clk), .D (new_AGEMA_signal_35351), .Q (new_AGEMA_signal_35352) ) ;
    buf_clk new_AGEMA_reg_buffer_14400 ( .C (clk), .D (new_AGEMA_signal_35355), .Q (new_AGEMA_signal_35356) ) ;
    buf_clk new_AGEMA_reg_buffer_14404 ( .C (clk), .D (new_AGEMA_signal_35359), .Q (new_AGEMA_signal_35360) ) ;
    buf_clk new_AGEMA_reg_buffer_14408 ( .C (clk), .D (new_AGEMA_signal_35363), .Q (new_AGEMA_signal_35364) ) ;
    buf_clk new_AGEMA_reg_buffer_14412 ( .C (clk), .D (new_AGEMA_signal_35367), .Q (new_AGEMA_signal_35368) ) ;
    buf_clk new_AGEMA_reg_buffer_14416 ( .C (clk), .D (new_AGEMA_signal_35371), .Q (new_AGEMA_signal_35372) ) ;
    buf_clk new_AGEMA_reg_buffer_14420 ( .C (clk), .D (new_AGEMA_signal_35375), .Q (new_AGEMA_signal_35376) ) ;
    buf_clk new_AGEMA_reg_buffer_14424 ( .C (clk), .D (new_AGEMA_signal_35379), .Q (new_AGEMA_signal_35380) ) ;
    buf_clk new_AGEMA_reg_buffer_14428 ( .C (clk), .D (new_AGEMA_signal_35383), .Q (new_AGEMA_signal_35384) ) ;
    buf_clk new_AGEMA_reg_buffer_14432 ( .C (clk), .D (new_AGEMA_signal_35387), .Q (new_AGEMA_signal_35388) ) ;
    buf_clk new_AGEMA_reg_buffer_14436 ( .C (clk), .D (new_AGEMA_signal_35391), .Q (new_AGEMA_signal_35392) ) ;
    buf_clk new_AGEMA_reg_buffer_14440 ( .C (clk), .D (new_AGEMA_signal_35395), .Q (new_AGEMA_signal_35396) ) ;
    buf_clk new_AGEMA_reg_buffer_14444 ( .C (clk), .D (new_AGEMA_signal_35399), .Q (new_AGEMA_signal_35400) ) ;
    buf_clk new_AGEMA_reg_buffer_14448 ( .C (clk), .D (new_AGEMA_signal_35403), .Q (new_AGEMA_signal_35404) ) ;
    buf_clk new_AGEMA_reg_buffer_14452 ( .C (clk), .D (new_AGEMA_signal_35407), .Q (new_AGEMA_signal_35408) ) ;
    buf_clk new_AGEMA_reg_buffer_14456 ( .C (clk), .D (new_AGEMA_signal_35411), .Q (new_AGEMA_signal_35412) ) ;
    buf_clk new_AGEMA_reg_buffer_14460 ( .C (clk), .D (new_AGEMA_signal_35415), .Q (new_AGEMA_signal_35416) ) ;
    buf_clk new_AGEMA_reg_buffer_14464 ( .C (clk), .D (new_AGEMA_signal_35419), .Q (new_AGEMA_signal_35420) ) ;
    buf_clk new_AGEMA_reg_buffer_14468 ( .C (clk), .D (new_AGEMA_signal_35423), .Q (new_AGEMA_signal_35424) ) ;
    buf_clk new_AGEMA_reg_buffer_14472 ( .C (clk), .D (new_AGEMA_signal_35427), .Q (new_AGEMA_signal_35428) ) ;
    buf_clk new_AGEMA_reg_buffer_14476 ( .C (clk), .D (new_AGEMA_signal_35431), .Q (new_AGEMA_signal_35432) ) ;
    buf_clk new_AGEMA_reg_buffer_14480 ( .C (clk), .D (new_AGEMA_signal_35435), .Q (new_AGEMA_signal_35436) ) ;
    buf_clk new_AGEMA_reg_buffer_14484 ( .C (clk), .D (new_AGEMA_signal_35439), .Q (new_AGEMA_signal_35440) ) ;
    buf_clk new_AGEMA_reg_buffer_14488 ( .C (clk), .D (new_AGEMA_signal_35443), .Q (new_AGEMA_signal_35444) ) ;
    buf_clk new_AGEMA_reg_buffer_14492 ( .C (clk), .D (new_AGEMA_signal_35447), .Q (new_AGEMA_signal_35448) ) ;
    buf_clk new_AGEMA_reg_buffer_14496 ( .C (clk), .D (new_AGEMA_signal_35451), .Q (new_AGEMA_signal_35452) ) ;
    buf_clk new_AGEMA_reg_buffer_14500 ( .C (clk), .D (new_AGEMA_signal_35455), .Q (new_AGEMA_signal_35456) ) ;
    buf_clk new_AGEMA_reg_buffer_14504 ( .C (clk), .D (new_AGEMA_signal_35459), .Q (new_AGEMA_signal_35460) ) ;
    buf_clk new_AGEMA_reg_buffer_14508 ( .C (clk), .D (new_AGEMA_signal_35463), .Q (new_AGEMA_signal_35464) ) ;
    buf_clk new_AGEMA_reg_buffer_14512 ( .C (clk), .D (new_AGEMA_signal_35467), .Q (new_AGEMA_signal_35468) ) ;
    buf_clk new_AGEMA_reg_buffer_14516 ( .C (clk), .D (new_AGEMA_signal_35471), .Q (new_AGEMA_signal_35472) ) ;
    buf_clk new_AGEMA_reg_buffer_14520 ( .C (clk), .D (new_AGEMA_signal_35475), .Q (new_AGEMA_signal_35476) ) ;
    buf_clk new_AGEMA_reg_buffer_14524 ( .C (clk), .D (new_AGEMA_signal_35479), .Q (new_AGEMA_signal_35480) ) ;
    buf_clk new_AGEMA_reg_buffer_14528 ( .C (clk), .D (new_AGEMA_signal_35483), .Q (new_AGEMA_signal_35484) ) ;
    buf_clk new_AGEMA_reg_buffer_14532 ( .C (clk), .D (new_AGEMA_signal_35487), .Q (new_AGEMA_signal_35488) ) ;
    buf_clk new_AGEMA_reg_buffer_14536 ( .C (clk), .D (new_AGEMA_signal_35491), .Q (new_AGEMA_signal_35492) ) ;
    buf_clk new_AGEMA_reg_buffer_14540 ( .C (clk), .D (new_AGEMA_signal_35495), .Q (new_AGEMA_signal_35496) ) ;
    buf_clk new_AGEMA_reg_buffer_14544 ( .C (clk), .D (new_AGEMA_signal_35499), .Q (new_AGEMA_signal_35500) ) ;
    buf_clk new_AGEMA_reg_buffer_14548 ( .C (clk), .D (new_AGEMA_signal_35503), .Q (new_AGEMA_signal_35504) ) ;
    buf_clk new_AGEMA_reg_buffer_14552 ( .C (clk), .D (new_AGEMA_signal_35507), .Q (new_AGEMA_signal_35508) ) ;
    buf_clk new_AGEMA_reg_buffer_14556 ( .C (clk), .D (new_AGEMA_signal_35511), .Q (new_AGEMA_signal_35512) ) ;
    buf_clk new_AGEMA_reg_buffer_14560 ( .C (clk), .D (new_AGEMA_signal_35515), .Q (new_AGEMA_signal_35516) ) ;
    buf_clk new_AGEMA_reg_buffer_14564 ( .C (clk), .D (new_AGEMA_signal_35519), .Q (new_AGEMA_signal_35520) ) ;
    buf_clk new_AGEMA_reg_buffer_14568 ( .C (clk), .D (new_AGEMA_signal_35523), .Q (new_AGEMA_signal_35524) ) ;
    buf_clk new_AGEMA_reg_buffer_14572 ( .C (clk), .D (new_AGEMA_signal_35527), .Q (new_AGEMA_signal_35528) ) ;
    buf_clk new_AGEMA_reg_buffer_14576 ( .C (clk), .D (new_AGEMA_signal_35531), .Q (new_AGEMA_signal_35532) ) ;
    buf_clk new_AGEMA_reg_buffer_14580 ( .C (clk), .D (new_AGEMA_signal_35535), .Q (new_AGEMA_signal_35536) ) ;
    buf_clk new_AGEMA_reg_buffer_14584 ( .C (clk), .D (new_AGEMA_signal_35539), .Q (new_AGEMA_signal_35540) ) ;
    buf_clk new_AGEMA_reg_buffer_14588 ( .C (clk), .D (new_AGEMA_signal_35543), .Q (new_AGEMA_signal_35544) ) ;
    buf_clk new_AGEMA_reg_buffer_14592 ( .C (clk), .D (new_AGEMA_signal_35547), .Q (new_AGEMA_signal_35548) ) ;
    buf_clk new_AGEMA_reg_buffer_14596 ( .C (clk), .D (new_AGEMA_signal_35551), .Q (new_AGEMA_signal_35552) ) ;
    buf_clk new_AGEMA_reg_buffer_14600 ( .C (clk), .D (new_AGEMA_signal_35555), .Q (new_AGEMA_signal_35556) ) ;
    buf_clk new_AGEMA_reg_buffer_14604 ( .C (clk), .D (new_AGEMA_signal_35559), .Q (new_AGEMA_signal_35560) ) ;
    buf_clk new_AGEMA_reg_buffer_14608 ( .C (clk), .D (new_AGEMA_signal_35563), .Q (new_AGEMA_signal_35564) ) ;
    buf_clk new_AGEMA_reg_buffer_14612 ( .C (clk), .D (new_AGEMA_signal_35567), .Q (new_AGEMA_signal_35568) ) ;
    buf_clk new_AGEMA_reg_buffer_14616 ( .C (clk), .D (new_AGEMA_signal_35571), .Q (new_AGEMA_signal_35572) ) ;
    buf_clk new_AGEMA_reg_buffer_14620 ( .C (clk), .D (new_AGEMA_signal_35575), .Q (new_AGEMA_signal_35576) ) ;
    buf_clk new_AGEMA_reg_buffer_14624 ( .C (clk), .D (new_AGEMA_signal_35579), .Q (new_AGEMA_signal_35580) ) ;
    buf_clk new_AGEMA_reg_buffer_14628 ( .C (clk), .D (new_AGEMA_signal_35583), .Q (new_AGEMA_signal_35584) ) ;
    buf_clk new_AGEMA_reg_buffer_14632 ( .C (clk), .D (new_AGEMA_signal_35587), .Q (new_AGEMA_signal_35588) ) ;
    buf_clk new_AGEMA_reg_buffer_14636 ( .C (clk), .D (new_AGEMA_signal_35591), .Q (new_AGEMA_signal_35592) ) ;
    buf_clk new_AGEMA_reg_buffer_14640 ( .C (clk), .D (new_AGEMA_signal_35595), .Q (new_AGEMA_signal_35596) ) ;
    buf_clk new_AGEMA_reg_buffer_14644 ( .C (clk), .D (new_AGEMA_signal_35599), .Q (new_AGEMA_signal_35600) ) ;
    buf_clk new_AGEMA_reg_buffer_14648 ( .C (clk), .D (new_AGEMA_signal_35603), .Q (new_AGEMA_signal_35604) ) ;
    buf_clk new_AGEMA_reg_buffer_14652 ( .C (clk), .D (new_AGEMA_signal_35607), .Q (new_AGEMA_signal_35608) ) ;
    buf_clk new_AGEMA_reg_buffer_14656 ( .C (clk), .D (new_AGEMA_signal_35611), .Q (new_AGEMA_signal_35612) ) ;
    buf_clk new_AGEMA_reg_buffer_14660 ( .C (clk), .D (new_AGEMA_signal_35615), .Q (new_AGEMA_signal_35616) ) ;
    buf_clk new_AGEMA_reg_buffer_14664 ( .C (clk), .D (new_AGEMA_signal_35619), .Q (new_AGEMA_signal_35620) ) ;
    buf_clk new_AGEMA_reg_buffer_14668 ( .C (clk), .D (new_AGEMA_signal_35623), .Q (new_AGEMA_signal_35624) ) ;
    buf_clk new_AGEMA_reg_buffer_14672 ( .C (clk), .D (new_AGEMA_signal_35627), .Q (new_AGEMA_signal_35628) ) ;
    buf_clk new_AGEMA_reg_buffer_14676 ( .C (clk), .D (new_AGEMA_signal_35631), .Q (new_AGEMA_signal_35632) ) ;
    buf_clk new_AGEMA_reg_buffer_14680 ( .C (clk), .D (new_AGEMA_signal_35635), .Q (new_AGEMA_signal_35636) ) ;
    buf_clk new_AGEMA_reg_buffer_14684 ( .C (clk), .D (new_AGEMA_signal_35639), .Q (new_AGEMA_signal_35640) ) ;
    buf_clk new_AGEMA_reg_buffer_14688 ( .C (clk), .D (new_AGEMA_signal_35643), .Q (new_AGEMA_signal_35644) ) ;
    buf_clk new_AGEMA_reg_buffer_14692 ( .C (clk), .D (new_AGEMA_signal_35647), .Q (new_AGEMA_signal_35648) ) ;
    buf_clk new_AGEMA_reg_buffer_14696 ( .C (clk), .D (new_AGEMA_signal_35651), .Q (new_AGEMA_signal_35652) ) ;
    buf_clk new_AGEMA_reg_buffer_14700 ( .C (clk), .D (new_AGEMA_signal_35655), .Q (new_AGEMA_signal_35656) ) ;
    buf_clk new_AGEMA_reg_buffer_14704 ( .C (clk), .D (new_AGEMA_signal_35659), .Q (new_AGEMA_signal_35660) ) ;
    buf_clk new_AGEMA_reg_buffer_14708 ( .C (clk), .D (new_AGEMA_signal_35663), .Q (new_AGEMA_signal_35664) ) ;
    buf_clk new_AGEMA_reg_buffer_14712 ( .C (clk), .D (new_AGEMA_signal_35667), .Q (new_AGEMA_signal_35668) ) ;
    buf_clk new_AGEMA_reg_buffer_14716 ( .C (clk), .D (new_AGEMA_signal_35671), .Q (new_AGEMA_signal_35672) ) ;
    buf_clk new_AGEMA_reg_buffer_14720 ( .C (clk), .D (new_AGEMA_signal_35675), .Q (new_AGEMA_signal_35676) ) ;
    buf_clk new_AGEMA_reg_buffer_14724 ( .C (clk), .D (new_AGEMA_signal_35679), .Q (new_AGEMA_signal_35680) ) ;
    buf_clk new_AGEMA_reg_buffer_14728 ( .C (clk), .D (new_AGEMA_signal_35683), .Q (new_AGEMA_signal_35684) ) ;
    buf_clk new_AGEMA_reg_buffer_14732 ( .C (clk), .D (new_AGEMA_signal_35687), .Q (new_AGEMA_signal_35688) ) ;
    buf_clk new_AGEMA_reg_buffer_14736 ( .C (clk), .D (new_AGEMA_signal_35691), .Q (new_AGEMA_signal_35692) ) ;
    buf_clk new_AGEMA_reg_buffer_14740 ( .C (clk), .D (new_AGEMA_signal_35695), .Q (new_AGEMA_signal_35696) ) ;
    buf_clk new_AGEMA_reg_buffer_14744 ( .C (clk), .D (new_AGEMA_signal_35699), .Q (new_AGEMA_signal_35700) ) ;
    buf_clk new_AGEMA_reg_buffer_14748 ( .C (clk), .D (new_AGEMA_signal_35703), .Q (new_AGEMA_signal_35704) ) ;
    buf_clk new_AGEMA_reg_buffer_14752 ( .C (clk), .D (new_AGEMA_signal_35707), .Q (new_AGEMA_signal_35708) ) ;
    buf_clk new_AGEMA_reg_buffer_14756 ( .C (clk), .D (new_AGEMA_signal_35711), .Q (new_AGEMA_signal_35712) ) ;
    buf_clk new_AGEMA_reg_buffer_14760 ( .C (clk), .D (new_AGEMA_signal_35715), .Q (new_AGEMA_signal_35716) ) ;
    buf_clk new_AGEMA_reg_buffer_14764 ( .C (clk), .D (new_AGEMA_signal_35719), .Q (new_AGEMA_signal_35720) ) ;
    buf_clk new_AGEMA_reg_buffer_14768 ( .C (clk), .D (new_AGEMA_signal_35723), .Q (new_AGEMA_signal_35724) ) ;
    buf_clk new_AGEMA_reg_buffer_14772 ( .C (clk), .D (new_AGEMA_signal_35727), .Q (new_AGEMA_signal_35728) ) ;
    buf_clk new_AGEMA_reg_buffer_14776 ( .C (clk), .D (new_AGEMA_signal_35731), .Q (new_AGEMA_signal_35732) ) ;
    buf_clk new_AGEMA_reg_buffer_14780 ( .C (clk), .D (new_AGEMA_signal_35735), .Q (new_AGEMA_signal_35736) ) ;
    buf_clk new_AGEMA_reg_buffer_14784 ( .C (clk), .D (new_AGEMA_signal_35739), .Q (new_AGEMA_signal_35740) ) ;
    buf_clk new_AGEMA_reg_buffer_14788 ( .C (clk), .D (new_AGEMA_signal_35743), .Q (new_AGEMA_signal_35744) ) ;
    buf_clk new_AGEMA_reg_buffer_14792 ( .C (clk), .D (new_AGEMA_signal_35747), .Q (new_AGEMA_signal_35748) ) ;
    buf_clk new_AGEMA_reg_buffer_14796 ( .C (clk), .D (new_AGEMA_signal_35751), .Q (new_AGEMA_signal_35752) ) ;
    buf_clk new_AGEMA_reg_buffer_14800 ( .C (clk), .D (new_AGEMA_signal_35755), .Q (new_AGEMA_signal_35756) ) ;
    buf_clk new_AGEMA_reg_buffer_14804 ( .C (clk), .D (new_AGEMA_signal_35759), .Q (new_AGEMA_signal_35760) ) ;
    buf_clk new_AGEMA_reg_buffer_14808 ( .C (clk), .D (new_AGEMA_signal_35763), .Q (new_AGEMA_signal_35764) ) ;
    buf_clk new_AGEMA_reg_buffer_14812 ( .C (clk), .D (new_AGEMA_signal_35767), .Q (new_AGEMA_signal_35768) ) ;
    buf_clk new_AGEMA_reg_buffer_14816 ( .C (clk), .D (new_AGEMA_signal_35771), .Q (new_AGEMA_signal_35772) ) ;
    buf_clk new_AGEMA_reg_buffer_14820 ( .C (clk), .D (new_AGEMA_signal_35775), .Q (new_AGEMA_signal_35776) ) ;
    buf_clk new_AGEMA_reg_buffer_14824 ( .C (clk), .D (new_AGEMA_signal_35779), .Q (new_AGEMA_signal_35780) ) ;
    buf_clk new_AGEMA_reg_buffer_14828 ( .C (clk), .D (new_AGEMA_signal_35783), .Q (new_AGEMA_signal_35784) ) ;
    buf_clk new_AGEMA_reg_buffer_14832 ( .C (clk), .D (new_AGEMA_signal_35787), .Q (new_AGEMA_signal_35788) ) ;
    buf_clk new_AGEMA_reg_buffer_15652 ( .C (clk), .D (new_AGEMA_signal_36607), .Q (new_AGEMA_signal_36608) ) ;
    buf_clk new_AGEMA_reg_buffer_15656 ( .C (clk), .D (new_AGEMA_signal_36611), .Q (new_AGEMA_signal_36612) ) ;
    buf_clk new_AGEMA_reg_buffer_15660 ( .C (clk), .D (new_AGEMA_signal_36615), .Q (new_AGEMA_signal_36616) ) ;
    buf_clk new_AGEMA_reg_buffer_15664 ( .C (clk), .D (new_AGEMA_signal_36619), .Q (new_AGEMA_signal_36620) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16200, new_AGEMA_signal_16199, new_AGEMA_signal_16198, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16722, new_AGEMA_signal_16721, new_AGEMA_signal_16720, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, RoundInput[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16206, new_AGEMA_signal_16205, new_AGEMA_signal_16204, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16728, new_AGEMA_signal_16727, new_AGEMA_signal_16726, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundInput[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16734, new_AGEMA_signal_16733, new_AGEMA_signal_16732, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16212, new_AGEMA_signal_16211, new_AGEMA_signal_16210, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, RoundInput[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16218, new_AGEMA_signal_16217, new_AGEMA_signal_16216, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, RoundInput[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16224, new_AGEMA_signal_16223, new_AGEMA_signal_16222, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, RoundInput[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16230, new_AGEMA_signal_16229, new_AGEMA_signal_16228, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, RoundInput[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16740, new_AGEMA_signal_16739, new_AGEMA_signal_16738, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundInput[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16236, new_AGEMA_signal_16235, new_AGEMA_signal_16234, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, RoundInput[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16746, new_AGEMA_signal_16745, new_AGEMA_signal_16744, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16752, new_AGEMA_signal_16751, new_AGEMA_signal_16750, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, RoundInput[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16242, new_AGEMA_signal_16241, new_AGEMA_signal_16240, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16248, new_AGEMA_signal_16247, new_AGEMA_signal_16246, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, RoundInput[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16254, new_AGEMA_signal_16253, new_AGEMA_signal_16252, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16260, new_AGEMA_signal_16259, new_AGEMA_signal_16258, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, RoundInput[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16758, new_AGEMA_signal_16757, new_AGEMA_signal_16756, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16266, new_AGEMA_signal_16265, new_AGEMA_signal_16264, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, RoundInput[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16764, new_AGEMA_signal_16763, new_AGEMA_signal_16762, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16770, new_AGEMA_signal_16769, new_AGEMA_signal_16768, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16272, new_AGEMA_signal_16271, new_AGEMA_signal_16270, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, RoundInput[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16278, new_AGEMA_signal_16277, new_AGEMA_signal_16276, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16284, new_AGEMA_signal_16283, new_AGEMA_signal_16282, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, RoundInput[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16290, new_AGEMA_signal_16289, new_AGEMA_signal_16288, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16776, new_AGEMA_signal_16775, new_AGEMA_signal_16774, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, RoundInput[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16296, new_AGEMA_signal_16295, new_AGEMA_signal_16294, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16782, new_AGEMA_signal_16781, new_AGEMA_signal_16780, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, RoundInput[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16788, new_AGEMA_signal_16787, new_AGEMA_signal_16786, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16302, new_AGEMA_signal_16301, new_AGEMA_signal_16300, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, RoundInput[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16308, new_AGEMA_signal_16307, new_AGEMA_signal_16306, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, RoundInput[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16314, new_AGEMA_signal_16313, new_AGEMA_signal_16312, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16320, new_AGEMA_signal_16319, new_AGEMA_signal_16318, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, RoundInput[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16794, new_AGEMA_signal_16793, new_AGEMA_signal_16792, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16326, new_AGEMA_signal_16325, new_AGEMA_signal_16324, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, RoundInput[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16800, new_AGEMA_signal_16799, new_AGEMA_signal_16798, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16806, new_AGEMA_signal_16805, new_AGEMA_signal_16804, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundInput[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16332, new_AGEMA_signal_16331, new_AGEMA_signal_16330, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16338, new_AGEMA_signal_16337, new_AGEMA_signal_16336, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundInput[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16344, new_AGEMA_signal_16343, new_AGEMA_signal_16342, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16350, new_AGEMA_signal_16349, new_AGEMA_signal_16348, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16812, new_AGEMA_signal_16811, new_AGEMA_signal_16810, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, RoundInput[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16356, new_AGEMA_signal_16355, new_AGEMA_signal_16354, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16818, new_AGEMA_signal_16817, new_AGEMA_signal_16816, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, RoundInput[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16824, new_AGEMA_signal_16823, new_AGEMA_signal_16822, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16362, new_AGEMA_signal_16361, new_AGEMA_signal_16360, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, RoundInput[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16368, new_AGEMA_signal_16367, new_AGEMA_signal_16366, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16374, new_AGEMA_signal_16373, new_AGEMA_signal_16372, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, RoundInput[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16380, new_AGEMA_signal_16379, new_AGEMA_signal_16378, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16830, new_AGEMA_signal_16829, new_AGEMA_signal_16828, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, RoundInput[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16386, new_AGEMA_signal_16385, new_AGEMA_signal_16384, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, RoundInput[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16836, new_AGEMA_signal_16835, new_AGEMA_signal_16834, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16842, new_AGEMA_signal_16841, new_AGEMA_signal_16840, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, RoundInput[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16392, new_AGEMA_signal_16391, new_AGEMA_signal_16390, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16398, new_AGEMA_signal_16397, new_AGEMA_signal_16396, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, RoundInput[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16404, new_AGEMA_signal_16403, new_AGEMA_signal_16402, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16410, new_AGEMA_signal_16409, new_AGEMA_signal_16408, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, RoundInput[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16848, new_AGEMA_signal_16847, new_AGEMA_signal_16846, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16416, new_AGEMA_signal_16415, new_AGEMA_signal_16414, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, RoundInput[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16854, new_AGEMA_signal_16853, new_AGEMA_signal_16852, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16860, new_AGEMA_signal_16859, new_AGEMA_signal_16858, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16422, new_AGEMA_signal_16421, new_AGEMA_signal_16420, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, RoundInput[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16428, new_AGEMA_signal_16427, new_AGEMA_signal_16426, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, RoundInput[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16434, new_AGEMA_signal_16433, new_AGEMA_signal_16432, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundInput[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16440, new_AGEMA_signal_16439, new_AGEMA_signal_16438, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, RoundInput[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16866, new_AGEMA_signal_16865, new_AGEMA_signal_16864, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundInput[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16446, new_AGEMA_signal_16445, new_AGEMA_signal_16444, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, RoundInput[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16872, new_AGEMA_signal_16871, new_AGEMA_signal_16870, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundInput[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16878, new_AGEMA_signal_16877, new_AGEMA_signal_16876, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, RoundInput[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16452, new_AGEMA_signal_16451, new_AGEMA_signal_16450, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundInput[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16458, new_AGEMA_signal_16457, new_AGEMA_signal_16456, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, RoundInput[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16464, new_AGEMA_signal_16463, new_AGEMA_signal_16462, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, RoundInput[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16470, new_AGEMA_signal_16469, new_AGEMA_signal_16468, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, RoundInput[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16884, new_AGEMA_signal_16883, new_AGEMA_signal_16882, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, RoundInput[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16476, new_AGEMA_signal_16475, new_AGEMA_signal_16474, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, RoundInput[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16890, new_AGEMA_signal_16889, new_AGEMA_signal_16888, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, RoundInput[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16896, new_AGEMA_signal_16895, new_AGEMA_signal_16894, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, RoundInput[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16482, new_AGEMA_signal_16481, new_AGEMA_signal_16480, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, RoundInput[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16488, new_AGEMA_signal_16487, new_AGEMA_signal_16486, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, RoundInput[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16494, new_AGEMA_signal_16493, new_AGEMA_signal_16492, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, RoundInput[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16500, new_AGEMA_signal_16499, new_AGEMA_signal_16498, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, RoundInput[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16902, new_AGEMA_signal_16901, new_AGEMA_signal_16900, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, RoundInput[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16506, new_AGEMA_signal_16505, new_AGEMA_signal_16504, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, RoundInput[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16908, new_AGEMA_signal_16907, new_AGEMA_signal_16906, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, RoundInput[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16914, new_AGEMA_signal_16913, new_AGEMA_signal_16912, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, RoundInput[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16512, new_AGEMA_signal_16511, new_AGEMA_signal_16510, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, RoundInput[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16518, new_AGEMA_signal_16517, new_AGEMA_signal_16516, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, RoundInput[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16524, new_AGEMA_signal_16523, new_AGEMA_signal_16522, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, RoundInput[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16530, new_AGEMA_signal_16529, new_AGEMA_signal_16528, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, RoundInput[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16920, new_AGEMA_signal_16919, new_AGEMA_signal_16918, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, RoundInput[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16536, new_AGEMA_signal_16535, new_AGEMA_signal_16534, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, RoundInput[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16926, new_AGEMA_signal_16925, new_AGEMA_signal_16924, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, RoundInput[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16932, new_AGEMA_signal_16931, new_AGEMA_signal_16930, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, RoundInput[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16542, new_AGEMA_signal_16541, new_AGEMA_signal_16540, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, RoundInput[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16548, new_AGEMA_signal_16547, new_AGEMA_signal_16546, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, RoundInput[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16554, new_AGEMA_signal_16553, new_AGEMA_signal_16552, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, RoundInput[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16560, new_AGEMA_signal_16559, new_AGEMA_signal_16558, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundInput[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16938, new_AGEMA_signal_16937, new_AGEMA_signal_16936, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, RoundInput[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16566, new_AGEMA_signal_16565, new_AGEMA_signal_16564, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundInput[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16944, new_AGEMA_signal_16943, new_AGEMA_signal_16942, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, RoundInput[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16950, new_AGEMA_signal_16949, new_AGEMA_signal_16948, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, RoundInput[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16572, new_AGEMA_signal_16571, new_AGEMA_signal_16570, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16578, new_AGEMA_signal_16577, new_AGEMA_signal_16576, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, RoundInput[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16584, new_AGEMA_signal_16583, new_AGEMA_signal_16582, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16590, new_AGEMA_signal_16589, new_AGEMA_signal_16588, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, RoundInput[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16956, new_AGEMA_signal_16955, new_AGEMA_signal_16954, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16596, new_AGEMA_signal_16595, new_AGEMA_signal_16594, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, RoundInput[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16962, new_AGEMA_signal_16961, new_AGEMA_signal_16960, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16968, new_AGEMA_signal_16967, new_AGEMA_signal_16966, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, RoundInput[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16602, new_AGEMA_signal_16601, new_AGEMA_signal_16600, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16608, new_AGEMA_signal_16607, new_AGEMA_signal_16606, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16614, new_AGEMA_signal_16613, new_AGEMA_signal_16612, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, RoundInput[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16620, new_AGEMA_signal_16619, new_AGEMA_signal_16618, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16974, new_AGEMA_signal_16973, new_AGEMA_signal_16972, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, RoundInput[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16626, new_AGEMA_signal_16625, new_AGEMA_signal_16624, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16980, new_AGEMA_signal_16979, new_AGEMA_signal_16978, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, RoundInput[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16986, new_AGEMA_signal_16985, new_AGEMA_signal_16984, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16632, new_AGEMA_signal_16631, new_AGEMA_signal_16630, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, RoundInput[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16638, new_AGEMA_signal_16637, new_AGEMA_signal_16636, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16644, new_AGEMA_signal_16643, new_AGEMA_signal_16642, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, RoundInput[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16650, new_AGEMA_signal_16649, new_AGEMA_signal_16648, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, RoundInput[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16992, new_AGEMA_signal_16991, new_AGEMA_signal_16990, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16656, new_AGEMA_signal_16655, new_AGEMA_signal_16654, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, RoundInput[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16998, new_AGEMA_signal_16997, new_AGEMA_signal_16996, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_17004, new_AGEMA_signal_17003, new_AGEMA_signal_17002, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, RoundInput[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16662, new_AGEMA_signal_16661, new_AGEMA_signal_16660, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16668, new_AGEMA_signal_16667, new_AGEMA_signal_16666, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, RoundInput[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16674, new_AGEMA_signal_16673, new_AGEMA_signal_16672, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[127]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15198, new_AGEMA_signal_15197, new_AGEMA_signal_15196, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15861, new_AGEMA_signal_15860, new_AGEMA_signal_15859, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15867, new_AGEMA_signal_15866, new_AGEMA_signal_15865, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15873, new_AGEMA_signal_15872, new_AGEMA_signal_15871, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15879, new_AGEMA_signal_15878, new_AGEMA_signal_15877, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15885, new_AGEMA_signal_15884, new_AGEMA_signal_15883, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15891, new_AGEMA_signal_15890, new_AGEMA_signal_15889, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15897, new_AGEMA_signal_15896, new_AGEMA_signal_15895, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15204, new_AGEMA_signal_15203, new_AGEMA_signal_15202, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15903, new_AGEMA_signal_15902, new_AGEMA_signal_15901, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15909, new_AGEMA_signal_15908, new_AGEMA_signal_15907, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15915, new_AGEMA_signal_15914, new_AGEMA_signal_15913, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15921, new_AGEMA_signal_15920, new_AGEMA_signal_15919, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15927, new_AGEMA_signal_15926, new_AGEMA_signal_15925, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15933, new_AGEMA_signal_15932, new_AGEMA_signal_15931, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15939, new_AGEMA_signal_15938, new_AGEMA_signal_15937, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15210, new_AGEMA_signal_15209, new_AGEMA_signal_15208, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15945, new_AGEMA_signal_15944, new_AGEMA_signal_15943, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15951, new_AGEMA_signal_15950, new_AGEMA_signal_15949, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15957, new_AGEMA_signal_15956, new_AGEMA_signal_15955, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15963, new_AGEMA_signal_15962, new_AGEMA_signal_15961, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15969, new_AGEMA_signal_15968, new_AGEMA_signal_15967, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15975, new_AGEMA_signal_15974, new_AGEMA_signal_15973, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15981, new_AGEMA_signal_15980, new_AGEMA_signal_15979, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15987, new_AGEMA_signal_15986, new_AGEMA_signal_15985, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16680, new_AGEMA_signal_16679, new_AGEMA_signal_16678, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16686, new_AGEMA_signal_16685, new_AGEMA_signal_16684, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16692, new_AGEMA_signal_16691, new_AGEMA_signal_16690, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16698, new_AGEMA_signal_16697, new_AGEMA_signal_16696, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16704, new_AGEMA_signal_16703, new_AGEMA_signal_16702, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16710, new_AGEMA_signal_16709, new_AGEMA_signal_16708, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16716, new_AGEMA_signal_16715, new_AGEMA_signal_16714, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14526, new_AGEMA_signal_14525, new_AGEMA_signal_14524, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundKey[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15216, new_AGEMA_signal_15215, new_AGEMA_signal_15214, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, RoundKey[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15222, new_AGEMA_signal_15221, new_AGEMA_signal_15220, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundKey[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15228, new_AGEMA_signal_15227, new_AGEMA_signal_15226, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKey[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15234, new_AGEMA_signal_15233, new_AGEMA_signal_15232, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundKey[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15240, new_AGEMA_signal_15239, new_AGEMA_signal_15238, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKey[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15246, new_AGEMA_signal_15245, new_AGEMA_signal_15244, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundKey[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15252, new_AGEMA_signal_15251, new_AGEMA_signal_15250, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKey[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14532, new_AGEMA_signal_14531, new_AGEMA_signal_14530, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, RoundKey[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15258, new_AGEMA_signal_15257, new_AGEMA_signal_15256, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundKey[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15264, new_AGEMA_signal_15263, new_AGEMA_signal_15262, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, RoundKey[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15270, new_AGEMA_signal_15269, new_AGEMA_signal_15268, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundKey[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15276, new_AGEMA_signal_15275, new_AGEMA_signal_15274, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, RoundKey[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15282, new_AGEMA_signal_15281, new_AGEMA_signal_15280, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundKey[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15288, new_AGEMA_signal_15287, new_AGEMA_signal_15286, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, RoundKey[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15294, new_AGEMA_signal_15293, new_AGEMA_signal_15292, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundKey[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14538, new_AGEMA_signal_14537, new_AGEMA_signal_14536, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, RoundKey[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15300, new_AGEMA_signal_15299, new_AGEMA_signal_15298, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundKey[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15306, new_AGEMA_signal_15305, new_AGEMA_signal_15304, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundKey[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15312, new_AGEMA_signal_15311, new_AGEMA_signal_15310, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, RoundKey[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15318, new_AGEMA_signal_15317, new_AGEMA_signal_15316, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundKey[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15324, new_AGEMA_signal_15323, new_AGEMA_signal_15322, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, RoundKey[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15330, new_AGEMA_signal_15329, new_AGEMA_signal_15328, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundKey[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15336, new_AGEMA_signal_15335, new_AGEMA_signal_15334, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, RoundKey[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15342, new_AGEMA_signal_15341, new_AGEMA_signal_15340, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundKey[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15993, new_AGEMA_signal_15992, new_AGEMA_signal_15991, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, RoundKey[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15999, new_AGEMA_signal_15998, new_AGEMA_signal_15997, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundKey[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, new_AGEMA_signal_16003, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, RoundKey[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, new_AGEMA_signal_16009, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, RoundKey[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16017, new_AGEMA_signal_16016, new_AGEMA_signal_16015, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, RoundKey[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16023, new_AGEMA_signal_16022, new_AGEMA_signal_16021, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, RoundKey[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, new_AGEMA_signal_16027, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, RoundKey[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13896, new_AGEMA_signal_13895, new_AGEMA_signal_13894, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKey[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14544, new_AGEMA_signal_14543, new_AGEMA_signal_14542, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, RoundKey[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14550, new_AGEMA_signal_14549, new_AGEMA_signal_14548, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKey[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14556, new_AGEMA_signal_14555, new_AGEMA_signal_14554, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, RoundKey[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14562, new_AGEMA_signal_14561, new_AGEMA_signal_14560, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKey[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14568, new_AGEMA_signal_14567, new_AGEMA_signal_14566, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, RoundKey[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14574, new_AGEMA_signal_14573, new_AGEMA_signal_14572, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, RoundKey[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14580, new_AGEMA_signal_14579, new_AGEMA_signal_14578, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, RoundKey[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13902, new_AGEMA_signal_13901, new_AGEMA_signal_13900, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, RoundKey[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14586, new_AGEMA_signal_14585, new_AGEMA_signal_14584, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, RoundKey[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14592, new_AGEMA_signal_14591, new_AGEMA_signal_14590, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, RoundKey[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14598, new_AGEMA_signal_14597, new_AGEMA_signal_14596, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, RoundKey[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14604, new_AGEMA_signal_14603, new_AGEMA_signal_14602, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, RoundKey[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14610, new_AGEMA_signal_14609, new_AGEMA_signal_14608, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, RoundKey[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14616, new_AGEMA_signal_14615, new_AGEMA_signal_14614, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, RoundKey[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14622, new_AGEMA_signal_14621, new_AGEMA_signal_14620, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, RoundKey[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13908, new_AGEMA_signal_13907, new_AGEMA_signal_13906, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, RoundKey[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14628, new_AGEMA_signal_14627, new_AGEMA_signal_14626, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, RoundKey[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14634, new_AGEMA_signal_14633, new_AGEMA_signal_14632, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, RoundKey[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14640, new_AGEMA_signal_14639, new_AGEMA_signal_14638, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, RoundKey[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14646, new_AGEMA_signal_14645, new_AGEMA_signal_14644, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, RoundKey[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14652, new_AGEMA_signal_14651, new_AGEMA_signal_14650, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, RoundKey[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14658, new_AGEMA_signal_14657, new_AGEMA_signal_14656, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, RoundKey[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14664, new_AGEMA_signal_14663, new_AGEMA_signal_14662, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, RoundKey[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14670, new_AGEMA_signal_14669, new_AGEMA_signal_14668, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, RoundKey[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15348, new_AGEMA_signal_15347, new_AGEMA_signal_15346, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, RoundKey[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15354, new_AGEMA_signal_15353, new_AGEMA_signal_15352, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, RoundKey[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15360, new_AGEMA_signal_15359, new_AGEMA_signal_15358, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, RoundKey[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15366, new_AGEMA_signal_15365, new_AGEMA_signal_15364, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, RoundKey[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15372, new_AGEMA_signal_15371, new_AGEMA_signal_15370, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, RoundKey[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15378, new_AGEMA_signal_15377, new_AGEMA_signal_15376, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, RoundKey[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_15384, new_AGEMA_signal_15383, new_AGEMA_signal_15382, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKey[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13398, new_AGEMA_signal_13397, new_AGEMA_signal_13396, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, RoundKey[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13914, new_AGEMA_signal_13913, new_AGEMA_signal_13912, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKey[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13920, new_AGEMA_signal_13919, new_AGEMA_signal_13918, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, RoundKey[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13926, new_AGEMA_signal_13925, new_AGEMA_signal_13924, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKey[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13932, new_AGEMA_signal_13931, new_AGEMA_signal_13930, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundKey[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13938, new_AGEMA_signal_13937, new_AGEMA_signal_13936, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, RoundKey[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13944, new_AGEMA_signal_13943, new_AGEMA_signal_13942, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundKey[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13950, new_AGEMA_signal_13949, new_AGEMA_signal_13948, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, RoundKey[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13404, new_AGEMA_signal_13403, new_AGEMA_signal_13402, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundKey[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13956, new_AGEMA_signal_13955, new_AGEMA_signal_13954, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, RoundKey[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13962, new_AGEMA_signal_13961, new_AGEMA_signal_13960, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundKey[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13968, new_AGEMA_signal_13967, new_AGEMA_signal_13966, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, RoundKey[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13974, new_AGEMA_signal_13973, new_AGEMA_signal_13972, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundKey[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13980, new_AGEMA_signal_13979, new_AGEMA_signal_13978, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, RoundKey[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13986, new_AGEMA_signal_13985, new_AGEMA_signal_13984, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, RoundKey[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13992, new_AGEMA_signal_13991, new_AGEMA_signal_13990, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundKey[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13410, new_AGEMA_signal_13409, new_AGEMA_signal_13408, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, RoundKey[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_13998, new_AGEMA_signal_13997, new_AGEMA_signal_13996, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundKey[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14004, new_AGEMA_signal_14003, new_AGEMA_signal_14002, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, RoundKey[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14010, new_AGEMA_signal_14009, new_AGEMA_signal_14008, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundKey[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14016, new_AGEMA_signal_14015, new_AGEMA_signal_14014, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, RoundKey[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14022, new_AGEMA_signal_14021, new_AGEMA_signal_14020, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundKey[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14028, new_AGEMA_signal_14027, new_AGEMA_signal_14026, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, RoundKey[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14034, new_AGEMA_signal_14033, new_AGEMA_signal_14032, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundKey[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14040, new_AGEMA_signal_14039, new_AGEMA_signal_14038, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundKey[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14676, new_AGEMA_signal_14675, new_AGEMA_signal_14674, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, RoundKey[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14682, new_AGEMA_signal_14681, new_AGEMA_signal_14680, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundKey[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14688, new_AGEMA_signal_14687, new_AGEMA_signal_14686, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, RoundKey[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14694, new_AGEMA_signal_14693, new_AGEMA_signal_14692, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundKey[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14700, new_AGEMA_signal_14699, new_AGEMA_signal_14698, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, RoundKey[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14706, new_AGEMA_signal_14705, new_AGEMA_signal_14704, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundKey[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_14712, new_AGEMA_signal_14711, new_AGEMA_signal_14710, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_36608), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_36612), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_36616), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_36620), .Q (RoundCounter[3]), .QN () ) ;
endmodule
