module LED_Top(x, y);
 input [193:0] x;
 output [64:0] y;

 wire [3862:0] t;
  FX FX_inst(.x({t[1354], t[1353], t[1352], t[1351], t[1350], t[1349], t[1348], t[1347], t[1346], t[1345], t[1344], t[1343], t[1342], t[1341], t[1340], t[1339], t[1338], t[1337], t[1336], t[1335], t[1334], t[1333], t[1332], t[1331], t[1330], t[1329], t[1328], t[1327], t[1326], t[1325], t[1324], t[1323], t[1322], t[1321], t[1320], t[1319], t[1318], t[1317], t[1316], t[1315], t[1314], t[1313], t[1312], t[1311], t[1310], t[1309], t[1308], t[1307], t[1306], t[1305], t[1304], t[1303], t[1302], t[1301], t[1300], t[1299], t[1298], t[1297], t[1296], t[1295], t[1294], t[1293], t[1292], t[1291], t[1290], t[1289], t[1288], t[1287], t[1286], t[1285], t[1284], t[1283], t[1282], t[1281], t[1280], t[1279], t[1278], t[1277], t[1276], t[1275], t[1274], t[1273], t[1272], t[1271], t[1270], t[1269], t[1268], t[1267], t[1266], t[1265], t[1264], t[1263], t[1262], t[1261], t[1260], t[1259], t[1258], t[1257], t[1256], t[1255], t[1254], t[1253], t[1252], t[1251], t[1250], t[1249], t[1248], t[1247], t[1246], t[1245], t[1244], t[1243], t[1242], t[1241], t[1240], t[1239], t[1238], t[1237], t[1236], t[1235], t[1234], t[1233], t[1232], t[1231], t[1230], t[1229], t[1228], t[1227], t[1226], t[1225], t[1224], t[1223], t[1222], t[1221], t[1220], t[1219], t[1218], t[1217], t[1216], t[1215], t[1214], t[1213], t[1212], t[1211], t[1210], t[1209], t[1208], t[1207], t[1206], t[1205], t[1204], t[1203], t[1202], t[1201], t[1200], t[1199], t[1198], t[1197], t[1196], t[1195], t[1194], t[1193], t[1192], t[1191], t[1190], t[1189], t[1188], t[1187], t[1186], t[1185], t[1184], t[1183], t[1182], t[1181], t[1180], t[1179], t[1178], t[1177], t[1176], t[1175], t[1174], t[1173], t[1172], t[1171], t[1170], t[1169], t[1168], t[1167], t[1166], t[1165], t[1164], t[1163], t[1162], t[1161], t[1160], t[1159], t[1158], t[1157], t[1156], t[1155], t[1154], t[1153], t[1152], t[1151], t[1150], t[1149], t[1148], t[1147], t[1146], t[1145], t[1144], t[1143], t[1142], t[1141], t[1140], t[1139], t[1138], t[1137], t[1136], t[1135], t[1134], t[1133], t[1132], t[1131], t[1130], t[1129], t[1128], t[1127], t[1126], t[1125], t[1124], t[1123], t[1122], t[1121], t[1120], t[1119], t[1118], t[1117], t[1116], t[1115], t[1114], t[1113], t[1112], t[1111], t[1110], t[1109], t[1108], t[1107], t[1106], t[1105], t[1104], t[1103], t[1102], t[1101], t[1100], t[1099], t[1098], t[1097], t[1096], t[1095], t[1094], t[1093], t[1092], t[1091], t[1090], t[1089], t[1088], t[1087], t[1086], t[1085], t[1084], t[1083], t[1082], t[1081], t[1080], t[1079], t[1078], t[1077], t[1076], t[1075], t[1074], t[1073], t[1072], t[1071], t[1070], t[1069], t[1068], t[1067], t[1066], t[1065], t[1064], t[1063], t[1062], t[1061], t[1060], t[1059], t[1058], t[1057], t[1056], t[1055], t[1054], t[1053], t[1052], t[1051], t[1050], t[1049], t[1048], t[1047], t[1046], t[1045], t[1044], t[1043], t[1042], t[1041], t[1040], t[1039], t[1038], t[1037], t[1036], t[1035], t[1034], t[1033], t[1032], t[1031], t[1030], t[1029], t[1028], t[1027], t[1026], t[1025], t[1024], t[1023], t[1022], t[1021], t[1020], t[1019], t[1018], t[1017], t[1016], t[1015], t[1014], t[1013], t[1012], t[1011], t[1010], t[1009], t[1008], t[1007], t[1006], t[1005], t[1004], t[1003], t[1002], t[1001], t[1000], t[999], t[998], t[997], t[996], t[995], t[994], t[993], t[992], t[991], t[990], t[989], t[988], t[987], t[986], t[985], t[984], t[983], t[982], t[981], t[980], t[979], t[978], t[977], t[976], t[975], t[974], t[973], t[972], t[971], t[970], t[969], t[968], t[967], t[966], t[965], t[964], t[963], t[962], t[961], t[960], t[959], t[958], t[957], t[956], t[955], t[954], t[953], t[952], t[951], t[950], t[949], t[948], t[947], t[946], t[945], t[944], t[943], t[942], t[941], t[940], t[939], t[938], t[937], t[936], t[935], t[934], t[933], t[932], t[931], t[930], t[929], t[928], t[927], t[926], t[925], t[924], t[923], t[922], t[921], t[920], t[919], t[918], t[917], t[916], t[915], t[914], t[913], t[912], t[911], t[910], t[909], t[908], t[907], t[906], t[905], t[904], t[903], t[902], t[901], t[900], t[899], t[898], t[897], t[896], t[895], t[894], t[893], t[892], t[891], t[890], t[889], t[888], t[887], t[886], t[885], t[884], t[883], t[882], t[881], t[880], t[879], t[878], t[877], t[876], t[875], t[874], t[873], t[872], t[871], t[870], t[869], t[868], t[867], t[866], t[865], t[864], t[863], t[862], t[861], t[860], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[852], t[851], t[850], t[849], t[848], t[847], t[846], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[803], t[802], t[801], t[800], t[799], t[798], t[797], t[796], t[795], t[794], t[793], t[792], t[791], t[790], t[789], t[788], t[787], t[786], t[785], t[784], t[783], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[761], t[760], t[759], t[758], t[757], t[756], t[755], t[754], t[753], t[752], t[751], t[750], t[749], t[748], t[747], t[746], t[745], t[744], t[743], t[742], t[741], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[719], t[718], t[717], t[716], t[715], t[714], t[713], t[712], t[711], t[710], t[709], t[708], t[707], t[706], t[705], t[704], t[703], t[702], t[701], t[700], t[699], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[684], t[683], t[682], t[681], t[680], t[679], t[678], t[677], t[676], t[675], t[674], t[673], t[672], t[671], t[670], t[669], t[668], t[667], t[666], t[665], t[664], t[663], t[662], t[661], t[660], t[659], t[658], t[657], t[656], t[655], t[654], t[653], t[652], t[651], t[650], t[649], t[648], t[647], t[646], t[645], t[644], t[643], t[642], t[641], t[640], t[639], t[638], t[637], t[636], t[635], t[634], t[633], t[632], t[631], t[630], t[629], t[628], t[627], t[626], t[625], t[624], t[623], t[622], t[621], t[620], t[619], t[618], t[617], t[616], t[615], t[614], t[613], t[612], t[611], t[610], t[609], t[608], t[607], t[606], t[605], t[604], t[603], t[602], t[601], t[600], t[599], t[598], t[597], t[596], t[595], t[594], t[593], t[592], t[591], t[590], t[589], t[588], t[587], t[586], t[585], t[584], t[583], t[582], t[581], t[580], t[579], t[578], t[577], t[576], t[575], t[574], t[573], t[572], t[571], t[570], t[569], t[568], t[567], t[566], t[565], t[564], t[563], t[562], t[561], t[560], t[559], t[558], t[557], t[556], t[555], t[554], t[553], t[552], t[551], t[550], t[549], t[548], t[547], t[546], t[545], t[544], t[543], t[542], t[541], t[540], t[539], t[538], t[537], t[536], t[535], t[534], t[533], t[532], t[531], t[530], t[529], t[528], t[527], t[526], t[525], t[524], t[523], t[522], t[521], t[520], t[519], t[518], t[517], t[516], t[515], t[514], t[513], t[512], t[511], t[510], t[509], t[508], t[507], t[506], t[505], t[504], t[503], t[502], t[501], t[500], t[499], t[498], t[497], t[496], t[495], t[494], t[493], t[492], t[491], t[490], t[489], t[488], t[487], t[486], t[485], t[484], t[483], t[482], t[481], t[480], t[479], t[478], t[477], t[476], t[475], t[474], t[473], t[472], t[471], t[470], t[469], t[468], t[467], t[466], t[465], t[464], t[463], t[462], t[461], t[460], t[459], t[458], t[457], t[456], t[455], t[454], t[453], t[452], t[451], t[450], t[449], t[448], t[447], t[446], t[445], t[444], t[443], t[442], t[441], t[440], t[439], t[438], t[437], t[436], t[435], t[434], t[433], t[432], t[431], t[430], t[429], t[428], t[427], t[426], t[425], t[424], t[423], t[422], t[421], t[420], t[419], t[418], t[417], t[416], t[415], t[414], t[413], t[412], t[411], t[410], t[409], t[408], t[407], t[406], t[405], t[404], t[403], t[402], t[401], t[400], t[399], t[398], t[397], t[396], t[395], t[394], t[393], t[392], t[391], t[390], t[389], t[388], t[387], t[386], t[385], t[384], t[383], t[382], t[381], t[380], t[379], t[378], t[377], t[376], t[375], t[374], t[373], t[372], t[371], t[370], t[369], t[368], t[367], t[366], t[365], t[364], t[363], t[362], t[361], t[360], t[359], t[358], t[357], t[356], t[355], t[354], t[353], t[352], t[351], t[350], t[349], t[348], t[347], t[346], t[345], t[344], t[343], t[342], t[341], t[340], t[339], t[338], t[337], t[336], t[335], t[334], t[333], t[332], t[331], t[330], t[329], t[328], t[327], t[326], t[325], t[324], t[323], t[322], t[321], t[320], t[319], t[318], t[317], t[316], t[315], t[314], t[313], t[312], t[311], t[310], t[309], t[308], t[307], t[306], t[305], t[304], t[303], t[302], t[301], t[300], t[299], t[298], t[297], t[296], t[295], t[294], t[293], t[292], t[291], t[290], t[289], t[288], t[287], t[286], t[285], t[284], t[283], t[282], t[281], t[280], t[279], t[278], t[277], t[276], t[275], t[274], t[273], t[272], t[271], t[270], t[269], t[268], t[267], t[266], t[265], t[264], t[263], t[262], t[261], t[260], t[259], t[258], t[257], t[256], t[255], t[254], t[253], t[252], t[251], t[250], t[249], t[248], t[247], t[246], t[245], t[244], t[243], t[242], t[241], t[240], t[239], t[238], t[237], t[236], t[235], t[234], t[233], t[232], t[231], t[230], t[229], t[228], t[227], t[226], t[225], t[224], t[223], t[222], t[221], t[220], t[219], t[218], t[217], t[216], t[215], t[214], t[213], t[212], t[211], t[210], t[209], t[208], t[207], t[206], t[205], t[204], t[203], t[202], t[201], t[200], t[199], t[198], t[197], t[196], t[195], t[194], t[193], t[192], t[191], t[190], t[189], t[188], t[187], t[186], t[185], t[184], t[183], t[182], t[181], t[180], t[179], t[178], t[177], t[176], t[175], t[174], t[173], t[172], t[171], t[170], t[169], t[168], t[167], t[166], t[165], t[164], t[163], t[162], t[161], t[160], t[159], t[158], t[157], t[156], t[155], t[154], t[153], t[152], t[151], t[150], t[149], t[148], t[147], t[146], t[145], t[144], t[143], t[142], t[141], t[140], t[139], t[138], t[137], t[136], t[135], t[134], t[133], t[132], t[131], t[130], t[129], t[128], t[127], t[126], t[125], t[124], t[123], t[122], t[121], t[120], t[119], t[118], t[117], t[116], t[115], t[114], t[113], t[112], t[111], t[110], t[109], t[108], t[107], t[106], t[105], t[104], t[103], t[102], t[101], t[100], t[99], t[98], t[97], t[96], t[95], t[94], t[93], t[92], t[91], t[90], t[89], t[88], t[87], t[86], t[85], t[84], t[83], t[82], t[81], t[80], t[79], t[78], t[77], t[76], t[75], t[74], t[73], t[72], t[71], t[70], t[69], t[68], t[67], t[66], t[65], t[64], t[63], t[62], t[61], t[60], t[59], t[58], t[57], t[56], t[55], t[54], t[53], t[52], t[51], t[50], t[49], t[48], t[47], t[46], t[45], t[44], t[43], t[42], t[41], t[40], t[39], t[38], t[37], t[36], t[35], t[34], t[33], t[32], t[31], t[30], t[29], t[28], t[27], t[26], t[25], t[24], t[23], t[22], t[21], t[20], t[19], t[18], t[17], t[16], t[15], t[14], t[13], t[12], t[11], t[10], t[9], t[8], t[7], t[6], t[5], t[4], t[3], t[2], t[1], t[0]}), .y({t[2438], t[2437], t[2436], t[2435], t[2434], t[2433], t[2432], t[2431], t[2430], t[2429], t[2428], t[2427], t[2426], t[2425], t[2424], t[2423], t[2422], t[2421], t[2420], t[2419], t[2418], t[2417], t[2416], t[2415], t[2414], t[2413], t[2412], t[2411], t[2410], t[2409], t[2408], t[2407], t[2406], t[2405], t[2404], t[2403], t[2402], t[2401], t[2400], t[2399], t[2398], t[2397], t[2396], t[2395], t[2394], t[2393], t[2392], t[2391], t[2390], t[2389], t[2388], t[2387], t[2386], t[2385], t[2384], t[2383], t[2382], t[2381], t[2380], t[2379], t[2378], t[2377], t[2376], t[2375], t[2374], t[2373], t[2372], t[2371], t[2370], t[2369], t[2368], t[2367], t[2366], t[2365], t[2364], t[2363], t[2362], t[2361], t[2360], t[2359], t[2358], t[2357], t[2356], t[2355], t[2354], t[2353], t[2352], t[2351], t[2350], t[2349], t[2348], t[2347], t[2346], t[2345], t[2344], t[2343], t[2342], t[2341], t[2340], t[2339], t[2338], t[2337], t[2336], t[2335], t[2334], t[2333], t[2332], t[2331], t[2330], t[2329], t[2328], t[2327], t[2326], t[2325], t[2324], t[2323], t[2322], t[2321], t[2320], t[2319], t[2318], t[2317], t[2316], t[2315], t[2314], t[2313], t[2312], t[2311], t[2310], t[2309], t[2308], t[2307], t[2306], t[2305], t[2304], t[2303], t[2302], t[2301], t[2300], t[2299], t[2298], t[2297], t[2296], t[2295], t[2294], t[2293], t[2292], t[2291], t[2290], t[2289], t[2288], t[2287], t[2286], t[2285], t[2284], t[2283], t[2282], t[2281], t[2280], t[2279], t[2278], t[2277], t[2276], t[2275], t[2274], t[2273], t[2272], t[2271], t[2270], t[2269], t[2268], t[2267], t[2266], t[2265], t[2264], t[2263], t[2262], t[2261], t[2260], t[2259], t[2258], t[2257], t[2256], t[2255], t[2254], t[2253], t[2252], t[2251], t[2250], t[2249], t[2248], t[2247], t[2246], t[2245], t[2244], t[2243], t[2242], t[2241], t[2240], t[2239], t[2238], t[2237], t[2236], t[2235], t[2234], t[2233], t[2232], t[2231], t[2230], t[2229], t[2228], t[2227], t[2226], t[2225], t[2224], t[2223], t[2222], t[2221], t[2220], t[2219], t[2218], t[2217], t[2216], t[2215], t[2214], t[2213], t[2212], t[2211], t[2210], t[2209], t[2208], t[2207], t[2206], t[2205], t[2204], t[2203], t[2202], t[2201], t[2200], t[2199], t[2198], t[2197], t[2196], t[2195], t[2194], t[2193], t[2192], t[2191], t[2190], t[2189], t[2188], t[2187], t[2186], t[2185], t[2184], t[2183], t[2182], t[2181], t[2180], t[2179], t[2178], t[2177], t[2176], t[2175], t[2174], t[2173], t[2172], t[2171], t[2170], t[2169], t[2168], t[2167], t[2166], t[2165], t[2164], t[2163], t[2162], t[2161], t[2160], t[2159], t[2158], t[2157], t[2156], t[2155], t[2154], t[2153], t[2152], t[2151], t[2150], t[2149], t[2148], t[2147], t[2146], t[2145], t[2144], t[2143], t[2142], t[2141], t[2140], t[2139], t[2138], t[2137], t[2136], t[2135], t[2134], t[2133], t[2132], t[2131], t[2130], t[2129], t[2128], t[2127], t[2126], t[2125], t[2124], t[2123], t[2122], t[2121], t[2120], t[2119], t[2118], t[2117], t[2116], t[2115], t[2114], t[2113], t[2112], t[2111], t[2110], t[2109], t[2108], t[2107], t[2106], t[2105], t[2104], t[2103], t[2102], t[2101], t[2100], t[2099], t[2098], t[2097], t[2096], t[2095], t[2094], t[2093], t[2092], t[2091], t[2090], t[2089], t[2088], t[2087], t[2086], t[2085], t[2084], t[2083], t[2082], t[2081], t[2080], t[2079], t[2078], t[2077], t[2076], t[2075], t[2074], t[2073], t[2072], t[2071], t[2070], t[2069], t[2068], t[2067], t[2066], t[2065], t[2064], t[2063], t[2062], t[2061], t[2060], t[2059], t[2058], t[2057], t[2056], t[2055], t[2054], t[2053], t[2052], t[2051], t[2050], t[2049], t[2048], t[2047], t[2046], t[2045], t[2044], t[2043], t[2042], t[2041], t[2040], t[2039], t[2038], t[2037], t[2036], t[2035], t[2034], t[2033], t[2032], t[2031], t[2030], t[2029], t[2028], t[2027], t[2026], t[2025], t[2024], t[2023], t[2022], t[2021], t[2020], t[2019], t[2018], t[2017], t[2016], t[2015], t[2014], t[2013], t[2012], t[2011], t[2010], t[2009], t[2008], t[2007], t[2006], t[2005], t[2004], t[2003], t[2002], t[2001], t[2000], t[1999], t[1998], t[1997], t[1996], t[1995], t[1994], t[1993], t[1992], t[1991], t[1990], t[1989], t[1988], t[1987], t[1986], t[1985], t[1984], t[1983], t[1982], t[1981], t[1980], t[1979], t[1978], t[1977], t[1976], t[1975], t[1974], t[1973], t[1972], t[1971], t[1970], t[1969], t[1968], t[1967], t[1966], t[1965], t[1964], t[1963], t[1962], t[1961], t[1960], t[1959], t[1958], t[1957], t[1956], t[1955], t[1954], t[1953], t[1952], t[1951], t[1950], t[1949], t[1948], t[1947], t[1946], t[1945], t[1944], t[1943], t[1942], t[1941], t[1940], t[1939], t[1938], t[1937], t[1936], t[1935], t[1934], t[1933], t[1932], t[1931], t[1930], t[1929], t[1928], t[1927], t[1926], t[1925], t[1924], t[1923], t[1922], t[1921], t[1920], t[1919], t[1918], t[1917], t[1916], t[1915], t[1914], t[1913], t[1912], t[1911], t[1910], t[1909], t[1908], t[1907], t[1906], t[1905], t[1904], t[1903], t[1902], t[1901], t[1900], t[1899], t[1898], t[1897], t[1896], t[1895], t[1894], t[1893], t[1892], t[1891], t[1890], t[1889], t[1888], t[1887], t[1886], t[1885], t[1884], t[1883], t[1882], t[1881], t[1880], t[1879], t[1878], t[1877], t[1876], t[1875], t[1874], t[1873], t[1872], t[1871], t[1870], t[1869], t[1868], t[1867], t[1866], t[1865], t[1864], t[1863], t[1862], t[1861], t[1860], t[1859], t[1858], t[1857], t[1856], t[1855], t[1854], t[1853], t[1852], t[1851], t[1850], t[1849], t[1848], t[1847], t[1846], t[1845], t[1844], t[1843], t[1842], t[1841], t[1840], t[1839], t[1838], t[1837], t[1836], t[1835], t[1834], t[1833], t[1832], t[1831], t[1830], t[1829], t[1828], t[1827], t[1826], t[1825], t[1824], t[1823], t[1822], t[1821], t[1820], t[1819], t[1818], t[1817], t[1816], t[1815], t[1814], t[1813], t[1812], t[1811], t[1810], t[1809], t[1808], t[1807], t[1806], t[1805], t[1804], t[1803], t[1802], t[1801], t[1800], t[1799], t[1798], t[1797], t[1796], t[1795], t[1794], t[1793], t[1792], t[1791], t[1790], t[1789], t[1788], t[1787], t[1786], t[1785], t[1784], t[1783], t[1782], t[1781], t[1780], t[1779], t[1778], t[1777], t[1776], t[1775], t[1774], t[1773], t[1772], t[1771], t[1770], t[1769], t[1768], t[1767], t[1766], t[1765], t[1764], t[1763], t[1762], t[1761], t[1760], t[1759], t[1758], t[1757], t[1756], t[1755], t[1754], t[1753], t[1752], t[1751], t[1750], t[1749], t[1748], t[1747], t[1746], t[1745], t[1744], t[1743], t[1742], t[1741], t[1740], t[1739], t[1738], t[1737], t[1736], t[1735], t[1734], t[1733], t[1732], t[1731], t[1730], t[1729], t[1728], t[1727], t[1726], t[1725], t[1724], t[1723], t[1722], t[1721], t[1720], t[1719], t[1718], t[1717], t[1716], t[1715], t[1714], t[1713], t[1712], t[1711], t[1710], t[1709], t[1708], t[1707], t[1706], t[1705], t[1704], t[1703], t[1702], t[1701], t[1700], t[1699], t[1698], t[1697], t[1696], t[1695], t[1694], t[1693], t[1692], t[1691], t[1690], t[1689], t[1688], t[1687], t[1686], t[1685], t[1684], t[1683], t[1682], t[1681], t[1680], t[1679], t[1678], t[1677], t[1676], t[1675], t[1674], t[1673], t[1672], t[1671], t[1670], t[1669], t[1668], t[1667], t[1666], t[1665], t[1664], t[1663], t[1662], t[1661], t[1660], t[1659], t[1658], t[1657], t[1656], t[1655], t[1654], t[1653], t[1652], t[1651], t[1650], t[1649], t[1648], t[1647], t[1646], t[1645], t[1644], t[1643], t[1642], t[1641], t[1640], t[1639], t[1638], t[1637], t[1636], t[1635], t[1634], t[1633], t[1632], t[1631], t[1630], t[1629], t[1628], t[1627], t[1626], t[1625], t[1624], t[1623], t[1622], t[1621], t[1620], t[1619], t[1618], t[1617], t[1616], t[1615], t[1614], t[1613], t[1612], t[1611], t[1610], t[1609], t[1608], t[1607], t[1606], t[1605], t[1604], t[1603], t[1602], t[1601], t[1600], t[1599], t[1598], t[1597], t[1596], t[1595], t[1594], t[1593], t[1592], t[1591], t[1590], t[1589], t[1588], t[1587], t[1586], t[1585], t[1584], t[1583], t[1582], t[1581], t[1580], t[1579], t[1578], t[1577], t[1576], t[1575], t[1574], t[1573], t[1572], t[1571], t[1570], t[1569], t[1568], t[1567], t[1566], t[1565], t[1564], t[1563], t[1562], t[1561], t[1560], t[1559], t[1558], t[1557], t[1556], t[1555], t[1554], t[1553], t[1552], t[1551], t[1550], t[1549], t[1548], t[1547], t[1546], t[1545], t[1544], t[1543], t[1542], t[1541], t[1540], t[1539], t[1538], t[1537], t[1536], t[1535], t[1534], t[1533], t[1532], t[1531], t[1530], t[1529], t[1528], t[1527], t[1526], t[1525], t[1524], t[1523], t[1522], t[1521], t[1520], t[1519], t[1518], t[1517], t[1516], t[1515], t[1514], t[1513], t[1512], t[1511], t[1510], t[1509], t[1508], t[1507], t[1506], t[1505], t[1504], t[1503], t[1502], t[1501], t[1500], t[1499], t[1498], t[1497], t[1496], t[1495], t[1494], t[1493], t[1492], t[1491], t[1490], t[1489], t[1488], t[1487], t[1486], t[1485], t[1484], t[1483], t[1482], t[1481], t[1480], t[1479], t[1478], t[1477], t[1476], t[1475], t[1474], t[1473], t[1472], t[1471], t[1470], t[1469], t[1468], t[1467], t[1466], t[1465], t[1464], t[1463], t[1462], t[1461], t[1460], t[1459], t[1458], t[1457], t[1456], t[1455], t[1454], t[1453], t[1452], t[1451], t[1450], t[1449], t[1448], t[1447], t[1446], t[1445], t[1444], t[1443], t[1442], t[1441], t[1440], t[1439], t[1438], t[1437], t[1436], t[1435], t[1434], t[1433], t[1432], t[1431], t[1430], t[1429], t[1428], t[1427], t[1426], t[1425], t[1424], t[1423], t[1422], t[1421], t[1420], t[1419], t[1418], t[1417], t[1416], t[1415], t[1414], t[1413], t[1412], t[1411], t[1410], t[1409], t[1408], t[1407], t[1406], t[1405], t[1404], t[1403], t[1402], t[1401], t[1400], t[1399], t[1398], t[1397], t[1396], t[1395], t[1394], t[1393], t[1392], t[1391], t[1390], t[1389], t[1388], t[1387], t[1386], t[1385], t[1384], t[1383], t[1382], t[1381], t[1380], t[1379], t[1378], t[1377], t[1376], t[1375], t[1374], t[1373], t[1372], t[1371], t[1370], t[1369], t[1368], t[1367], t[1366], t[1365], t[1364], t[1363], t[1362], t[1361], t[1360], t[1359], t[1358], t[1357], t[1356], t[1355]}));
  R1_ind R1_ind_inst(.x({x[184], x[120], x[183], x[119], x[182], x[118], x[181], x[117], x[180], x[116], x[179], x[115], x[178], x[114], x[177], x[113], x[176], x[112], x[168], x[104], x[167], x[103], x[166], x[102], x[165], x[101], x[164], x[100], x[163], x[99], x[162], x[98], x[161], x[97], x[160], x[96], x[152], x[88], x[151], x[87], x[150], x[86], x[149], x[85], x[148], x[84], x[147], x[83], x[146], x[82], x[145], x[81], x[144], x[80], x[136], x[72], x[135], x[71], x[134], x[70], x[133], x[69], x[132], x[68], x[131], x[67], x[130], x[66], x[129], x[65], x[128], x[64], x[191], x[127], x[190], x[126], x[189], x[125], x[188], x[124], x[187], x[123], x[186], x[122], x[185], x[121], t[430], t[1702], t[1701], t[1700], t[1699], t[435], t[1706], t[1705], t[1704], t[1703], t[440], t[1710], t[1709], t[1708], t[1707], t[445], t[1714], t[1713], t[1712], t[1711], t[450], t[1718], t[1717], t[1716], t[1715], t[455], t[1722], t[1721], t[1720], t[1719], t[460], t[1726], t[1725], t[1724], t[1723], t[465], t[1730], t[1729], t[1728], t[1727], t[470], t[1734], t[1733], t[1732], t[1731], x[175], x[111], x[174], x[110], x[173], x[109], x[172], x[108], x[171], x[107], x[170], x[106], x[169], x[105], t[510], t[1766], t[1765], t[1764], t[1763], t[515], t[1770], t[1769], t[1768], t[1767], t[520], t[1774], t[1773], t[1772], t[1771], t[525], t[1778], t[1777], t[1776], t[1775], t[530], t[1782], t[1781], t[1780], t[1779], t[535], t[1786], t[1785], t[1784], t[1783], t[540], t[1790], t[1789], t[1788], t[1787], t[545], t[1794], t[1793], t[1792], t[1791], t[550], t[1798], t[1797], t[1796], t[1795], x[159], x[95], x[158], x[94], x[157], x[93], x[156], x[92], x[155], x[91], x[154], x[90], x[153], x[89], t[590], t[1830], t[1829], t[1828], t[1827], t[595], t[1834], t[1833], t[1832], t[1831], t[600], t[1838], t[1837], t[1836], t[1835], t[605], t[1842], t[1841], t[1840], t[1839], t[610], t[1846], t[1845], t[1844], t[1843], t[615], t[1850], t[1849], t[1848], t[1847], t[620], t[1854], t[1853], t[1852], t[1851], t[625], t[1858], t[1857], t[1856], t[1855], t[630], t[1862], t[1861], t[1860], t[1859], x[143], x[79], x[142], x[78], x[141], x[77], t[715], t[1930], t[1929], t[1928], t[1927], t[725], t[1938], t[1937], t[1936], t[1935], t[720], t[1934], t[1933], t[1932], t[1931], t[730], t[1942], t[1941], t[1940], t[1939], t[820], t[2014], t[2013], t[2012], t[2011], t[825], t[2018], t[2017], t[2016], t[2015], t[815], t[2010], t[2009], t[2008], t[2007], x[140], x[76], x[139], x[75], x[138], x[74], x[137], x[73], t[735], t[1946], t[1945], t[1944], t[1943], t[745], t[1954], t[1953], t[1952], t[1951], t[740], t[1950], t[1949], t[1948], t[1947], t[955], t[2122], t[2121], t[2120], t[2119], t[965], t[2130], t[2129], t[2128], t[2127], t[960], t[2126], t[2125], t[2124], t[2123], t[970], t[2134], t[2133], t[2132], t[2131], t[670], t[1894], t[1893], t[1892], t[1891], t[675], t[1898], t[1897], t[1896], t[1895], t[680], t[1902], t[1901], t[1900], t[1899], t[685], t[1906], t[1905], t[1904], t[1903], t[890], t[2070], t[2069], t[2068], t[2067], t[885], t[2066], t[2065], t[2064], t[2063], t[875], t[2058], t[2057], t[2056], t[2055], t[880], t[2062], t[2061], t[2060], t[2059], t[975], t[2138], t[2137], t[2136], t[2135], t[985], t[2146], t[2145], t[2144], t[2143], t[980], t[2142], t[2141], t[2140], t[2139], t[690], t[1910], t[1909], t[1908], t[1907], t[695], t[1914], t[1913], t[1912], t[1911], t[700], t[1918], t[1917], t[1916], t[1915], t[705], t[1922], t[1921], t[1920], t[1919], t[905], t[2082], t[2081], t[2080], t[2079], t[895], t[2074], t[2073], t[2072], t[2071], t[900], t[2078], t[2077], t[2076], t[2075], t[800], t[1998], t[1997], t[1996], t[1995], t[805], t[2002], t[2001], t[2000], t[1999], t[795], t[1994], t[1993], t[1992], t[1991], t[810], t[2006], t[2005], t[2004], t[2003], t[710], t[1926], t[1925], t[1924], t[1923], t[55], t[1402], t[1401], t[1400], t[1399], t[395], t[1674], t[1673], t[1672], t[1671], x[63], t[400], t[1678], t[1677], t[1676], t[1675], x[62], t[405], t[1682], t[1681], t[1680], t[1679], x[61], t[410], t[1686], t[1685], t[1684], t[1683], x[60], t[415], t[1690], t[1689], t[1688], t[1687], x[59], t[420], t[1694], t[1693], t[1692], t[1691], x[58], t[425], t[1698], t[1697], t[1696], t[1695], x[57], t[750], t[1958], t[1957], t[1956], t[1955], x[56], t[755], t[1962], t[1961], t[1960], t[1959], x[55], t[760], t[1966], t[1965], t[1964], t[1963], x[54], t[765], t[1970], t[1969], t[1968], t[1967], x[53], t[770], t[1974], t[1973], t[1972], t[1971], x[52], t[775], t[1978], t[1977], t[1976], t[1975], x[51], t[780], t[1982], t[1981], t[1980], t[1979], x[50], t[785], t[1986], t[1985], t[1984], t[1983], x[49], t[790], t[1990], t[1989], t[1988], t[1987], x[48], t[475], t[1738], t[1737], t[1736], t[1735], x[47], t[480], t[1742], t[1741], t[1740], t[1739], x[46], t[485], t[1746], t[1745], t[1744], t[1743], x[45], t[490], t[1750], t[1749], t[1748], t[1747], x[44], t[495], t[1754], t[1753], t[1752], t[1751], x[43], t[500], t[1758], t[1757], t[1756], t[1755], x[42], t[505], t[1762], t[1761], t[1760], t[1759], x[41], t[830], t[2022], t[2021], t[2020], t[2019], x[40], t[835], t[2026], t[2025], t[2024], t[2023], x[39], t[840], t[2030], t[2029], t[2028], t[2027], x[38], t[845], t[2034], t[2033], t[2032], t[2031], x[37], t[850], t[2038], t[2037], t[2036], t[2035], x[36], t[855], t[2042], t[2041], t[2040], t[2039], x[35], t[860], t[2046], t[2045], t[2044], t[2043], x[34], t[865], t[2050], t[2049], t[2048], t[2047], x[33], t[870], t[2054], t[2053], t[2052], t[2051], x[32], t[555], t[1802], t[1801], t[1800], t[1799], x[31], t[560], t[1806], t[1805], t[1804], t[1803], x[30], t[565], t[1810], t[1809], t[1808], t[1807], x[29], t[570], t[1814], t[1813], t[1812], t[1811], x[28], t[575], t[1818], t[1817], t[1816], t[1815], x[27], t[580], t[1822], t[1821], t[1820], t[1819], x[26], t[585], t[1826], t[1825], t[1824], t[1823], x[25], t[910], t[2086], t[2085], t[2084], t[2083], x[24], t[915], t[2090], t[2089], t[2088], t[2087], x[23], t[920], t[2094], t[2093], t[2092], t[2091], x[22], t[925], t[2098], t[2097], t[2096], t[2095], x[21], t[930], t[2102], t[2101], t[2100], t[2099], x[20], t[935], t[2106], t[2105], t[2104], t[2103], x[19], t[940], t[2110], t[2109], t[2108], t[2107], x[18], t[945], t[2114], t[2113], t[2112], t[2111], x[17], t[950], t[2118], t[2117], t[2116], t[2115], x[16], t[635], t[1866], t[1865], t[1864], t[1863], x[15], t[640], t[1870], t[1869], t[1868], t[1867], x[14], t[1035], t[2186], t[2185], t[2184], t[2183], t[645], t[1874], t[1873], t[1872], t[1871], x[13], t[1335], t[2426], t[2425], t[2424], t[2423], t[1350], t[2438], t[2437], t[2436], t[2435], t[1250], t[2358], t[2357], t[2356], t[2355], t[1235], t[2346], t[2345], t[2344], t[2343], t[1240], t[2350], t[2349], t[2348], t[2347], t[1145], t[2274], t[2273], t[2272], t[2271], t[1050], t[2198], t[2197], t[2196], t[2195], t[1140], t[2270], t[2269], t[2268], t[2267], t[1245], t[2354], t[2353], t[2352], t[2351], t[1150], t[2278], t[2277], t[2276], t[2275], t[1045], t[2194], t[2193], t[2192], t[2191], t[1040], t[2190], t[2189], t[2188], t[2187], t[1135], t[2266], t[2265], t[2264], t[2263], t[1345], t[2434], t[2433], t[2432], t[2431], t[1340], t[2430], t[2429], t[2428], t[2427], t[650], t[1878], t[1877], t[1876], t[1875], x[12], t[655], t[1882], t[1881], t[1880], t[1879], x[11], t[660], t[1886], t[1885], t[1884], t[1883], x[10], t[35], t[1386], t[1385], t[1384], t[1383], t[40], t[1390], t[1389], t[1388], t[1387], t[45], t[1394], t[1393], t[1392], t[1391], t[50], t[1398], t[1397], t[1396], t[1395], t[1055], t[2202], t[2201], t[2200], t[2199], t[665], t[1890], t[1889], t[1888], t[1887], x[9], t[1275], t[2378], t[2377], t[2376], t[2375], t[1290], t[2390], t[2389], t[2388], t[2387], t[1270], t[2374], t[2373], t[2372], t[2371], t[1255], t[2362], t[2361], t[2360], t[2359], t[1260], t[2366], t[2365], t[2364], t[2363], t[1165], t[2290], t[2289], t[2288], t[2287], t[1070], t[2214], t[2213], t[2212], t[2211], t[1160], t[2286], t[2285], t[2284], t[2283], t[1265], t[2370], t[2369], t[2368], t[2367], t[1170], t[2294], t[2293], t[2292], t[2291], t[1065], t[2210], t[2209], t[2208], t[2207], t[1060], t[2206], t[2205], t[2204], t[2203], t[1155], t[2282], t[2281], t[2280], t[2279], t[1285], t[2386], t[2385], t[2384], t[2383], t[1280], t[2382], t[2381], t[2380], t[2379], t[990], t[2150], t[2149], t[2148], t[2147], x[8], t[995], t[2154], t[2153], t[2152], t[2151], x[7], t[1000], t[2158], t[2157], t[2156], t[2155], x[6], t[1075], t[2218], t[2217], t[2216], t[2215], t[1005], t[2162], t[2161], t[2160], t[2159], x[5], t[1295], t[2394], t[2393], t[2392], t[2391], t[1310], t[2406], t[2405], t[2404], t[2403], t[1210], t[2326], t[2325], t[2324], t[2323], t[1195], t[2314], t[2313], t[2312], t[2311], t[1200], t[2318], t[2317], t[2316], t[2315], t[1185], t[2306], t[2305], t[2304], t[2303], t[1090], t[2230], t[2229], t[2228], t[2227], t[1180], t[2302], t[2301], t[2300], t[2299], t[1205], t[2322], t[2321], t[2320], t[2319], t[1190], t[2310], t[2309], t[2308], t[2307], t[1085], t[2226], t[2225], t[2224], t[2223], t[1080], t[2222], t[2221], t[2220], t[2219], t[1175], t[2298], t[2297], t[2296], t[2295], t[1305], t[2402], t[2401], t[2400], t[2399], t[1300], t[2398], t[2397], t[2396], t[2395], t[1010], t[2166], t[2165], t[2164], t[2163], x[4], t[1015], t[2170], t[2169], t[2168], t[2167], t[65], t[1410], t[1409], t[1408], t[1407], x[3], t[1020], t[2174], t[2173], t[2172], t[2171], t[70], t[1414], t[1413], t[1412], t[1411], x[2], t[1095], t[2234], t[2233], t[2232], t[2231], t[1025], t[2178], t[2177], t[2176], t[2175], x[1], t[1315], t[2410], t[2409], t[2408], t[2407], t[1330], t[2422], t[2421], t[2420], t[2419], t[1230], t[2342], t[2341], t[2340], t[2339], t[1215], t[2330], t[2329], t[2328], t[2327], t[1220], t[2334], t[2333], t[2332], t[2331], t[1125], t[2258], t[2257], t[2256], t[2255], t[1110], t[2246], t[2245], t[2244], t[2243], t[1120], t[2254], t[2253], t[2252], t[2251], t[1225], t[2338], t[2337], t[2336], t[2335], t[1130], t[2262], t[2261], t[2260], t[2259], t[1105], t[2242], t[2241], t[2240], t[2239], t[1100], t[2238], t[2237], t[2236], t[2235], t[1115], t[2250], t[2249], t[2248], t[2247], t[1325], t[2418], t[2417], t[2416], t[2415], t[1320], t[2414], t[2413], t[2412], t[2411], t[1030], t[2182], t[2181], t[2180], t[2179], t[60], t[1406], t[1405], t[1404], t[1403], x[0], t[10], t[1366], t[1365], t[1364], t[1363], t[25], t[1378], t[1377], t[1376], t[1375], t[5], t[1362], t[1361], t[1360], t[1359], t[30], t[1382], t[1381], t[1380], t[1379], t[20], t[1374], t[1373], t[1372], t[1371], t[15], t[1370], t[1369], t[1368], t[1367], x[192], t[390], t[1670], t[1669], t[1668], t[1667], t[385], t[1666], t[1665], t[1664], t[1663], t[380], t[1662], t[1661], t[1660], t[1659], t[375], t[1658], t[1657], t[1656], t[1655], t[370], t[1654], t[1653], t[1652], t[1651], t[365], t[1650], t[1649], t[1648], t[1647], t[360], t[1646], t[1645], t[1644], t[1643], t[355], t[1642], t[1641], t[1640], t[1639], t[350], t[1638], t[1637], t[1636], t[1635], t[345], t[1634], t[1633], t[1632], t[1631], t[340], t[1630], t[1629], t[1628], t[1627], t[335], t[1626], t[1625], t[1624], t[1623], t[330], t[1622], t[1621], t[1620], t[1619], t[325], t[1618], t[1617], t[1616], t[1615], t[320], t[1614], t[1613], t[1612], t[1611], t[315], t[1610], t[1609], t[1608], t[1607], t[310], t[1606], t[1605], t[1604], t[1603], t[305], t[1602], t[1601], t[1600], t[1599], t[300], t[1598], t[1597], t[1596], t[1595], t[295], t[1594], t[1593], t[1592], t[1591], t[290], t[1590], t[1589], t[1588], t[1587], t[285], t[1586], t[1585], t[1584], t[1583], t[280], t[1582], t[1581], t[1580], t[1579], t[275], t[1578], t[1577], t[1576], t[1575], t[270], t[1574], t[1573], t[1572], t[1571], t[265], t[1570], t[1569], t[1568], t[1567], t[260], t[1566], t[1565], t[1564], t[1563], t[255], t[1562], t[1561], t[1560], t[1559], t[250], t[1558], t[1557], t[1556], t[1555], t[245], t[1554], t[1553], t[1552], t[1551], t[240], t[1550], t[1549], t[1548], t[1547], t[235], t[1546], t[1545], t[1544], t[1543], t[230], t[1542], t[1541], t[1540], t[1539], t[225], t[1538], t[1537], t[1536], t[1535], t[220], t[1534], t[1533], t[1532], t[1531], t[215], t[1530], t[1529], t[1528], t[1527], t[210], t[1526], t[1525], t[1524], t[1523], t[205], t[1522], t[1521], t[1520], t[1519], t[200], t[1518], t[1517], t[1516], t[1515], t[195], t[1514], t[1513], t[1512], t[1511], t[190], t[1510], t[1509], t[1508], t[1507], t[185], t[1506], t[1505], t[1504], t[1503], t[180], t[1502], t[1501], t[1500], t[1499], t[175], t[1498], t[1497], t[1496], t[1495], t[170], t[1494], t[1493], t[1492], t[1491], t[165], t[1490], t[1489], t[1488], t[1487], t[160], t[1486], t[1485], t[1484], t[1483], t[155], t[1482], t[1481], t[1480], t[1479], t[150], t[1478], t[1477], t[1476], t[1475], t[145], t[1474], t[1473], t[1472], t[1471], t[140], t[1470], t[1469], t[1468], t[1467], t[135], t[1466], t[1465], t[1464], t[1463], t[130], t[1462], t[1461], t[1460], t[1459], t[125], t[1458], t[1457], t[1456], t[1455], t[120], t[1454], t[1453], t[1452], t[1451], t[115], t[1450], t[1449], t[1448], t[1447], t[110], t[1446], t[1445], t[1444], t[1443], t[105], t[1442], t[1441], t[1440], t[1439], t[100], t[1438], t[1437], t[1436], t[1435], t[95], t[1434], t[1433], t[1432], t[1431], t[90], t[1430], t[1429], t[1428], t[1427], t[85], t[1426], t[1425], t[1424], t[1423], t[80], t[1422], t[1421], t[1420], t[1419], t[75], t[1418], t[1417], t[1416], t[1415], t[0], t[1358], t[1357], t[1356], t[1355]}), .y({t[2774], t[2773], t[2772], t[2771], t[2770], t[2769], t[2768], t[2767], t[2766], t[2765], t[2764], t[2763], t[2762], t[2761], t[2760], t[2759], t[2758], t[2757], t[2756], t[2755], t[2754], t[2753], t[2752], t[2751], t[2750], t[2749], t[2748], t[2747], t[2746], t[2745], t[2744], t[2743], t[2742], t[2741], t[2740], t[2739], t[2738], t[2737], t[2736], t[2735], t[2734], t[2733], t[2732], t[2731], t[2730], t[2729], t[2728], t[2727], t[2726], t[2725], t[2724], t[2723], t[2722], t[2721], t[2720], t[2719], t[2718], t[2717], t[2716], t[2715], t[2714], t[2713], t[2712], t[2711], t[2710], t[2709], t[2708], t[2707], t[2706], t[2705], t[2704], t[2703], t[2702], t[2701], t[2700], t[2699], t[2698], t[2697], t[2696], t[2695], t[2694], t[2693], t[2692], t[2691], t[2690], t[2689], t[2688], t[2687], t[2686], t[2685], t[2684], t[2683], t[2682], t[2681], t[2680], t[2679], t[2678], t[2677], t[2676], t[2675], t[2674], t[2673], t[2672], t[2671], t[2670], t[2669], t[2668], t[2667], t[2666], t[2665], t[2664], t[2663], t[2662], t[2661], t[2660], t[2659], t[2658], t[2657], t[2656], t[2655], t[2654], t[2653], t[2652], t[2651], t[2650], t[2649], t[2648], t[2647], t[2646], t[2645], t[2644], t[2643], t[2642], t[2641], t[2640], t[2639], t[2638], t[2637], t[2636], t[2635], t[2634], t[2633], t[2632], t[2631], t[2630], t[2629], t[2628], t[2627], t[2626], t[2625], t[2624], t[2623], t[2622], t[2621], t[2620], t[2619], t[2618], t[2617], t[2616], t[2615], t[2614], t[2613], t[2612], t[2611], t[2610], t[2609], t[2608], t[2607], t[2606], t[2605], t[2604], t[2603], t[2602], t[2601], t[2600], t[2599], t[2598], t[2597], t[2596], t[2595], t[2594], t[2593], t[2592], t[2591], t[2590], t[2589], t[2588], t[2587], t[2586], t[2585], t[2584], t[2583], t[2582], t[2581], t[2580], t[2579], t[2578], t[2577], t[2576], t[2575], t[2574], t[2573], t[2572], t[2571], t[2570], t[2569], t[2568], t[2567], t[2566], t[2565], t[2564], t[2563], t[2562], t[2561], t[2560], t[2559], t[2558], t[2557], t[2556], t[2555], t[2554], t[2553], t[2552], t[2551], t[2550], t[2549], t[2548], t[2547], t[2546], t[2545], t[2544], t[2543], t[2542], t[2541], t[2540], t[2539], t[2538], t[2537], t[2536], t[2535], t[2534], t[2533], t[2532], t[2531], t[2530], t[2529], t[2528], t[2527], t[2526], t[2525], t[2524], t[2523], t[2522], t[2521], t[2520], t[2519], t[2518], t[2517], t[2516], t[2515], t[2514], t[2513], t[2512], t[2511], t[2510], t[2509], t[2508], t[2507], t[2506], t[2505], t[2504], t[2503], t[2502], t[2501], t[2500], t[2499], t[2498], t[2497], t[2496], t[2495], t[2494], t[2493], t[2492], t[2491], t[2490], t[2489], t[2488], t[2487], t[2486], t[2485], t[2484], t[2483], t[2482], t[2481], t[2480], t[2479], t[2478], t[2477], t[2476], t[2475], t[2474], t[2473], t[2472], t[2471], t[2470], t[2469], t[2468], t[2467], t[2466], t[2465], t[2464], t[2463], t[2462], t[2461], t[2460], t[2459], t[2458], t[2457], t[2456], t[2455], t[2454], t[2453], t[2452], t[2451], t[2450], t[2449], t[2448], t[2447], t[2446], t[2445], t[2444], t[2443], t[2442], t[2441], t[2440], t[2439]}));
  R2_ind R2_ind_inst(.x({t[981], t[984], t[983], t[982], t[980], t[986], t[989], t[988], t[987], t[985], t[976], t[979], t[978], t[977], t[975], t[961], t[964], t[963], t[962], t[960], t[966], t[969], t[968], t[967], t[965], t[956], t[959], t[958], t[957], t[955], t[971], t[974], t[973], t[972], t[970], t[901], t[904], t[903], t[902], t[900], t[906], t[909], t[908], t[907], t[905], t[896], t[899], t[898], t[897], t[895], t[881], t[884], t[883], t[882], t[880], t[886], t[889], t[888], t[887], t[885], t[876], t[879], t[878], t[877], t[875], t[891], t[894], t[893], t[892], t[890], t[821], t[824], t[823], t[822], t[820], t[826], t[829], t[828], t[827], t[825], t[816], t[819], t[818], t[817], t[815], t[801], t[804], t[803], t[802], t[800], t[806], t[809], t[808], t[807], t[805], t[796], t[799], t[798], t[797], t[795], t[811], t[814], t[813], t[812], t[810], t[741], t[744], t[743], t[742], t[740], t[746], t[749], t[748], t[747], t[745], t[736], t[739], t[738], t[737], t[735], t[721], t[724], t[723], t[722], t[720], t[726], t[729], t[728], t[727], t[725], t[716], t[719], t[718], t[717], t[715], t[731], t[734], t[733], t[732], t[730], t[711], t[714], t[713], t[712], t[710], t[706], t[709], t[708], t[707], t[705], t[701], t[704], t[703], t[702], t[700], t[696], t[699], t[698], t[697], t[695], t[691], t[694], t[693], t[692], t[690], t[686], t[689], t[688], t[687], t[685], t[681], t[684], t[683], t[682], t[680], t[676], t[679], t[678], t[677], t[675], t[671], t[674], t[673], t[672], t[670], t[631], t[634], t[633], t[632], t[630], t[626], t[629], t[628], t[627], t[625], t[621], t[624], t[623], t[622], t[620], t[616], t[619], t[618], t[617], t[615], t[611], t[614], t[613], t[612], t[610], t[606], t[609], t[608], t[607], t[605], t[601], t[604], t[603], t[602], t[600], t[596], t[599], t[598], t[597], t[595], t[591], t[594], t[593], t[592], t[590], t[551], t[554], t[553], t[552], t[550], t[546], t[549], t[548], t[547], t[545], t[541], t[544], t[543], t[542], t[540], t[536], t[539], t[538], t[537], t[535], t[531], t[534], t[533], t[532], t[530], t[526], t[529], t[528], t[527], t[525], t[521], t[524], t[523], t[522], t[520], t[516], t[519], t[518], t[517], t[515], t[511], t[514], t[513], t[512], t[510], t[471], t[474], t[473], t[472], t[470], t[466], t[469], t[468], t[467], t[465], t[461], t[464], t[463], t[462], t[460], t[456], t[459], t[458], t[457], t[455], t[451], t[454], t[453], t[452], t[450], t[446], t[449], t[448], t[447], t[445], t[441], t[444], t[443], t[442], t[440], t[436], t[439], t[438], t[437], t[435], t[431], t[434], t[433], t[432], t[430], x[128], x[64], t[391], t[394], t[393], t[392], t[390], x[129], x[65], t[386], t[389], t[388], t[387], t[385], x[130], x[66], t[381], t[384], t[383], t[382], t[380], x[131], x[67], t[376], t[379], t[378], t[377], t[375], x[132], x[68], t[371], t[374], t[373], t[372], t[370], x[133], x[69], t[366], t[369], t[368], t[367], t[365], x[134], x[70], t[361], t[364], t[363], t[362], t[360], x[135], x[71], t[356], t[359], t[358], t[357], t[355], x[136], x[72], t[351], t[354], t[353], t[352], t[350], x[137], x[73], x[138], x[74], x[139], x[75], x[140], x[76], x[141], x[77], x[142], x[78], x[143], x[79], x[144], x[80], t[311], t[314], t[313], t[312], t[310], x[145], x[81], t[306], t[309], t[308], t[307], t[305], x[146], x[82], t[301], t[304], t[303], t[302], t[300], x[147], x[83], t[296], t[299], t[298], t[297], t[295], x[148], x[84], t[291], t[294], t[293], t[292], t[290], x[149], x[85], t[286], t[289], t[288], t[287], t[285], x[150], x[86], t[281], t[284], t[283], t[282], t[280], x[151], x[87], t[276], t[279], t[278], t[277], t[275], x[152], x[88], t[271], t[274], t[273], t[272], t[270], x[153], x[89], x[154], x[90], x[155], x[91], x[156], x[92], x[157], x[93], x[158], x[94], x[159], x[95], x[160], x[96], t[231], t[234], t[233], t[232], t[230], x[161], x[97], t[226], t[229], t[228], t[227], t[225], x[162], x[98], t[221], t[224], t[223], t[222], t[220], x[163], x[99], t[216], t[219], t[218], t[217], t[215], x[164], x[100], t[211], t[214], t[213], t[212], t[210], x[165], x[101], t[206], t[209], t[208], t[207], t[205], x[166], x[102], t[201], t[204], t[203], t[202], t[200], x[167], x[103], t[196], t[199], t[198], t[197], t[195], x[168], x[104], t[191], t[194], t[193], t[192], t[190], x[169], x[105], x[170], x[106], x[171], x[107], x[172], x[108], x[173], x[109], x[174], x[110], x[175], x[111], x[176], x[112], t[151], t[154], t[153], t[152], t[150], x[177], x[113], t[146], t[149], t[148], t[147], t[145], x[178], x[114], t[141], t[144], t[143], t[142], t[140], x[179], x[115], t[136], t[139], t[138], t[137], t[135], x[180], x[116], t[131], t[134], t[133], t[132], t[130], x[181], x[117], t[126], t[129], t[128], t[127], t[125], x[182], x[118], t[121], t[124], t[123], t[122], t[120], x[183], x[119], t[116], t[119], t[118], t[117], t[115], x[184], x[120], t[111], t[114], t[113], t[112], t[110], x[185], x[121], x[186], x[122], x[187], x[123], x[188], x[124], x[189], x[125], x[190], x[126], x[191], x[127], t[1031], t[1034], t[1033], t[1032], t[1030], x[0], t[1026], t[1029], t[1028], t[1027], t[1025], x[1], t[1021], t[1024], t[1023], t[1022], t[1020], x[2], t[1016], t[1019], t[1018], t[1017], t[1015], x[3], t[1011], t[1014], t[1013], t[1012], t[1010], x[4], t[1006], t[1009], t[1008], t[1007], t[1005], x[5], t[1001], t[1004], t[1003], t[1002], t[1000], x[6], t[996], t[999], t[998], t[997], t[995], x[7], t[991], t[994], t[993], t[992], t[990], x[8], t[666], t[669], t[668], t[667], t[665], t[346], t[349], t[348], t[347], t[345], x[9], t[661], t[664], t[663], t[662], t[660], t[341], t[344], t[343], t[342], t[340], x[10], t[656], t[659], t[658], t[657], t[655], t[336], t[339], t[338], t[337], t[335], x[11], t[651], t[654], t[653], t[652], t[650], t[331], t[334], t[333], t[332], t[330], x[12], t[646], t[649], t[648], t[647], t[645], t[326], t[329], t[328], t[327], t[325], x[13], t[641], t[644], t[643], t[642], t[640], t[321], t[324], t[323], t[322], t[320], x[14], t[636], t[639], t[638], t[637], t[635], t[316], t[319], t[318], t[317], t[315], x[15], t[951], t[954], t[953], t[952], t[950], x[16], t[946], t[949], t[948], t[947], t[945], x[17], t[941], t[944], t[943], t[942], t[940], x[18], t[936], t[939], t[938], t[937], t[935], x[19], t[931], t[934], t[933], t[932], t[930], x[20], t[926], t[929], t[928], t[927], t[925], x[21], t[921], t[924], t[923], t[922], t[920], x[22], t[916], t[919], t[918], t[917], t[915], x[23], t[911], t[914], t[913], t[912], t[910], x[24], t[586], t[589], t[588], t[587], t[585], t[266], t[269], t[268], t[267], t[265], x[25], t[581], t[584], t[583], t[582], t[580], t[261], t[264], t[263], t[262], t[260], x[26], t[576], t[579], t[578], t[577], t[575], t[256], t[259], t[258], t[257], t[255], x[27], t[571], t[574], t[573], t[572], t[570], t[251], t[254], t[253], t[252], t[250], x[28], t[566], t[569], t[568], t[567], t[565], t[246], t[249], t[248], t[247], t[245], x[29], t[561], t[564], t[563], t[562], t[560], t[241], t[244], t[243], t[242], t[240], x[30], t[556], t[559], t[558], t[557], t[555], t[236], t[239], t[238], t[237], t[235], x[31], t[871], t[874], t[873], t[872], t[870], x[32], t[866], t[869], t[868], t[867], t[865], x[33], t[861], t[864], t[863], t[862], t[860], x[34], t[856], t[859], t[858], t[857], t[855], x[35], t[851], t[854], t[853], t[852], t[850], x[36], t[846], t[849], t[848], t[847], t[845], x[37], t[841], t[844], t[843], t[842], t[840], x[38], t[836], t[839], t[838], t[837], t[835], x[39], t[831], t[834], t[833], t[832], t[830], x[40], t[506], t[509], t[508], t[507], t[505], t[186], t[189], t[188], t[187], t[185], x[41], t[501], t[504], t[503], t[502], t[500], t[181], t[184], t[183], t[182], t[180], x[42], t[496], t[499], t[498], t[497], t[495], t[176], t[179], t[178], t[177], t[175], x[43], t[491], t[494], t[493], t[492], t[490], t[171], t[174], t[173], t[172], t[170], x[44], t[486], t[489], t[488], t[487], t[485], t[166], t[169], t[168], t[167], t[165], x[45], t[481], t[484], t[483], t[482], t[480], t[161], t[164], t[163], t[162], t[160], x[46], t[476], t[479], t[478], t[477], t[475], t[156], t[159], t[158], t[157], t[155], x[47], t[1131], t[1134], t[1133], t[1132], t[1130], t[1226], t[1229], t[1228], t[1227], t[1225], t[1101], t[1104], t[1103], t[1102], t[1100], t[1326], t[1329], t[1328], t[1327], t[1325], t[791], t[794], t[793], t[792], t[790], x[48], t[1221], t[1224], t[1223], t[1222], t[1220], t[1126], t[1129], t[1128], t[1127], t[1125], t[1321], t[1324], t[1323], t[1322], t[1320], t[1096], t[1099], t[1098], t[1097], t[1095], t[786], t[789], t[788], t[787], t[785], x[49], t[1111], t[1114], t[1113], t[1112], t[1110], t[1121], t[1124], t[1123], t[1122], t[1120], t[1316], t[1319], t[1318], t[1317], t[1315], t[1216], t[1219], t[1218], t[1217], t[1215], t[781], t[784], t[783], t[782], t[780], x[50], t[1231], t[1234], t[1233], t[1232], t[1230], t[1331], t[1334], t[1333], t[1332], t[1330], t[1116], t[1119], t[1118], t[1117], t[1115], t[1106], t[1109], t[1108], t[1107], t[1105], t[776], t[779], t[778], t[777], t[775], x[51], t[1191], t[1194], t[1193], t[1192], t[1190], t[1206], t[1209], t[1208], t[1207], t[1205], t[1081], t[1084], t[1083], t[1082], t[1080], t[1306], t[1309], t[1308], t[1307], t[1305], t[771], t[774], t[773], t[772], t[770], x[52], t[1201], t[1204], t[1203], t[1202], t[1200], t[1186], t[1189], t[1188], t[1187], t[1185], t[1301], t[1304], t[1303], t[1302], t[1300], t[1076], t[1079], t[1078], t[1077], t[1075], t[766], t[769], t[768], t[767], t[765], x[53], t[1091], t[1094], t[1093], t[1092], t[1090], t[1181], t[1184], t[1183], t[1182], t[1180], t[1296], t[1299], t[1298], t[1297], t[1295], t[1196], t[1199], t[1198], t[1197], t[1195], t[761], t[764], t[763], t[762], t[760], x[54], t[1211], t[1214], t[1213], t[1212], t[1210], t[1311], t[1314], t[1313], t[1312], t[1310], t[1176], t[1179], t[1178], t[1177], t[1175], t[1086], t[1089], t[1088], t[1087], t[1085], t[756], t[759], t[758], t[757], t[755], x[55], t[1171], t[1174], t[1173], t[1172], t[1170], t[1266], t[1269], t[1268], t[1267], t[1265], t[1061], t[1064], t[1063], t[1062], t[1060], t[1286], t[1289], t[1288], t[1287], t[1285], t[751], t[754], t[753], t[752], t[750], x[56], t[1261], t[1264], t[1263], t[1262], t[1260], t[1166], t[1169], t[1168], t[1167], t[1165], t[1281], t[1284], t[1283], t[1282], t[1280], t[1056], t[1059], t[1058], t[1057], t[1055], t[426], t[429], t[428], t[427], t[425], t[106], t[109], t[108], t[107], t[105], x[57], t[1071], t[1074], t[1073], t[1072], t[1070], t[1161], t[1164], t[1163], t[1162], t[1160], t[1276], t[1279], t[1278], t[1277], t[1275], t[1256], t[1259], t[1258], t[1257], t[1255], t[421], t[424], t[423], t[422], t[420], t[101], t[104], t[103], t[102], t[100], x[58], t[1271], t[1274], t[1273], t[1272], t[1270], t[1291], t[1294], t[1293], t[1292], t[1290], t[1156], t[1159], t[1158], t[1157], t[1155], t[1066], t[1069], t[1068], t[1067], t[1065], t[416], t[419], t[418], t[417], t[415], t[96], t[99], t[98], t[97], t[95], x[59], t[1151], t[1154], t[1153], t[1152], t[1150], t[1246], t[1249], t[1248], t[1247], t[1245], t[1041], t[1044], t[1043], t[1042], t[1040], t[411], t[414], t[413], t[412], t[410], t[91], t[94], t[93], t[92], t[90], t[1346], t[1349], t[1348], t[1347], t[1345], t[71], t[74], t[73], t[72], t[70], x[60], t[1241], t[1244], t[1243], t[1242], t[1240], t[1146], t[1149], t[1148], t[1147], t[1145], t[1341], t[1344], t[1343], t[1342], t[1340], t[1036], t[1039], t[1038], t[1037], t[1035], t[406], t[409], t[408], t[407], t[405], t[86], t[89], t[88], t[87], t[85], t[61], t[64], t[63], t[62], t[60], x[61], t[1051], t[1054], t[1053], t[1052], t[1050], t[1141], t[1144], t[1143], t[1142], t[1140], t[1336], t[1339], t[1338], t[1337], t[1335], t[1236], t[1239], t[1238], t[1237], t[1235], t[401], t[404], t[403], t[402], t[400], t[81], t[84], t[83], t[82], t[80], x[62], t[1251], t[1254], t[1253], t[1252], t[1250], t[1351], t[1354], t[1353], t[1352], t[1350], t[1136], t[1139], t[1138], t[1137], t[1135], t[1046], t[1049], t[1048], t[1047], t[1045], t[396], t[399], t[398], t[397], t[395], t[76], t[79], t[78], t[77], t[75], t[66], t[69], t[68], t[67], t[65], x[63], t[56], t[59], t[58], t[57], t[55], t[46], t[49], t[48], t[47], t[45], t[41], t[44], t[43], t[42], t[40], t[36], t[39], t[38], t[37], t[35], t[51], t[54], t[53], t[52], t[50], t[11], t[14], t[13], t[12], t[10], t[26], t[29], t[28], t[27], t[25], t[6], t[9], t[8], t[7], t[5], t[31], t[34], t[33], t[32], t[30], t[21], t[24], t[23], t[22], t[20], t[16], t[19], t[18], t[17], t[15], x[192], t[1], t[4], t[3], t[2], t[0]}), .y({t[3862], t[3861], t[3860], t[3859], t[3858], t[3857], t[3856], t[3855], t[3854], t[3853], t[3852], t[3851], t[3850], t[3849], t[3848], t[3847], t[3846], t[3845], t[3844], t[3843], t[3842], t[3841], t[3840], t[3839], t[3838], t[3837], t[3836], t[3835], t[3834], t[3833], t[3832], t[3831], t[3830], t[3829], t[3828], t[3827], t[3826], t[3825], t[3824], t[3823], t[3822], t[3821], t[3820], t[3819], t[3818], t[3817], t[3816], t[3815], t[3814], t[3813], t[3812], t[3811], t[3810], t[3809], t[3808], t[3807], t[3806], t[3805], t[3804], t[3803], t[3802], t[3801], t[3800], t[3799], t[3798], t[3797], t[3796], t[3795], t[3794], t[3793], t[3792], t[3791], t[3790], t[3789], t[3788], t[3787], t[3786], t[3785], t[3784], t[3783], t[3782], t[3781], t[3780], t[3779], t[3778], t[3777], t[3776], t[3775], t[3774], t[3773], t[3772], t[3771], t[3770], t[3769], t[3768], t[3767], t[3766], t[3765], t[3764], t[3763], t[3762], t[3761], t[3760], t[3759], t[3758], t[3757], t[3756], t[3755], t[3754], t[3753], t[3752], t[3751], t[3750], t[3749], t[3748], t[3747], t[3746], t[3745], t[3744], t[3743], t[3742], t[3741], t[3740], t[3739], t[3738], t[3737], t[3736], t[3735], t[3734], t[3733], t[3732], t[3731], t[3730], t[3729], t[3728], t[3727], t[3726], t[3725], t[3724], t[3723], t[3722], t[3721], t[3720], t[3719], t[3718], t[3717], t[3716], t[3715], t[3714], t[3713], t[3712], t[3711], t[3710], t[3709], t[3708], t[3707], t[3706], t[3705], t[3704], t[3703], t[3702], t[3701], t[3700], t[3699], t[3698], t[3697], t[3696], t[3695], t[3694], t[3693], t[3692], t[3691], t[3690], t[3689], t[3688], t[3687], t[3686], t[3685], t[3684], t[3683], t[3682], t[3681], t[3680], t[3679], t[3678], t[3677], t[3676], t[3675], t[3674], t[3673], t[3672], t[3671], t[3670], t[3669], t[3668], t[3667], t[3666], t[3665], t[3664], t[3663], t[3662], t[3661], t[3660], t[3659], t[3658], t[3657], t[3656], t[3655], t[3654], t[3653], t[3652], t[3651], t[3650], t[3649], t[3648], t[3647], t[3646], t[3645], t[3644], t[3643], t[3642], t[3641], t[3640], t[3639], t[3638], t[3637], t[3636], t[3635], t[3634], t[3633], t[3632], t[3631], t[3630], t[3629], t[3628], t[3627], t[3626], t[3625], t[3624], t[3623], t[3622], t[3621], t[3620], t[3619], t[3618], t[3617], t[3616], t[3615], t[3614], t[3613], t[3612], t[3611], t[3610], t[3609], t[3608], t[3607], t[3606], t[3605], t[3604], t[3603], t[3602], t[3601], t[3600], t[3599], t[3598], t[3597], t[3596], t[3595], t[3594], t[3593], t[3592], t[3591], t[3590], t[3589], t[3588], t[3587], t[3586], t[3585], t[3584], t[3583], t[3582], t[3581], t[3580], t[3579], t[3578], t[3577], t[3576], t[3575], t[3574], t[3573], t[3572], t[3571], t[3570], t[3569], t[3568], t[3567], t[3566], t[3565], t[3564], t[3563], t[3562], t[3561], t[3560], t[3559], t[3558], t[3557], t[3556], t[3555], t[3554], t[3553], t[3552], t[3551], t[3550], t[3549], t[3548], t[3547], t[3546], t[3545], t[3544], t[3543], t[3542], t[3541], t[3540], t[3539], t[3538], t[3537], t[3536], t[3535], t[3534], t[3533], t[3532], t[3531], t[3530], t[3529], t[3528], t[3527], t[3526], t[3525], t[3524], t[3523], t[3522], t[3521], t[3520], t[3519], t[3518], t[3517], t[3516], t[3515], t[3514], t[3513], t[3512], t[3511], t[3510], t[3509], t[3508], t[3507], t[3506], t[3505], t[3504], t[3503], t[3502], t[3501], t[3500], t[3499], t[3498], t[3497], t[3496], t[3495], t[3494], t[3493], t[3492], t[3491], t[3490], t[3489], t[3488], t[3487], t[3486], t[3485], t[3484], t[3483], t[3482], t[3481], t[3480], t[3479], t[3478], t[3477], t[3476], t[3475], t[3474], t[3473], t[3472], t[3471], t[3470], t[3469], t[3468], t[3467], t[3466], t[3465], t[3464], t[3463], t[3462], t[3461], t[3460], t[3459], t[3458], t[3457], t[3456], t[3455], t[3454], t[3453], t[3452], t[3451], t[3450], t[3449], t[3448], t[3447], t[3446], t[3445], t[3444], t[3443], t[3442], t[3441], t[3440], t[3439], t[3438], t[3437], t[3436], t[3435], t[3434], t[3433], t[3432], t[3431], t[3430], t[3429], t[3428], t[3427], t[3426], t[3425], t[3424], t[3423], t[3422], t[3421], t[3420], t[3419], t[3418], t[3417], t[3416], t[3415], t[3414], t[3413], t[3412], t[3411], t[3410], t[3409], t[3408], t[3407], t[3406], t[3405], t[3404], t[3403], t[3402], t[3401], t[3400], t[3399], t[3398], t[3397], t[3396], t[3395], t[3394], t[3393], t[3392], t[3391], t[3390], t[3389], t[3388], t[3387], t[3386], t[3385], t[3384], t[3383], t[3382], t[3381], t[3380], t[3379], t[3378], t[3377], t[3376], t[3375], t[3374], t[3373], t[3372], t[3371], t[3370], t[3369], t[3368], t[3367], t[3366], t[3365], t[3364], t[3363], t[3362], t[3361], t[3360], t[3359], t[3358], t[3357], t[3356], t[3355], t[3354], t[3353], t[3352], t[3351], t[3350], t[3349], t[3348], t[3347], t[3346], t[3345], t[3344], t[3343], t[3342], t[3341], t[3340], t[3339], t[3338], t[3337], t[3336], t[3335], t[3334], t[3333], t[3332], t[3331], t[3330], t[3329], t[3328], t[3327], t[3326], t[3325], t[3324], t[3323], t[3322], t[3321], t[3320], t[3319], t[3318], t[3317], t[3316], t[3315], t[3314], t[3313], t[3312], t[3311], t[3310], t[3309], t[3308], t[3307], t[3306], t[3305], t[3304], t[3303], t[3302], t[3301], t[3300], t[3299], t[3298], t[3297], t[3296], t[3295], t[3294], t[3293], t[3292], t[3291], t[3290], t[3289], t[3288], t[3287], t[3286], t[3285], t[3284], t[3283], t[3282], t[3281], t[3280], t[3279], t[3278], t[3277], t[3276], t[3275], t[3274], t[3273], t[3272], t[3271], t[3270], t[3269], t[3268], t[3267], t[3266], t[3265], t[3264], t[3263], t[3262], t[3261], t[3260], t[3259], t[3258], t[3257], t[3256], t[3255], t[3254], t[3253], t[3252], t[3251], t[3250], t[3249], t[3248], t[3247], t[3246], t[3245], t[3244], t[3243], t[3242], t[3241], t[3240], t[3239], t[3238], t[3237], t[3236], t[3235], t[3234], t[3233], t[3232], t[3231], t[3230], t[3229], t[3228], t[3227], t[3226], t[3225], t[3224], t[3223], t[3222], t[3221], t[3220], t[3219], t[3218], t[3217], t[3216], t[3215], t[3214], t[3213], t[3212], t[3211], t[3210], t[3209], t[3208], t[3207], t[3206], t[3205], t[3204], t[3203], t[3202], t[3201], t[3200], t[3199], t[3198], t[3197], t[3196], t[3195], t[3194], t[3193], t[3192], t[3191], t[3190], t[3189], t[3188], t[3187], t[3186], t[3185], t[3184], t[3183], t[3182], t[3181], t[3180], t[3179], t[3178], t[3177], t[3176], t[3175], t[3174], t[3173], t[3172], t[3171], t[3170], t[3169], t[3168], t[3167], t[3166], t[3165], t[3164], t[3163], t[3162], t[3161], t[3160], t[3159], t[3158], t[3157], t[3156], t[3155], t[3154], t[3153], t[3152], t[3151], t[3150], t[3149], t[3148], t[3147], t[3146], t[3145], t[3144], t[3143], t[3142], t[3141], t[3140], t[3139], t[3138], t[3137], t[3136], t[3135], t[3134], t[3133], t[3132], t[3131], t[3130], t[3129], t[3128], t[3127], t[3126], t[3125], t[3124], t[3123], t[3122], t[3121], t[3120], t[3119], t[3118], t[3117], t[3116], t[3115], t[3114], t[3113], t[3112], t[3111], t[3110], t[3109], t[3108], t[3107], t[3106], t[3105], t[3104], t[3103], t[3102], t[3101], t[3100], t[3099], t[3098], t[3097], t[3096], t[3095], t[3094], t[3093], t[3092], t[3091], t[3090], t[3089], t[3088], t[3087], t[3086], t[3085], t[3084], t[3083], t[3082], t[3081], t[3080], t[3079], t[3078], t[3077], t[3076], t[3075], t[3074], t[3073], t[3072], t[3071], t[3070], t[3069], t[3068], t[3067], t[3066], t[3065], t[3064], t[3063], t[3062], t[3061], t[3060], t[3059], t[3058], t[3057], t[3056], t[3055], t[3054], t[3053], t[3052], t[3051], t[3050], t[3049], t[3048], t[3047], t[3046], t[3045], t[3044], t[3043], t[3042], t[3041], t[3040], t[3039], t[3038], t[3037], t[3036], t[3035], t[3034], t[3033], t[3032], t[3031], t[3030], t[3029], t[3028], t[3027], t[3026], t[3025], t[3024], t[3023], t[3022], t[3021], t[3020], t[3019], t[3018], t[3017], t[3016], t[3015], t[3014], t[3013], t[3012], t[3011], t[3010], t[3009], t[3008], t[3007], t[3006], t[3005], t[3004], t[3003], t[3002], t[3001], t[3000], t[2999], t[2998], t[2997], t[2996], t[2995], t[2994], t[2993], t[2992], t[2991], t[2990], t[2989], t[2988], t[2987], t[2986], t[2985], t[2984], t[2983], t[2982], t[2981], t[2980], t[2979], t[2978], t[2977], t[2976], t[2975], t[2974], t[2973], t[2972], t[2971], t[2970], t[2969], t[2968], t[2967], t[2966], t[2965], t[2964], t[2963], t[2962], t[2961], t[2960], t[2959], t[2958], t[2957], t[2956], t[2955], t[2954], t[2953], t[2952], t[2951], t[2950], t[2949], t[2948], t[2947], t[2946], t[2945], t[2944], t[2943], t[2942], t[2941], t[2940], t[2939], t[2938], t[2937], t[2936], t[2935], t[2934], t[2933], t[2932], t[2931], t[2930], t[2929], t[2928], t[2927], t[2926], t[2925], t[2924], t[2923], t[2922], t[2921], t[2920], t[2919], t[2918], t[2917], t[2916], t[2915], t[2914], t[2913], t[2912], t[2911], t[2910], t[2909], t[2908], t[2907], t[2906], t[2905], t[2904], t[2903], t[2902], t[2901], t[2900], t[2899], t[2898], t[2897], t[2896], t[2895], t[2894], t[2893], t[2892], t[2891], t[2890], t[2889], t[2888], t[2887], t[2886], t[2885], t[2884], t[2883], t[2882], t[2881], t[2880], t[2879], t[2878], t[2877], t[2876], t[2875], t[2874], t[2873], t[2872], t[2871], t[2870], t[2869], t[2868], t[2867], t[2866], t[2865], t[2864], t[2863], t[2862], t[2861], t[2860], t[2859], t[2858], t[2857], t[2856], t[2855], t[2854], t[2853], t[2852], t[2851], t[2850], t[2849], t[2848], t[2847], t[2846], t[2845], t[2844], t[2843], t[2842], t[2841], t[2840], t[2839], t[2838], t[2837], t[2836], t[2835], t[2834], t[2833], t[2832], t[2831], t[2830], t[2829], t[2828], t[2827], t[2826], t[2825], t[2824], t[2823], t[2822], t[2821], t[2820], t[2819], t[2818], t[2817], t[2816], t[2815], t[2814], t[2813], t[2812], t[2811], t[2810], t[2809], t[2808], t[2807], t[2806], t[2805], t[2804], t[2803], t[2802], t[2801], t[2800], t[2799], t[2798], t[2797], t[2796], t[2795], t[2794], t[2793], t[2792], t[2791], t[2790], t[2789], t[2788], t[2787], t[2786], t[2785], t[2784], t[2783], t[2782], t[2781], t[2780], t[2779], t[2778], t[2777], t[2776], t[2775]}));
  Reg1 Reg1_inst(.x({t[2504], t[2606], t[2619], t[2631], t[2627], t[2656], t[2644], t[2643], t[2657], t[2626], t[2594], t[2582], t[2581], t[2595], t[2616], t[2604], t[2603], t[2617], t[2636], t[2624], t[2639], t[2623], t[2637], t[2635], t[2629], t[2633], t[2634], t[2655], t[2649], t[2653], t[2654], t[2651], t[2593], t[2587], t[2591], t[2592], t[2615], t[2609], t[2613], t[2614], t[2608], t[2612], t[2647], t[2610], t[2605], t[2628], t[2632], t[2630], t[2625], t[2648], t[2652], t[2650], t[2645], t[2646], t[2586], t[2590], t[2588], t[2583], t[2589], t[2585], t[2584], t[2597], t[2611], t[2607], t[2659], t[2559], t[2560], t[2561], t[2562], t[2505], t[2506], t[2507], t[2508], t[2563], t[2509], t[2510], t[2511], t[2512], t[2513], t[2514], t[2515], t[2516], t[2517], t[2518], t[2564], t[2519], t[2520], t[2521], t[2522], t[2523], t[2524], t[2525], t[2526], t[2527], t[2528], t[2565], t[2529], t[2530], t[2531], t[2532], t[2533], t[2534], t[2535], t[2536], t[2537], t[2538], t[2566], t[2539], t[2540], t[2541], t[2542], t[2543], t[2544], t[2545], t[2546], t[2547], t[2548], t[2567], t[2549], t[2550], t[2551], t[2552], t[2553], t[2554], t[2555], t[2556], t[2557], t[2558], t[2568], t[2772], t[2773], t[2774], t[2703], t[2711], t[2719], t[2720], t[2721], t[2704], t[2722], t[2730], t[2731], t[2732], t[2733], t[2638], t[2640], t[2641], t[2642], t[2658], t[2705], t[2660], t[2661], t[2748], t[2749], t[2750], t[2751], t[2752], t[2753], t[2754], t[2755], t[2706], t[2756], t[2671], t[2672], t[2673], t[2674], t[2675], t[2676], t[2677], t[2757], t[2758], t[2707], t[2759], t[2760], t[2761], t[2762], t[2763], t[2764], t[2765], t[2687], t[2688], t[2689], t[2708], t[2690], t[2691], t[2692], t[2693], t[2766], t[2767], t[2768], t[2769], t[2770], t[2771], t[2709], t[2700], t[2701], t[2702], t[2739], t[2580], t[2596], t[2599], t[2601], t[2738], t[2602], t[2618], t[2620], t[2621], t[2622], t[2724], t[2723], t[2725], t[2734], t[2736], t[2740], t[2735], t[2737], t[2662], t[2663], t[2664], t[2665], t[2666], t[2667], t[2668], t[2669], t[2744], t[2670], t[2718], t[2716], t[2717], t[2729], t[2728], t[2726], t[2727], t[2678], t[2679], t[2746], t[2680], t[2681], t[2682], t[2683], t[2684], t[2685], t[2686], t[2742], t[2743], t[2741], t[2745], t[2712], t[2714], t[2715], t[2713], t[2694], t[2695], t[2696], t[2697], t[2698], t[2699], t[2747], t[2569], t[2570], t[2571], t[2572], t[2573], t[2574], t[2575], t[2576], t[2577], t[2578], t[2600], t[2579], t[2710], t[2598], x[193]}), .y({t[1350], t[1345], t[1340], t[1335], t[1330], t[1325], t[1320], t[1315], t[1310], t[1305], t[1300], t[1295], t[1290], t[1285], t[1280], t[1275], t[1270], t[1265], t[1260], t[1255], t[1250], t[1245], t[1240], t[1235], t[1230], t[1225], t[1220], t[1215], t[1210], t[1205], t[1200], t[1195], t[1190], t[1185], t[1180], t[1175], t[1170], t[1165], t[1160], t[1155], t[1150], t[1145], t[1140], t[1135], t[1130], t[1125], t[1120], t[1115], t[1110], t[1105], t[1100], t[1095], t[1090], t[1085], t[1080], t[1075], t[1070], t[1065], t[1060], t[1055], t[1050], t[1045], t[1040], t[1035], t[1030], t[1025], t[1020], t[1015], t[1010], t[1005], t[1000], t[995], t[990], t[985], t[980], t[975], t[970], t[965], t[960], t[955], t[950], t[945], t[940], t[935], t[930], t[925], t[920], t[915], t[910], t[905], t[900], t[895], t[890], t[885], t[880], t[875], t[870], t[865], t[860], t[855], t[850], t[845], t[840], t[835], t[830], t[825], t[820], t[815], t[810], t[805], t[800], t[795], t[790], t[785], t[780], t[775], t[770], t[765], t[760], t[755], t[750], t[745], t[740], t[735], t[730], t[725], t[720], t[715], t[710], t[705], t[700], t[695], t[690], t[685], t[680], t[675], t[670], t[665], t[660], t[655], t[650], t[645], t[640], t[635], t[630], t[625], t[620], t[615], t[610], t[605], t[600], t[595], t[590], t[585], t[580], t[575], t[570], t[565], t[560], t[555], t[550], t[545], t[540], t[535], t[530], t[525], t[520], t[515], t[510], t[505], t[500], t[495], t[490], t[485], t[480], t[475], t[470], t[465], t[460], t[455], t[450], t[445], t[440], t[435], t[430], t[425], t[420], t[415], t[410], t[405], t[400], t[395], t[390], t[385], t[380], t[375], t[370], t[365], t[360], t[355], t[350], t[345], t[340], t[335], t[330], t[325], t[320], t[315], t[310], t[305], t[300], t[295], t[290], t[285], t[280], t[275], t[270], t[265], t[260], t[255], t[250], t[245], t[240], t[235], t[230], t[225], t[220], t[215], t[210], t[205], t[200], t[195], t[190], t[185], t[180], t[175], t[170], t[165], t[160], t[155], t[150], t[145], t[140], t[135], t[130], t[125], t[120], t[115], t[110], t[105], t[100], t[95], t[90], t[85], t[80], t[75], t[70], t[65], t[60], t[55], t[50], t[45], t[40], t[35], t[30], t[25], t[20], t[15], t[10], t[5], t[0]}));
  Reg2 Reg2_inst(.x({t[2782], t[2781], t[2780], t[2779], t[3646], t[3645], t[3644], t[3643], t[3642], t[3641], t[3640], t[3639], t[3638], t[3637], t[3636], t[3635], t[3634], t[3633], t[3632], t[3631], t[3862], t[3861], t[3860], t[3859], t[3858], t[3857], t[3856], t[3855], t[3854], t[3853], t[3852], t[3851], t[3850], t[3849], t[3848], t[3847], t[3630], t[3629], t[3628], t[3627], t[3846], t[3845], t[3844], t[3843], t[3842], t[3841], t[3840], t[3839], t[3838], t[3837], t[3836], t[3835], t[3834], t[3833], t[3832], t[3831], t[3830], t[3829], t[3828], t[3827], t[3826], t[3825], t[3824], t[3823], t[3822], t[3821], t[3820], t[3819], t[3818], t[3817], t[3816], t[3815], t[3814], t[3813], t[3812], t[3811], t[3810], t[3809], t[3808], t[3807], t[3626], t[3625], t[3624], t[3623], t[3806], t[3805], t[3804], t[3803], t[3802], t[3801], t[3800], t[3799], t[3798], t[3797], t[3796], t[3795], t[3794], t[3793], t[3792], t[3791], t[3790], t[3789], t[3788], t[3787], t[3786], t[3785], t[3784], t[3783], t[3782], t[3781], t[3780], t[3779], t[3778], t[3777], t[3776], t[3775], t[3774], t[3773], t[3772], t[3771], t[3770], t[3769], t[3768], t[3767], t[3622], t[3621], t[3620], t[3619], t[3766], t[3765], t[3764], t[3763], t[3762], t[3761], t[3760], t[3759], t[3758], t[3757], t[3756], t[3755], t[3754], t[3753], t[3752], t[3751], t[3750], t[3749], t[3748], t[3747], t[3746], t[3745], t[3744], t[3743], t[3742], t[3741], t[3740], t[3739], t[3738], t[3737], t[3736], t[3735], t[3734], t[3733], t[3732], t[3731], t[3730], t[3729], t[3728], t[3727], t[3618], t[3617], t[3616], t[3615], t[3726], t[3725], t[3724], t[3723], t[3722], t[3721], t[3720], t[3719], t[3718], t[3717], t[3716], t[3715], t[3714], t[3713], t[3712], t[3711], t[3710], t[3709], t[3708], t[3707], t[3706], t[3705], t[3704], t[3703], t[3702], t[3701], t[3700], t[3699], t[3698], t[3697], t[3696], t[3695], t[3694], t[3693], t[3692], t[3691], t[3690], t[3689], t[3688], t[3687], t[3614], t[3613], t[3612], t[3611], t[3686], t[3685], t[3684], t[3683], t[3682], t[3681], t[3680], t[3679], t[3678], t[3677], t[3676], t[3675], t[3674], t[3673], t[3672], t[3671], t[3670], t[3669], t[3668], t[3667], t[3666], t[3665], t[3664], t[3663], t[3662], t[3661], t[3660], t[3659], t[3658], t[3657], t[3656], t[3655], t[3654], t[3653], t[3652], t[3651], t[3650], t[3649], t[3648], t[3647], t[3610], t[3609], t[3608], t[3607], t[2878], t[2877], t[2876], t[2875], t[2874], t[2873], t[2872], t[2871], t[2870], t[2869], t[2868], t[2867], t[2866], t[2865], t[2864], t[2863], t[3094], t[3093], t[3092], t[3091], t[3090], t[3089], t[3088], t[3087], t[3086], t[3085], t[3084], t[3083], t[3082], t[3081], t[3080], t[3079], t[2862], t[2861], t[2860], t[2859], t[3078], t[3077], t[3076], t[3075], t[3074], t[3073], t[3072], t[3071], t[3070], t[3069], t[3068], t[3067], t[3066], t[3065], t[3064], t[3063], t[3062], t[3061], t[3060], t[3059], t[3058], t[3057], t[3056], t[3055], t[3054], t[3053], t[3052], t[3051], t[3050], t[3049], t[3048], t[3047], t[3046], t[3045], t[3044], t[3043], t[3042], t[3041], t[3040], t[3039], t[2858], t[2857], t[2856], t[2855], t[3038], t[3037], t[3036], t[3035], t[3034], t[3033], t[3032], t[3031], t[3030], t[3029], t[3028], t[3027], t[3026], t[3025], t[3024], t[3023], t[3022], t[3021], t[3020], t[3019], t[3018], t[3017], t[3016], t[3015], t[3014], t[3013], t[3012], t[3011], t[3010], t[3009], t[3008], t[3007], t[3006], t[3005], t[3004], t[3003], t[3002], t[3001], t[3000], t[2999], t[2854], t[2853], t[2852], t[2851], t[2998], t[2997], t[2996], t[2995], t[2994], t[2993], t[2992], t[2991], t[2990], t[2989], t[2988], t[2987], t[2986], t[2985], t[2984], t[2983], t[2982], t[2981], t[2980], t[2979], t[2978], t[2977], t[2976], t[2975], t[2974], t[2973], t[2972], t[2971], t[2970], t[2969], t[2968], t[2967], t[2966], t[2965], t[2964], t[2963], t[2962], t[2961], t[2960], t[2959], t[2850], t[2849], t[2848], t[2847], t[2958], t[2957], t[2956], t[2955], t[2954], t[2953], t[2952], t[2951], t[2950], t[2949], t[2948], t[2947], t[2946], t[2945], t[2944], t[2943], t[2942], t[2941], t[2940], t[2939], t[2938], t[2937], t[2936], t[2935], t[2934], t[2933], t[2932], t[2931], t[2930], t[2929], t[2928], t[2927], t[2926], t[2925], t[2924], t[2923], t[2922], t[2921], t[2920], t[2919], t[2846], t[2845], t[2844], t[2843], t[2918], t[2917], t[2916], t[2915], t[2914], t[2913], t[2912], t[2911], t[2910], t[2909], t[2908], t[2907], t[2906], t[2905], t[2904], t[2903], t[2902], t[2901], t[2900], t[2899], t[2898], t[2897], t[2896], t[2895], t[2894], t[2893], t[2892], t[2891], t[2890], t[2889], t[2888], t[2887], t[2886], t[2885], t[2884], t[2883], t[2882], t[2881], t[2880], t[2879], t[2842], t[2841], t[2840], t[2839], t[3134], t[3133], t[3132], t[3131], t[3130], t[3129], t[3128], t[3127], t[3126], t[3125], t[3124], t[3123], t[3122], t[3121], t[3120], t[3119], t[3350], t[3349], t[3348], t[3347], t[3346], t[3345], t[3344], t[3343], t[3342], t[3341], t[3340], t[3339], t[3338], t[3337], t[3336], t[3335], t[3118], t[3117], t[3116], t[3115], t[3334], t[3333], t[3332], t[3331], t[3330], t[3329], t[3328], t[3327], t[3326], t[3325], t[3324], t[3323], t[3322], t[3321], t[3320], t[3319], t[3318], t[3317], t[3316], t[3315], t[3314], t[3313], t[3312], t[3311], t[3310], t[3309], t[3308], t[3307], t[3306], t[3305], t[3304], t[3303], t[3302], t[3301], t[3300], t[3299], t[3298], t[3297], t[3296], t[3295], t[3114], t[3113], t[3112], t[3111], t[3294], t[3293], t[3292], t[3291], t[3290], t[3289], t[3288], t[3287], t[3286], t[3285], t[3284], t[3283], t[3282], t[3281], t[3280], t[3279], t[3278], t[3277], t[3276], t[3275], t[3274], t[3273], t[3272], t[3271], t[3270], t[3269], t[3268], t[3267], t[3266], t[3265], t[3264], t[3263], t[3262], t[3261], t[3260], t[3259], t[3258], t[3257], t[3256], t[3255], t[3110], t[3109], t[3108], t[3107], t[3254], t[3253], t[3252], t[3251], t[3250], t[3249], t[3248], t[3247], t[3246], t[3245], t[3244], t[3243], t[3242], t[3241], t[3240], t[3239], t[3238], t[3237], t[3236], t[3235], t[3234], t[3233], t[3232], t[3231], t[3230], t[3229], t[3228], t[3227], t[3226], t[3225], t[3224], t[3223], t[3222], t[3221], t[3220], t[3219], t[3218], t[3217], t[3216], t[3215], t[3106], t[3105], t[3104], t[3103], t[3214], t[3213], t[3212], t[3211], t[3210], t[3209], t[3208], t[3207], t[3206], t[3205], t[3204], t[3203], t[3202], t[3201], t[3200], t[3199], t[3198], t[3197], t[3196], t[3195], t[3194], t[3193], t[3192], t[3191], t[3190], t[3189], t[3188], t[3187], t[3186], t[3185], t[3184], t[3183], t[3182], t[3181], t[3180], t[3179], t[3178], t[3177], t[3176], t[3175], t[3102], t[3101], t[3100], t[3099], t[3174], t[3173], t[3172], t[3171], t[3170], t[3169], t[3168], t[3167], t[3166], t[3165], t[3164], t[3163], t[3162], t[3161], t[3160], t[3159], t[3158], t[3157], t[3156], t[3155], t[3154], t[3153], t[3152], t[3151], t[3150], t[3149], t[3148], t[3147], t[3146], t[3145], t[3144], t[3143], t[3142], t[3141], t[3140], t[3139], t[3138], t[3137], t[3136], t[3135], t[3098], t[3097], t[3096], t[3095], t[3390], t[3389], t[3388], t[3387], t[3386], t[3385], t[3384], t[3383], t[3382], t[3381], t[3380], t[3379], t[3378], t[3377], t[3376], t[3375], t[3606], t[3605], t[3604], t[3603], t[3602], t[3601], t[3600], t[3599], t[3598], t[3597], t[3596], t[3595], t[3594], t[3593], t[3592], t[3591], t[3374], t[3373], t[3372], t[3371], t[3590], t[3589], t[3588], t[3587], t[3586], t[3585], t[3584], t[3583], t[3582], t[3581], t[3580], t[3579], t[3578], t[3577], t[3576], t[3575], t[3574], t[3573], t[3572], t[3571], t[3570], t[3569], t[3568], t[3567], t[3566], t[3565], t[3564], t[3563], t[3562], t[3561], t[3560], t[3559], t[3558], t[3557], t[3556], t[3555], t[3554], t[3553], t[3552], t[3551], t[3370], t[3369], t[3368], t[3367], t[3550], t[3549], t[3548], t[3547], t[3546], t[3545], t[3544], t[3543], t[3542], t[3541], t[3540], t[3539], t[3538], t[3537], t[3536], t[3535], t[3534], t[3533], t[3532], t[3531], t[3530], t[3529], t[3528], t[3527], t[3526], t[3525], t[3524], t[3523], t[3522], t[3521], t[3520], t[3519], t[3518], t[3517], t[3516], t[3515], t[3514], t[3513], t[3512], t[3511], t[3366], t[3365], t[3364], t[3363], t[3510], t[3509], t[3508], t[3507], t[3506], t[3505], t[3504], t[3503], t[3502], t[3501], t[3500], t[3499], t[3498], t[3497], t[3496], t[3495], t[3494], t[3493], t[3492], t[3491], t[3490], t[3489], t[3488], t[3487], t[3486], t[3485], t[3484], t[3483], t[3482], t[3481], t[3480], t[3479], t[3478], t[3477], t[3476], t[3475], t[3474], t[3473], t[3472], t[3471], t[3362], t[3361], t[3360], t[3359], t[3470], t[3469], t[3468], t[3467], t[3466], t[3465], t[3464], t[3463], t[3462], t[3461], t[3460], t[3459], t[3458], t[3457], t[3456], t[3455], t[3454], t[3453], t[3452], t[3451], t[3450], t[3449], t[3448], t[3447], t[3446], t[3445], t[3444], t[3443], t[3442], t[3441], t[3440], t[3439], t[3438], t[3437], t[3436], t[3435], t[3434], t[3433], t[3432], t[3431], t[3358], t[3357], t[3356], t[3355], t[3430], t[3429], t[3428], t[3427], t[3426], t[3425], t[3424], t[3423], t[3422], t[3421], t[3420], t[3419], t[3418], t[3417], t[3416], t[3415], t[3414], t[3413], t[3412], t[3411], t[3410], t[3409], t[3408], t[3407], t[3406], t[3405], t[3404], t[3403], t[3402], t[3401], t[3400], t[3399], t[3398], t[3397], t[3396], t[3395], t[3394], t[3393], t[3392], t[3391], t[3354], t[3353], t[3352], t[3351], t[2806], t[2805], t[2804], t[2803], t[2802], t[2801], t[2800], t[2799], t[2798], t[2797], t[2796], t[2795], t[2794], t[2793], t[2792], t[2791], t[2790], t[2789], t[2788], t[2787], t[2786], t[2785], t[2784], t[2783], t[2822], t[2821], t[2820], t[2819], t[2818], t[2817], t[2816], t[2815], t[2814], t[2813], t[2812], t[2811], t[2810], t[2809], t[2808], t[2807], t[2834], t[2833], t[2832], t[2831], t[2830], t[2829], t[2828], t[2827], t[2826], t[2825], t[2824], t[2823], t[2838], t[2837], t[2836], t[2835], x[193]}), .y({t[1354], t[1353], t[1352], t[1351], t[1349], t[1348], t[1347], t[1346], t[1344], t[1343], t[1342], t[1341], t[1339], t[1338], t[1337], t[1336], t[1334], t[1333], t[1332], t[1331], t[1329], t[1328], t[1327], t[1326], t[1324], t[1323], t[1322], t[1321], t[1319], t[1318], t[1317], t[1316], t[1314], t[1313], t[1312], t[1311], t[1309], t[1308], t[1307], t[1306], t[1304], t[1303], t[1302], t[1301], t[1299], t[1298], t[1297], t[1296], t[1294], t[1293], t[1292], t[1291], t[1289], t[1288], t[1287], t[1286], t[1284], t[1283], t[1282], t[1281], t[1279], t[1278], t[1277], t[1276], t[1274], t[1273], t[1272], t[1271], t[1269], t[1268], t[1267], t[1266], t[1264], t[1263], t[1262], t[1261], t[1259], t[1258], t[1257], t[1256], t[1254], t[1253], t[1252], t[1251], t[1249], t[1248], t[1247], t[1246], t[1244], t[1243], t[1242], t[1241], t[1239], t[1238], t[1237], t[1236], t[1234], t[1233], t[1232], t[1231], t[1229], t[1228], t[1227], t[1226], t[1224], t[1223], t[1222], t[1221], t[1219], t[1218], t[1217], t[1216], t[1214], t[1213], t[1212], t[1211], t[1209], t[1208], t[1207], t[1206], t[1204], t[1203], t[1202], t[1201], t[1199], t[1198], t[1197], t[1196], t[1194], t[1193], t[1192], t[1191], t[1189], t[1188], t[1187], t[1186], t[1184], t[1183], t[1182], t[1181], t[1179], t[1178], t[1177], t[1176], t[1174], t[1173], t[1172], t[1171], t[1169], t[1168], t[1167], t[1166], t[1164], t[1163], t[1162], t[1161], t[1159], t[1158], t[1157], t[1156], t[1154], t[1153], t[1152], t[1151], t[1149], t[1148], t[1147], t[1146], t[1144], t[1143], t[1142], t[1141], t[1139], t[1138], t[1137], t[1136], t[1134], t[1133], t[1132], t[1131], t[1129], t[1128], t[1127], t[1126], t[1124], t[1123], t[1122], t[1121], t[1119], t[1118], t[1117], t[1116], t[1114], t[1113], t[1112], t[1111], t[1109], t[1108], t[1107], t[1106], t[1104], t[1103], t[1102], t[1101], t[1099], t[1098], t[1097], t[1096], t[1094], t[1093], t[1092], t[1091], t[1089], t[1088], t[1087], t[1086], t[1084], t[1083], t[1082], t[1081], t[1079], t[1078], t[1077], t[1076], t[1074], t[1073], t[1072], t[1071], t[1069], t[1068], t[1067], t[1066], t[1064], t[1063], t[1062], t[1061], t[1059], t[1058], t[1057], t[1056], t[1054], t[1053], t[1052], t[1051], t[1049], t[1048], t[1047], t[1046], t[1044], t[1043], t[1042], t[1041], t[1039], t[1038], t[1037], t[1036], t[1034], t[1033], t[1032], t[1031], t[1029], t[1028], t[1027], t[1026], t[1024], t[1023], t[1022], t[1021], t[1019], t[1018], t[1017], t[1016], t[1014], t[1013], t[1012], t[1011], t[1009], t[1008], t[1007], t[1006], t[1004], t[1003], t[1002], t[1001], t[999], t[998], t[997], t[996], t[994], t[993], t[992], t[991], t[989], t[988], t[987], t[986], t[984], t[983], t[982], t[981], t[979], t[978], t[977], t[976], t[974], t[973], t[972], t[971], t[969], t[968], t[967], t[966], t[964], t[963], t[962], t[961], t[959], t[958], t[957], t[956], t[954], t[953], t[952], t[951], t[949], t[948], t[947], t[946], t[944], t[943], t[942], t[941], t[939], t[938], t[937], t[936], t[934], t[933], t[932], t[931], t[929], t[928], t[927], t[926], t[924], t[923], t[922], t[921], t[919], t[918], t[917], t[916], t[914], t[913], t[912], t[911], t[909], t[908], t[907], t[906], t[904], t[903], t[902], t[901], t[899], t[898], t[897], t[896], t[894], t[893], t[892], t[891], t[889], t[888], t[887], t[886], t[884], t[883], t[882], t[881], t[879], t[878], t[877], t[876], t[874], t[873], t[872], t[871], t[869], t[868], t[867], t[866], t[864], t[863], t[862], t[861], t[859], t[858], t[857], t[856], t[854], t[853], t[852], t[851], t[849], t[848], t[847], t[846], t[844], t[843], t[842], t[841], t[839], t[838], t[837], t[836], t[834], t[833], t[832], t[831], t[829], t[828], t[827], t[826], t[824], t[823], t[822], t[821], t[819], t[818], t[817], t[816], t[814], t[813], t[812], t[811], t[809], t[808], t[807], t[806], t[804], t[803], t[802], t[801], t[799], t[798], t[797], t[796], t[794], t[793], t[792], t[791], t[789], t[788], t[787], t[786], t[784], t[783], t[782], t[781], t[779], t[778], t[777], t[776], t[774], t[773], t[772], t[771], t[769], t[768], t[767], t[766], t[764], t[763], t[762], t[761], t[759], t[758], t[757], t[756], t[754], t[753], t[752], t[751], t[749], t[748], t[747], t[746], t[744], t[743], t[742], t[741], t[739], t[738], t[737], t[736], t[734], t[733], t[732], t[731], t[729], t[728], t[727], t[726], t[724], t[723], t[722], t[721], t[719], t[718], t[717], t[716], t[714], t[713], t[712], t[711], t[709], t[708], t[707], t[706], t[704], t[703], t[702], t[701], t[699], t[698], t[697], t[696], t[694], t[693], t[692], t[691], t[689], t[688], t[687], t[686], t[684], t[683], t[682], t[681], t[679], t[678], t[677], t[676], t[674], t[673], t[672], t[671], t[669], t[668], t[667], t[666], t[664], t[663], t[662], t[661], t[659], t[658], t[657], t[656], t[654], t[653], t[652], t[651], t[649], t[648], t[647], t[646], t[644], t[643], t[642], t[641], t[639], t[638], t[637], t[636], t[634], t[633], t[632], t[631], t[629], t[628], t[627], t[626], t[624], t[623], t[622], t[621], t[619], t[618], t[617], t[616], t[614], t[613], t[612], t[611], t[609], t[608], t[607], t[606], t[604], t[603], t[602], t[601], t[599], t[598], t[597], t[596], t[594], t[593], t[592], t[591], t[589], t[588], t[587], t[586], t[584], t[583], t[582], t[581], t[579], t[578], t[577], t[576], t[574], t[573], t[572], t[571], t[569], t[568], t[567], t[566], t[564], t[563], t[562], t[561], t[559], t[558], t[557], t[556], t[554], t[553], t[552], t[551], t[549], t[548], t[547], t[546], t[544], t[543], t[542], t[541], t[539], t[538], t[537], t[536], t[534], t[533], t[532], t[531], t[529], t[528], t[527], t[526], t[524], t[523], t[522], t[521], t[519], t[518], t[517], t[516], t[514], t[513], t[512], t[511], t[509], t[508], t[507], t[506], t[504], t[503], t[502], t[501], t[499], t[498], t[497], t[496], t[494], t[493], t[492], t[491], t[489], t[488], t[487], t[486], t[484], t[483], t[482], t[481], t[479], t[478], t[477], t[476], t[474], t[473], t[472], t[471], t[469], t[468], t[467], t[466], t[464], t[463], t[462], t[461], t[459], t[458], t[457], t[456], t[454], t[453], t[452], t[451], t[449], t[448], t[447], t[446], t[444], t[443], t[442], t[441], t[439], t[438], t[437], t[436], t[434], t[433], t[432], t[431], t[429], t[428], t[427], t[426], t[424], t[423], t[422], t[421], t[419], t[418], t[417], t[416], t[414], t[413], t[412], t[411], t[409], t[408], t[407], t[406], t[404], t[403], t[402], t[401], t[399], t[398], t[397], t[396], t[394], t[393], t[392], t[391], t[389], t[388], t[387], t[386], t[384], t[383], t[382], t[381], t[379], t[378], t[377], t[376], t[374], t[373], t[372], t[371], t[369], t[368], t[367], t[366], t[364], t[363], t[362], t[361], t[359], t[358], t[357], t[356], t[354], t[353], t[352], t[351], t[349], t[348], t[347], t[346], t[344], t[343], t[342], t[341], t[339], t[338], t[337], t[336], t[334], t[333], t[332], t[331], t[329], t[328], t[327], t[326], t[324], t[323], t[322], t[321], t[319], t[318], t[317], t[316], t[314], t[313], t[312], t[311], t[309], t[308], t[307], t[306], t[304], t[303], t[302], t[301], t[299], t[298], t[297], t[296], t[294], t[293], t[292], t[291], t[289], t[288], t[287], t[286], t[284], t[283], t[282], t[281], t[279], t[278], t[277], t[276], t[274], t[273], t[272], t[271], t[269], t[268], t[267], t[266], t[264], t[263], t[262], t[261], t[259], t[258], t[257], t[256], t[254], t[253], t[252], t[251], t[249], t[248], t[247], t[246], t[244], t[243], t[242], t[241], t[239], t[238], t[237], t[236], t[234], t[233], t[232], t[231], t[229], t[228], t[227], t[226], t[224], t[223], t[222], t[221], t[219], t[218], t[217], t[216], t[214], t[213], t[212], t[211], t[209], t[208], t[207], t[206], t[204], t[203], t[202], t[201], t[199], t[198], t[197], t[196], t[194], t[193], t[192], t[191], t[189], t[188], t[187], t[186], t[184], t[183], t[182], t[181], t[179], t[178], t[177], t[176], t[174], t[173], t[172], t[171], t[169], t[168], t[167], t[166], t[164], t[163], t[162], t[161], t[159], t[158], t[157], t[156], t[154], t[153], t[152], t[151], t[149], t[148], t[147], t[146], t[144], t[143], t[142], t[141], t[139], t[138], t[137], t[136], t[134], t[133], t[132], t[131], t[129], t[128], t[127], t[126], t[124], t[123], t[122], t[121], t[119], t[118], t[117], t[116], t[114], t[113], t[112], t[111], t[109], t[108], t[107], t[106], t[104], t[103], t[102], t[101], t[99], t[98], t[97], t[96], t[94], t[93], t[92], t[91], t[89], t[88], t[87], t[86], t[84], t[83], t[82], t[81], t[79], t[78], t[77], t[76], t[74], t[73], t[72], t[71], t[69], t[68], t[67], t[66], t[64], t[63], t[62], t[61], t[59], t[58], t[57], t[56], t[54], t[53], t[52], t[51], t[49], t[48], t[47], t[46], t[44], t[43], t[42], t[41], t[39], t[38], t[37], t[36], t[34], t[33], t[32], t[31], t[29], t[28], t[27], t[26], t[24], t[23], t[22], t[21], t[19], t[18], t[17], t[16], t[14], t[13], t[12], t[11], t[9], t[8], t[7], t[6], t[4], t[3], t[2], t[1]}));
  multiplexer #(.WIDTH(65)) multiplexer_inst(.s({t[2775], t[2776], t[2777], t[2778], t[2439]}), .d({t[2503], t[2502], t[2501], t[2500], t[2499], t[2498], t[2497], t[2496], t[2495], t[2494], t[2493], t[2492], t[2491], t[2490], t[2489], t[2488], t[2487], t[2486], t[2485], t[2484], t[2483], t[2482], t[2481], t[2480], t[2479], t[2478], t[2477], t[2476], t[2475], t[2474], t[2473], t[2472], t[2471], t[2470], t[2469], t[2468], t[2467], t[2466], t[2465], t[2464], t[2463], t[2462], t[2461], t[2460], t[2459], t[2458], t[2457], t[2456], t[2455], t[2454], t[2453], t[2452], t[2451], t[2450], t[2449], t[2448], t[2447], t[2446], t[2445], t[2444], t[2443], t[2442], t[2441], t[2440], t[2775]}), .q({y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], y[8], y[9], y[10], y[11], y[12], y[13], y[14], y[15], y[16], y[17], y[18], y[19], y[20], y[21], y[22], y[23], y[24], y[25], y[26], y[27], y[28], y[29], y[30], y[31], y[32], y[33], y[34], y[35], y[36], y[37], y[38], y[39], y[40], y[41], y[42], y[43], y[44], y[45], y[46], y[47], y[48], y[49], y[50], y[51], y[52], y[53], y[54], y[55], y[56], y[57], y[58], y[59], y[60], y[61], y[62], y[63], y[64]}));
endmodule

module register_stage(clk, D, Q);
  parameter WIDTH = 8;
  input clk;
  input [WIDTH-1:0] D;
  output [WIDTH-1:0] Q;

  reg [WIDTH-1:0] s_current_state;
  wire [WIDTH-1:0] s_next_state;
  assign s_next_state = D;
  always @ (posedge clk)
  begin
      s_current_state <= s_next_state;
  end
  assign Q = s_current_state;
endmodule

module multiplexer(s, d, q);
  parameter WIDTH = 8;
  input [4:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  muxtree #(.WIDTH(65)) inst_0(.s(s), .d({d[0],d[1],d[2],d[3],d[4],d[5],d[6],d[7],d[8],d[9],d[10],d[11],d[12],d[13],d[14],d[15],d[16],d[17],d[18],d[19],d[20],d[21],d[22],d[23],d[24],d[25],d[26],d[27],d[28],d[29],d[30],d[31],d[32],d[33],d[34],d[35],d[36],d[37],d[38],d[39],d[40],d[41],d[42],d[43],d[44],d[45],d[46],d[47],d[48],d[49],d[50],d[51],d[52],d[53],d[54],d[55],d[56],d[57],d[58],d[59],d[60],d[61],d[62],d[63],d[64]}), .q({q[0],q[1],q[2],q[3],q[4],q[5],q[6],q[7],q[8],q[9],q[10],q[11],q[12],q[13],q[14],q[15],q[16],q[17],q[18],q[19],q[20],q[21],q[22],q[23],q[24],q[25],q[26],q[27],q[28],q[29],q[30],q[31],q[32],q[33],q[34],q[35],q[36],q[37],q[38],q[39],q[40],q[41],q[42],q[43],q[44],q[45],q[46],q[47],q[48],q[49],q[50],q[51],q[52],q[53],q[54],q[55],q[56],q[57],q[58],q[59],q[60],q[61],q[62],q[63],q[64]}));
endmodule

module muxtree(s, d, q);
  parameter WIDTH = 8;
  input [4:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  wire [WIDTH-1:0] v0_0;
  wire [WIDTH-1:0] v0_1;
  wire [WIDTH-1:0] v1_0;
  wire [WIDTH-1:0] v1_1;
  wire [WIDTH-1:0] v1_2;
  wire [WIDTH-1:0] v1_3;
  wire [WIDTH-1:0] v2_0;
  wire [WIDTH-1:0] v2_1;
  wire [WIDTH-1:0] v2_2;
  wire [WIDTH-1:0] v2_3;
  wire [WIDTH-1:0] v2_4;
  wire [WIDTH-1:0] v2_5;
  wire [WIDTH-1:0] v2_6;
  wire [WIDTH-1:0] v2_7;
  wire [WIDTH-1:0] v3_0;
  wire [WIDTH-1:0] v3_1;
  wire [WIDTH-1:0] v3_2;
  wire [WIDTH-1:0] v3_3;
  wire [WIDTH-1:0] v3_4;
  wire [WIDTH-1:0] v3_5;
  wire [WIDTH-1:0] v3_6;
  wire [WIDTH-1:0] v3_7;
  wire [WIDTH-1:0] v3_8;
  wire [WIDTH-1:0] v3_9;
  wire [WIDTH-1:0] v3_10;
  wire [WIDTH-1:0] v3_11;
  wire [WIDTH-1:0] v3_12;
  wire [WIDTH-1:0] v3_13;
  wire [WIDTH-1:0] v3_14;
  wire [WIDTH-1:0] v3_15;

  assign q = s[0] ? v0_1 : {WIDTH{1'b0}};

  assign v0_0 = s[1] ? v1_1 : {WIDTH{1'b0}};
  assign v0_1 = s[1] ? v1_3 : {WIDTH{1'b0}};

  assign v1_0 = s[2] ? v2_1 : {WIDTH{1'b0}};
  assign v1_1 = s[2] ? v2_3 : {WIDTH{1'b0}};
  assign v1_2 = s[2] ? v2_5 : {WIDTH{1'b0}};
  assign v1_3 = s[2] ? v2_7 : {WIDTH{1'b0}};

  assign v2_0 = s[3] ? v3_1 : {WIDTH{1'b0}};
  assign v2_1 = s[3] ? v3_3 : {WIDTH{1'b0}};
  assign v2_2 = s[3] ? v3_5 : {WIDTH{1'b0}};
  assign v2_3 = s[3] ? v3_7 : {WIDTH{1'b0}};
  assign v2_4 = s[3] ? v3_9 : {WIDTH{1'b0}};
  assign v2_5 = s[3] ? v3_11 : {WIDTH{1'b0}};
  assign v2_6 = s[3] ? v3_13 : {WIDTH{1'b0}};
  assign v2_7 = s[3] ? v3_15 : {WIDTH{1'b0}};

  assign v3_0 = {WIDTH{1'b0}};
  assign v3_1 = {WIDTH{1'b0}};
  assign v3_2 = {WIDTH{1'b0}};
  assign v3_3 = {WIDTH{1'b0}};
  assign v3_4 = {WIDTH{1'b0}};
  assign v3_5 = {WIDTH{1'b0}};
  assign v3_6 = {WIDTH{1'b0}};
  assign v3_7 = {WIDTH{1'b0}};
  assign v3_8 = {WIDTH{1'b0}};
  assign v3_9 = {WIDTH{1'b0}};
  assign v3_10 = {WIDTH{1'b0}};
  assign v3_11 = {WIDTH{1'b0}};
  assign v3_12 = {WIDTH{1'b0}};
  assign v3_13 = {WIDTH{1'b0}};
  assign v3_14 = {WIDTH{1'b0}};
  assign v3_15 = s[4] ? d : {WIDTH{1'b0}};

endmodule

