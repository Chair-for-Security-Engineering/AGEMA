/* modified netlist. Source: module CRAFT in file ../CaseStudies/09_CRAFT_round_based_encryption/FPGA_based/CRAFT_synthesis.v */
/* clock gating is added to the circuit, the latency increased 1 time(s)  */

module CRAFT_GHPCLL_ClockGating_d1 (clk, rst, Input_s0, Key_s0, Key_s1, Input_s1, Fresh, done, Output_s0, Output_s1, Synch);
    input clk ;
    input rst ;
    input [63:0] Input_s0 ;
    input [127:0] Key_s0 ;
    input [127:0] Key_s1 ;
    input [63:0] Input_s1 ;
    input [1023:0] Fresh ;
    output done ;
    output [63:0] Output_s0 ;
    output [63:0] Output_s1 ;
    output Synch ;
    wire [6:1] \FSM ;
    wire [6:2] \FSMUpdate ;
    wire done_internal ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N10 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N30 ;
    wire N32 ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N50 ;
    wire N52 ;
    wire N54 ;
    wire N55 ;
    wire N57 ;
    wire N58 ;
    wire N60 ;
    wire N61 ;
    wire N63 ;
    wire N64 ;
    wire N66 ;
    wire N67 ;
    wire N69 ;
    wire N70 ;
    wire N72 ;
    wire N73 ;
    wire N75 ;
    wire N77 ;
    wire N79 ;
    wire N81 ;
    wire N83 ;
    wire N85 ;
    wire N87 ;
    wire N89 ;
    wire N91 ;
    wire N93 ;
    wire N95 ;
    wire N97 ;
    wire N99 ;
    wire N101 ;
    wire N103 ;
    wire N105 ;
    wire N107 ;
    wire [6:0] \FSMRegInst/s_current_state ;
    wire [0:0] \selectsRegInst/s_current_state ;
    wire [0:0] selectsNext ;
    wire [63:0] Feedback ;
    wire [63:0] AddRoundKeyOutput ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_739 ;
    wire new_AGEMA_signal_740 ;
    wire new_AGEMA_signal_741 ;
    wire new_AGEMA_signal_742 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_749 ;
    wire new_AGEMA_signal_750 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_782 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[1].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [1]), .O (\FSM [1]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[2].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [2]), .O (\FSM [2]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[4].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [4]), .O (\FSM [4]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[5].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [5]), .O (\FSM [5]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[6].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [6]), .O (\FSM [6]) ) ;
    LUT3 #( .INIT ( 8'h54 ) ) \FSMSignalsInst/done<6>_SW0 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [5]), .I2 (\FSMRegInst/s_current_state [4]), .O (N2) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[0].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[32], Key_s0[32]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[96], Key_s0[96]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_857, N4}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[1].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[33], Key_s0[33]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[97], Key_s0[97]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_860, N6}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[2].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[34], Key_s0[34]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[98], Key_s0[98]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_863, N8}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[3].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[35], Key_s0[35]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[99], Key_s0[99]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_866, N10}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[4].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[36], Key_s0[36]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[100], Key_s0[100]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_869, N12}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[5].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[37], Key_s0[37]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[101], Key_s0[101]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_872, N14}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[6].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[38], Key_s0[38]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[102], Key_s0[102]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_875, N16}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[7].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[39], Key_s0[39]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[103], Key_s0[103]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_878, N18}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[11].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[43], Key_s0[43]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[107], Key_s0[107]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_881, N20}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[0].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[48], Key_s0[48]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[112], Key_s0[112]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_884, N22}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[1].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[49], Key_s0[49]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[113], Key_s0[113]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_887, N24}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[2].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[50], Key_s0[50]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[114], Key_s0[114]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_890, N26}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[3].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[51], Key_s0[51]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[115], Key_s0[115]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_893, N28}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[4].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[52], Key_s0[52]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[116], Key_s0[116]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_896, N30}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[5].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[53], Key_s0[53]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[117], Key_s0[117]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_899, N32}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[6].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[54], Key_s0[54]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[118], Key_s0[118]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_902, N34}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[7].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[55], Key_s0[55]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[119], Key_s0[119]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_905, N36}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[8].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[56], Key_s0[56]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[120], Key_s0[120]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_908, N38}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[9].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[57], Key_s0[57]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[121], Key_s0[121]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_911, N40}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[10].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[58], Key_s0[58]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[122], Key_s0[122]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_914, N42}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[11].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[59], Key_s0[59]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[123], Key_s0[123]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_917, N44}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[12].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[60], Key_s0[60]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[124], Key_s0[124]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_920, N46}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[13].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[61], Key_s0[61]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[125], Key_s0[125]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_923, N48}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[14].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[62], Key_s0[62]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[126], Key_s0[126]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_926, N50}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[15].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[63], Key_s0[63]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[127], Key_s0[127]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_929, N52}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[46], Key_s0[46]}), .I1 ({Key_s1[110], Key_s0[110]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_932, N54}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[110], Key_s0[110]}), .I1 ({Input_s1[46], Input_s0[46]}), .I2 ({Input_s1[14], Input_s0[14]}), .O ({new_AGEMA_signal_935, N55}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[45], Key_s0[45]}), .I1 ({Key_s1[109], Key_s0[109]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_938, N57}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[109], Key_s0[109]}), .I1 ({Input_s1[45], Input_s0[45]}), .I2 ({Input_s1[13], Input_s0[13]}), .O ({new_AGEMA_signal_941, N58}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[47], Key_s0[47]}), .I1 ({Key_s1[111], Key_s0[111]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_944, N60}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[111], Key_s0[111]}), .I1 ({Input_s1[47], Input_s0[47]}), .I2 ({Input_s1[15], Input_s0[15]}), .O ({new_AGEMA_signal_947, N61}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[44], Key_s0[44]}), .I1 ({Key_s1[108], Key_s0[108]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_950, N63}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[108], Key_s0[108]}), .I1 ({Input_s1[44], Input_s0[44]}), .I2 ({Input_s1[12], Input_s0[12]}), .O ({new_AGEMA_signal_953, N64}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[42], Key_s0[42]}), .I1 ({Key_s1[106], Key_s0[106]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_956, N66}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[106], Key_s0[106]}), .I1 ({Input_s1[42], Input_s0[42]}), .I2 ({Input_s1[10], Input_s0[10]}), .O ({new_AGEMA_signal_959, N67}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[41], Key_s0[41]}), .I1 ({Key_s1[105], Key_s0[105]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_962, N69}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[105], Key_s0[105]}), .I1 ({Input_s1[9], Input_s0[9]}), .I2 ({Input_s1[41], Input_s0[41]}), .O ({new_AGEMA_signal_965, N70}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[40], Key_s0[40]}), .I1 ({Key_s1[104], Key_s0[104]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_968, N72}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[104], Key_s0[104]}), .I1 ({Input_s1[8], Input_s0[8]}), .I2 ({Input_s1[40], Input_s0[40]}), .O ({new_AGEMA_signal_971, N73}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[48], Input_s0[48]}), .I1 ({Input_s1[16], Input_s0[16]}), .I2 ({Input_s1[0], Input_s0[0]}), .O ({new_AGEMA_signal_975, N75}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[49], Input_s0[49]}), .I1 ({Input_s1[1], Input_s0[1]}), .I2 ({Input_s1[17], Input_s0[17]}), .O ({new_AGEMA_signal_979, N77}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[50], Input_s0[50]}), .I1 ({Input_s1[2], Input_s0[2]}), .I2 ({Input_s1[18], Input_s0[18]}), .O ({new_AGEMA_signal_983, N79}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[51], Input_s0[51]}), .I1 ({Input_s1[3], Input_s0[3]}), .I2 ({Input_s1[19], Input_s0[19]}), .O ({new_AGEMA_signal_987, N81}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[52], Input_s0[52]}), .I1 ({Input_s1[4], Input_s0[4]}), .I2 ({Input_s1[20], Input_s0[20]}), .O ({new_AGEMA_signal_991, N83}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[5], Input_s0[5]}), .I1 ({Input_s1[53], Input_s0[53]}), .I2 ({Input_s1[21], Input_s0[21]}), .O ({new_AGEMA_signal_995, N85}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[6], Input_s0[6]}), .I1 ({Input_s1[54], Input_s0[54]}), .I2 ({Input_s1[22], Input_s0[22]}), .O ({new_AGEMA_signal_999, N87}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[7], Input_s0[7]}), .I1 ({Input_s1[55], Input_s0[55]}), .I2 ({Input_s1[23], Input_s0[23]}), .O ({new_AGEMA_signal_1003, N89}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[8], Input_s0[8]}), .I1 ({Input_s1[56], Input_s0[56]}), .I2 ({Input_s1[24], Input_s0[24]}), .O ({new_AGEMA_signal_1006, N91}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[9], Input_s0[9]}), .I1 ({Input_s1[57], Input_s0[57]}), .I2 ({Input_s1[25], Input_s0[25]}), .O ({new_AGEMA_signal_1009, N93}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[58], Input_s0[58]}), .I1 ({Input_s1[26], Input_s0[26]}), .I2 ({Input_s1[10], Input_s0[10]}), .O ({new_AGEMA_signal_1012, N95}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[59], Input_s0[59]}), .I1 ({Input_s1[27], Input_s0[27]}), .I2 ({Input_s1[11], Input_s0[11]}), .O ({new_AGEMA_signal_1016, N97}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[60], Input_s0[60]}), .I1 ({Input_s1[28], Input_s0[28]}), .I2 ({Input_s1[12], Input_s0[12]}), .O ({new_AGEMA_signal_1019, N99}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[61], Input_s0[61]}), .I1 ({Input_s1[29], Input_s0[29]}), .I2 ({Input_s1[13], Input_s0[13]}), .O ({new_AGEMA_signal_1022, N101}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[62], Input_s0[62]}), .I1 ({Input_s1[30], Input_s0[30]}), .I2 ({Input_s1[14], Input_s0[14]}), .O ({new_AGEMA_signal_1025, N103}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[63], Input_s0[63]}), .I1 ({Input_s1[31], Input_s0[31]}), .I2 ({Input_s1[15], Input_s0[15]}), .O ({new_AGEMA_signal_1028, N105}) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \selectsUpdateInst/selectsNext<0>1 ( .I0 (\selectsRegInst/s_current_state [0]), .I1 (rst), .O (selectsNext[0]) ) ;
    LUT3 #( .INIT ( 8'hBE ) ) \FSMUpdateInst/Mxor_FSMUpdate<2>_xo<0>1 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [1]), .I2 (\FSMRegInst/s_current_state [0]), .O (\FSMUpdate [2]) ) ;
    LUT3 #( .INIT ( 8'hBE ) ) \FSMUpdateInst/Mxor_FSMUpdate<6>_xo<0>1 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [4]), .I2 (\FSMRegInst/s_current_state [3]), .O (\FSMUpdate [6]) ) ;
    MUXF7 \FSMSignalsInst/done<6> ( .S (N2), .I0 (N107), .I1 (1'b0), .O (done_internal) ) ;
    LUT6 #( .INIT ( 64'h0000000000000080 ) ) \FSMSignalsInst/done<6>_F ( .I0 (\FSMRegInst/s_current_state [0]), .I1 (\FSMRegInst/s_current_state [6]), .I2 (\FSMRegInst/s_current_state [2]), .I3 (rst), .I4 (\FSMRegInst/s_current_state [1]), .I5 (\FSMRegInst/s_current_state [3]), .O (N107) ) ;
    ClockGatingController #(2) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[0].SboxInst/y_0 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .O ({new_AGEMA_signal_731, Feedback[0]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[0].SboxInst/y_1 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .O ({new_AGEMA_signal_732, Feedback[1]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[0].SboxInst/y_2 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .O ({new_AGEMA_signal_733, Feedback[2]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[0].SboxInst/y_3 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .O ({new_AGEMA_signal_734, Feedback[3]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[1].SboxInst/y_0 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .O ({new_AGEMA_signal_739, Feedback[4]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[1].SboxInst/y_1 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .O ({new_AGEMA_signal_740, Feedback[5]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[1].SboxInst/y_2 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .O ({new_AGEMA_signal_741, Feedback[6]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[1].SboxInst/y_3 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .O ({new_AGEMA_signal_742, Feedback[7]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[2].SboxInst/y_0 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .O ({new_AGEMA_signal_747, Feedback[8]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[2].SboxInst/y_1 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .O ({new_AGEMA_signal_748, Feedback[9]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[2].SboxInst/y_2 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r ({Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .O ({new_AGEMA_signal_749, Feedback[10]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[2].SboxInst/y_3 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176]}), .O ({new_AGEMA_signal_750, Feedback[11]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[3].SboxInst/y_0 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r ({Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .O ({new_AGEMA_signal_755, Feedback[12]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[3].SboxInst/y_1 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r ({Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208]}), .O ({new_AGEMA_signal_756, Feedback[13]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[3].SboxInst/y_2 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224]}), .O ({new_AGEMA_signal_757, Feedback[14]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[3].SboxInst/y_3 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .O ({new_AGEMA_signal_758, Feedback[15]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[4].SboxInst/y_0 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r ({Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .O ({new_AGEMA_signal_763, Feedback[16]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[4].SboxInst/y_1 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272]}), .O ({new_AGEMA_signal_764, Feedback[17]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[4].SboxInst/y_2 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r ({Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .O ({new_AGEMA_signal_765, Feedback[18]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[4].SboxInst/y_3 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304]}), .O ({new_AGEMA_signal_766, Feedback[19]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[5].SboxInst/y_0 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .O ({new_AGEMA_signal_771, Feedback[20]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[5].SboxInst/y_1 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r ({Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .O ({new_AGEMA_signal_772, Feedback[21]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[5].SboxInst/y_2 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r ({Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352]}), .O ({new_AGEMA_signal_773, Feedback[22]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[5].SboxInst/y_3 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368]}), .O ({new_AGEMA_signal_774, Feedback[23]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[6].SboxInst/y_0 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .O ({new_AGEMA_signal_779, Feedback[24]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[6].SboxInst/y_1 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r ({Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .O ({new_AGEMA_signal_780, Feedback[25]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[6].SboxInst/y_2 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416]}), .O ({new_AGEMA_signal_781, Feedback[26]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[6].SboxInst/y_3 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .O ({new_AGEMA_signal_782, Feedback[27]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[7].SboxInst/y_0 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r ({Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .O ({new_AGEMA_signal_787, Feedback[28]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[7].SboxInst/y_1 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464]}), .O ({new_AGEMA_signal_788, Feedback[29]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[7].SboxInst/y_2 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r ({Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .O ({new_AGEMA_signal_789, Feedback[30]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[7].SboxInst/y_3 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496]}), .O ({new_AGEMA_signal_790, Feedback[31]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[8].SboxInst/y_0 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .O ({new_AGEMA_signal_795, Feedback[32]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[8].SboxInst/y_1 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r ({Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .O ({new_AGEMA_signal_796, Feedback[33]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[8].SboxInst/y_2 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544]}), .O ({new_AGEMA_signal_797, Feedback[34]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[8].SboxInst/y_3 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .O ({new_AGEMA_signal_798, Feedback[35]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[9].SboxInst/y_0 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r ({Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .O ({new_AGEMA_signal_803, Feedback[36]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[9].SboxInst/y_1 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r ({Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592]}), .O ({new_AGEMA_signal_804, Feedback[37]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[9].SboxInst/y_2 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608]}), .O ({new_AGEMA_signal_805, Feedback[38]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[9].SboxInst/y_3 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .O ({new_AGEMA_signal_806, Feedback[39]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[10].SboxInst/y_0 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r ({Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .O ({new_AGEMA_signal_811, Feedback[40]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[10].SboxInst/y_1 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656]}), .O ({new_AGEMA_signal_812, Feedback[41]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[10].SboxInst/y_2 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r ({Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .O ({new_AGEMA_signal_813, Feedback[42]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[10].SboxInst/y_3 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688]}), .O ({new_AGEMA_signal_814, Feedback[43]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[11].SboxInst/y_0 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .O ({new_AGEMA_signal_819, Feedback[44]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[11].SboxInst/y_1 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r ({Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .O ({new_AGEMA_signal_820, Feedback[45]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[11].SboxInst/y_2 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r ({Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736]}), .O ({new_AGEMA_signal_821, Feedback[46]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[11].SboxInst/y_3 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752]}), .O ({new_AGEMA_signal_822, Feedback[47]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[12].SboxInst/y_0 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r ({Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .O ({new_AGEMA_signal_827, Feedback[48]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[12].SboxInst/y_1 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784]}), .O ({new_AGEMA_signal_828, Feedback[49]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[12].SboxInst/y_2 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .O ({new_AGEMA_signal_829, Feedback[50]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[12].SboxInst/y_3 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .O ({new_AGEMA_signal_830, Feedback[51]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[13].SboxInst/y_0 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r ({Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .O ({new_AGEMA_signal_835, Feedback[52]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[13].SboxInst/y_1 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848]}), .O ({new_AGEMA_signal_836, Feedback[53]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[13].SboxInst/y_2 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .O ({new_AGEMA_signal_837, Feedback[54]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[13].SboxInst/y_3 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .O ({new_AGEMA_signal_838, Feedback[55]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[14].SboxInst/y_0 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .O ({new_AGEMA_signal_843, Feedback[56]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[14].SboxInst/y_1 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r ({Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .O ({new_AGEMA_signal_844, Feedback[57]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[14].SboxInst/y_2 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r ({Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928]}), .O ({new_AGEMA_signal_845, Feedback[58]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[14].SboxInst/y_3 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944]}), .O ({new_AGEMA_signal_846, Feedback[59]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[15].SboxInst/y_0 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r ({Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .O ({new_AGEMA_signal_851, Feedback[60]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[15].SboxInst/y_1 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r ({Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976]}), .O ({new_AGEMA_signal_852, Feedback[61]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[15].SboxInst/y_2 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992]}), .O ({new_AGEMA_signal_853, Feedback[62]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[15].SboxInst/y_3 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .O ({new_AGEMA_signal_854, Feedback[63]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[0], Input_s0[0]}), .I1 ({Key_s1[0], Key_s0[0]}), .I2 ({Key_s1[64], Key_s0[64]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1031, AddRoundKeyOutput[0]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[10], Input_s0[10]}), .I1 ({Key_s1[10], Key_s0[10]}), .I2 ({Key_s1[74], Key_s0[74]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1034, AddRoundKeyOutput[10]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[11], Input_s0[11]}), .I1 ({Key_s1[11], Key_s0[11]}), .I2 ({Key_s1[75], Key_s0[75]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1037, AddRoundKeyOutput[11]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[12], Input_s0[12]}), .I1 ({Key_s1[12], Key_s0[12]}), .I2 ({Key_s1[76], Key_s0[76]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1040, AddRoundKeyOutput[12]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[13], Input_s0[13]}), .I1 ({Key_s1[13], Key_s0[13]}), .I2 ({Key_s1[77], Key_s0[77]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1043, AddRoundKeyOutput[13]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[14], Input_s0[14]}), .I1 ({Key_s1[14], Key_s0[14]}), .I2 ({Key_s1[78], Key_s0[78]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1046, AddRoundKeyOutput[14]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[15], Input_s0[15]}), .I1 ({Key_s1[15], Key_s0[15]}), .I2 ({Key_s1[79], Key_s0[79]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1049, AddRoundKeyOutput[15]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[16], Input_s0[16]}), .I1 ({Key_s1[16], Key_s0[16]}), .I2 ({Key_s1[80], Key_s0[80]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_763, Feedback[16]}), .O ({new_AGEMA_signal_1052, AddRoundKeyOutput[16]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[17], Input_s0[17]}), .I1 ({Key_s1[17], Key_s0[17]}), .I2 ({Key_s1[81], Key_s0[81]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_764, Feedback[17]}), .O ({new_AGEMA_signal_1055, AddRoundKeyOutput[17]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[18], Input_s0[18]}), .I1 ({Key_s1[18], Key_s0[18]}), .I2 ({Key_s1[82], Key_s0[82]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_765, Feedback[18]}), .O ({new_AGEMA_signal_1058, AddRoundKeyOutput[18]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[19], Input_s0[19]}), .I1 ({Key_s1[19], Key_s0[19]}), .I2 ({Key_s1[83], Key_s0[83]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_766, Feedback[19]}), .O ({new_AGEMA_signal_1061, AddRoundKeyOutput[19]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[1], Input_s0[1]}), .I1 ({Key_s1[1], Key_s0[1]}), .I2 ({Key_s1[65], Key_s0[65]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1064, AddRoundKeyOutput[1]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[20], Input_s0[20]}), .I1 ({Key_s1[20], Key_s0[20]}), .I2 ({Key_s1[84], Key_s0[84]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_771, Feedback[20]}), .O ({new_AGEMA_signal_1067, AddRoundKeyOutput[20]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[21], Input_s0[21]}), .I1 ({Key_s1[21], Key_s0[21]}), .I2 ({Key_s1[85], Key_s0[85]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_772, Feedback[21]}), .O ({new_AGEMA_signal_1070, AddRoundKeyOutput[21]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[22], Input_s0[22]}), .I1 ({Key_s1[22], Key_s0[22]}), .I2 ({Key_s1[86], Key_s0[86]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_773, Feedback[22]}), .O ({new_AGEMA_signal_1073, AddRoundKeyOutput[22]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[23], Input_s0[23]}), .I1 ({Key_s1[23], Key_s0[23]}), .I2 ({Key_s1[87], Key_s0[87]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_774, Feedback[23]}), .O ({new_AGEMA_signal_1076, AddRoundKeyOutput[23]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[24], Input_s0[24]}), .I1 ({Key_s1[24], Key_s0[24]}), .I2 ({Key_s1[88], Key_s0[88]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_779, Feedback[24]}), .O ({new_AGEMA_signal_1079, AddRoundKeyOutput[24]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[25], Input_s0[25]}), .I1 ({Key_s1[25], Key_s0[25]}), .I2 ({Key_s1[89], Key_s0[89]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_780, Feedback[25]}), .O ({new_AGEMA_signal_1082, AddRoundKeyOutput[25]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[26], Input_s0[26]}), .I1 ({Key_s1[26], Key_s0[26]}), .I2 ({Key_s1[90], Key_s0[90]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_781, Feedback[26]}), .O ({new_AGEMA_signal_1085, AddRoundKeyOutput[26]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[27], Input_s0[27]}), .I1 ({Key_s1[27], Key_s0[27]}), .I2 ({Key_s1[91], Key_s0[91]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_782, Feedback[27]}), .O ({new_AGEMA_signal_1088, AddRoundKeyOutput[27]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[28], Input_s0[28]}), .I1 ({Key_s1[28], Key_s0[28]}), .I2 ({Key_s1[92], Key_s0[92]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_787, Feedback[28]}), .O ({new_AGEMA_signal_1091, AddRoundKeyOutput[28]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[29], Input_s0[29]}), .I1 ({Key_s1[29], Key_s0[29]}), .I2 ({Key_s1[93], Key_s0[93]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_788, Feedback[29]}), .O ({new_AGEMA_signal_1094, AddRoundKeyOutput[29]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[2], Input_s0[2]}), .I1 ({Key_s1[2], Key_s0[2]}), .I2 ({Key_s1[66], Key_s0[66]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1097, AddRoundKeyOutput[2]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[30], Input_s0[30]}), .I1 ({Key_s1[30], Key_s0[30]}), .I2 ({Key_s1[94], Key_s0[94]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_789, Feedback[30]}), .O ({new_AGEMA_signal_1100, AddRoundKeyOutput[30]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[31], Input_s0[31]}), .I1 ({Key_s1[31], Key_s0[31]}), .I2 ({Key_s1[95], Key_s0[95]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_790, Feedback[31]}), .O ({new_AGEMA_signal_1103, AddRoundKeyOutput[31]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[3], Input_s0[3]}), .I1 ({Key_s1[3], Key_s0[3]}), .I2 ({Key_s1[67], Key_s0[67]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1106, AddRoundKeyOutput[3]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[4], Input_s0[4]}), .I1 ({Key_s1[4], Key_s0[4]}), .I2 ({Key_s1[68], Key_s0[68]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1109, AddRoundKeyOutput[4]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[5], Input_s0[5]}), .I1 ({Key_s1[5], Key_s0[5]}), .I2 ({Key_s1[69], Key_s0[69]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1112, AddRoundKeyOutput[5]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[6], Input_s0[6]}), .I1 ({Key_s1[6], Key_s0[6]}), .I2 ({Key_s1[70], Key_s0[70]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1115, AddRoundKeyOutput[6]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[7], Input_s0[7]}), .I1 ({Key_s1[7], Key_s0[7]}), .I2 ({Key_s1[71], Key_s0[71]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1118, AddRoundKeyOutput[7]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[8], Input_s0[8]}), .I1 ({Key_s1[8], Key_s0[8]}), .I2 ({Key_s1[72], Key_s0[72]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1121, AddRoundKeyOutput[8]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[9], Input_s0[9]}), .I1 ({Key_s1[9], Key_s0[9]}), .I2 ({Key_s1[73], Key_s0[73]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1124, AddRoundKeyOutput[9]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_935, N55}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [5]}), .I3 ({new_AGEMA_signal_932, N54}), .I4 ({new_AGEMA_signal_821, Feedback[46]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1125, AddRoundKeyOutput[46]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_941, N58}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [4]}), .I3 ({new_AGEMA_signal_938, N57}), .I4 ({new_AGEMA_signal_820, Feedback[45]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1126, AddRoundKeyOutput[45]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[32], Input_s0[32]}), .I1 ({Input_s1[0], Input_s0[0]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_857, N4}), .I4 ({new_AGEMA_signal_795, Feedback[32]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1128, AddRoundKeyOutput[32]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[33], Input_s0[33]}), .I1 ({Input_s1[1], Input_s0[1]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_860, N6}), .I4 ({new_AGEMA_signal_796, Feedback[33]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1130, AddRoundKeyOutput[33]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[34], Input_s0[34]}), .I1 ({Input_s1[2], Input_s0[2]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_863, N8}), .I4 ({new_AGEMA_signal_797, Feedback[34]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1132, AddRoundKeyOutput[34]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[35], Input_s0[35]}), .I1 ({Input_s1[3], Input_s0[3]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_866, N10}), .I4 ({new_AGEMA_signal_798, Feedback[35]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1134, AddRoundKeyOutput[35]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[36], Input_s0[36]}), .I1 ({Input_s1[4], Input_s0[4]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_869, N12}), .I4 ({new_AGEMA_signal_803, Feedback[36]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1136, AddRoundKeyOutput[36]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[37], Input_s0[37]}), .I1 ({Input_s1[5], Input_s0[5]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_872, N14}), .I4 ({new_AGEMA_signal_804, Feedback[37]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1138, AddRoundKeyOutput[37]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[38], Input_s0[38]}), .I1 ({Input_s1[6], Input_s0[6]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_875, N16}), .I4 ({new_AGEMA_signal_805, Feedback[38]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1140, AddRoundKeyOutput[38]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[39], Input_s0[39]}), .I1 ({Input_s1[7], Input_s0[7]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_878, N18}), .I4 ({new_AGEMA_signal_806, Feedback[39]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1142, AddRoundKeyOutput[39]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyConstXOR/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[43], Input_s0[43]}), .I1 ({Input_s1[11], Input_s0[11]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_881, N20}), .I4 ({new_AGEMA_signal_814, Feedback[43]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1144, AddRoundKeyOutput[43]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_975, N75}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_884, N22}), .I3 ({new_AGEMA_signal_827, Feedback[48]}), .I4 ({new_AGEMA_signal_763, Feedback[16]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1145, AddRoundKeyOutput[48]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_979, N77}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_887, N24}), .I3 ({new_AGEMA_signal_828, Feedback[49]}), .I4 ({new_AGEMA_signal_764, Feedback[17]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1146, AddRoundKeyOutput[49]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_983, N79}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_890, N26}), .I3 ({new_AGEMA_signal_829, Feedback[50]}), .I4 ({new_AGEMA_signal_765, Feedback[18]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1147, AddRoundKeyOutput[50]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_987, N81}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_893, N28}), .I3 ({new_AGEMA_signal_830, Feedback[51]}), .I4 ({new_AGEMA_signal_766, Feedback[19]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1148, AddRoundKeyOutput[51]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_991, N83}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_896, N30}), .I3 ({new_AGEMA_signal_835, Feedback[52]}), .I4 ({new_AGEMA_signal_771, Feedback[20]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1149, AddRoundKeyOutput[52]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_995, N85}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_899, N32}), .I3 ({new_AGEMA_signal_836, Feedback[53]}), .I4 ({new_AGEMA_signal_772, Feedback[21]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1150, AddRoundKeyOutput[53]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_999, N87}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_902, N34}), .I3 ({new_AGEMA_signal_837, Feedback[54]}), .I4 ({new_AGEMA_signal_773, Feedback[22]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1151, AddRoundKeyOutput[54]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1003, N89}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_905, N36}), .I3 ({new_AGEMA_signal_838, Feedback[55]}), .I4 ({new_AGEMA_signal_774, Feedback[23]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1152, AddRoundKeyOutput[55]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1006, N91}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_908, N38}), .I3 ({new_AGEMA_signal_843, Feedback[56]}), .I4 ({new_AGEMA_signal_779, Feedback[24]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1153, AddRoundKeyOutput[56]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1009, N93}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_911, N40}), .I3 ({new_AGEMA_signal_844, Feedback[57]}), .I4 ({new_AGEMA_signal_780, Feedback[25]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1154, AddRoundKeyOutput[57]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1012, N95}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_914, N42}), .I3 ({new_AGEMA_signal_845, Feedback[58]}), .I4 ({new_AGEMA_signal_781, Feedback[26]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1155, AddRoundKeyOutput[58]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1016, N97}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_917, N44}), .I3 ({new_AGEMA_signal_846, Feedback[59]}), .I4 ({new_AGEMA_signal_782, Feedback[27]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1156, AddRoundKeyOutput[59]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1019, N99}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_920, N46}), .I3 ({new_AGEMA_signal_851, Feedback[60]}), .I4 ({new_AGEMA_signal_787, Feedback[28]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1157, AddRoundKeyOutput[60]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1022, N101}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_923, N48}), .I3 ({new_AGEMA_signal_852, Feedback[61]}), .I4 ({new_AGEMA_signal_788, Feedback[29]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1158, AddRoundKeyOutput[61]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1025, N103}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_926, N50}), .I3 ({new_AGEMA_signal_853, Feedback[62]}), .I4 ({new_AGEMA_signal_789, Feedback[30]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1159, AddRoundKeyOutput[62]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1028, N105}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_929, N52}), .I3 ({new_AGEMA_signal_854, Feedback[63]}), .I4 ({new_AGEMA_signal_790, Feedback[31]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1160, AddRoundKeyOutput[63]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_947, N61}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [6]}), .I3 ({new_AGEMA_signal_944, N60}), .I4 ({new_AGEMA_signal_822, Feedback[47]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1161, AddRoundKeyOutput[47]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h4774744774474774 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_953, N64}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [3]}), .I3 ({new_AGEMA_signal_950, N63}), .I4 ({new_AGEMA_signal_819, Feedback[44]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1162, AddRoundKeyOutput[44]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_959, N67}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [2]}), .I3 ({new_AGEMA_signal_956, N66}), .I4 ({new_AGEMA_signal_813, Feedback[42]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1163, AddRoundKeyOutput[42]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_965, N70}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [1]}), .I3 ({new_AGEMA_signal_962, N69}), .I4 ({new_AGEMA_signal_812, Feedback[41]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1164, AddRoundKeyOutput[41]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h4774744774474774 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_971, N73}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [0]}), .I3 ({new_AGEMA_signal_968, N72}), .I4 ({new_AGEMA_signal_811, Feedback[40]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1165, AddRoundKeyOutput[40]}) ) ;

    /* register cells */
    FD done_2 ( .D (done_internal), .C (clk_gated), .Q (done) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_6 ( .D (\FSMUpdate [6]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [6]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_5 ( .D (\FSM [6]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [5]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_4 ( .D (\FSM [5]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [4]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_3 ( .D (\FSM [4]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [3]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_2 ( .D (\FSMUpdate [2]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [2]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_1 ( .D (\FSM [2]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [1]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_0 ( .D (\FSM [1]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [0]) ) ;
    FD #( .INIT ( 1'b0 ) ) \selectsRegInst/s_current_state_0 ( .D (selectsNext[0]), .C (clk_gated), .Q (\selectsRegInst/s_current_state [0]) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_63 ( .D ({new_AGEMA_signal_1160, AddRoundKeyOutput[63]}), .clk (clk_gated), .Q ({Output_s1[63], Output_s0[63]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_62 ( .D ({new_AGEMA_signal_1159, AddRoundKeyOutput[62]}), .clk (clk_gated), .Q ({Output_s1[62], Output_s0[62]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_61 ( .D ({new_AGEMA_signal_1158, AddRoundKeyOutput[61]}), .clk (clk_gated), .Q ({Output_s1[61], Output_s0[61]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_60 ( .D ({new_AGEMA_signal_1157, AddRoundKeyOutput[60]}), .clk (clk_gated), .Q ({Output_s1[60], Output_s0[60]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_59 ( .D ({new_AGEMA_signal_1156, AddRoundKeyOutput[59]}), .clk (clk_gated), .Q ({Output_s1[59], Output_s0[59]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_58 ( .D ({new_AGEMA_signal_1155, AddRoundKeyOutput[58]}), .clk (clk_gated), .Q ({Output_s1[58], Output_s0[58]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_57 ( .D ({new_AGEMA_signal_1154, AddRoundKeyOutput[57]}), .clk (clk_gated), .Q ({Output_s1[57], Output_s0[57]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_56 ( .D ({new_AGEMA_signal_1153, AddRoundKeyOutput[56]}), .clk (clk_gated), .Q ({Output_s1[56], Output_s0[56]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_55 ( .D ({new_AGEMA_signal_1152, AddRoundKeyOutput[55]}), .clk (clk_gated), .Q ({Output_s1[55], Output_s0[55]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_54 ( .D ({new_AGEMA_signal_1151, AddRoundKeyOutput[54]}), .clk (clk_gated), .Q ({Output_s1[54], Output_s0[54]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_53 ( .D ({new_AGEMA_signal_1150, AddRoundKeyOutput[53]}), .clk (clk_gated), .Q ({Output_s1[53], Output_s0[53]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_52 ( .D ({new_AGEMA_signal_1149, AddRoundKeyOutput[52]}), .clk (clk_gated), .Q ({Output_s1[52], Output_s0[52]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_51 ( .D ({new_AGEMA_signal_1148, AddRoundKeyOutput[51]}), .clk (clk_gated), .Q ({Output_s1[51], Output_s0[51]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_50 ( .D ({new_AGEMA_signal_1147, AddRoundKeyOutput[50]}), .clk (clk_gated), .Q ({Output_s1[50], Output_s0[50]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_49 ( .D ({new_AGEMA_signal_1146, AddRoundKeyOutput[49]}), .clk (clk_gated), .Q ({Output_s1[49], Output_s0[49]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_48 ( .D ({new_AGEMA_signal_1145, AddRoundKeyOutput[48]}), .clk (clk_gated), .Q ({Output_s1[48], Output_s0[48]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_47 ( .D ({new_AGEMA_signal_1161, AddRoundKeyOutput[47]}), .clk (clk_gated), .Q ({Output_s1[47], Output_s0[47]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_46 ( .D ({new_AGEMA_signal_1125, AddRoundKeyOutput[46]}), .clk (clk_gated), .Q ({Output_s1[46], Output_s0[46]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_45 ( .D ({new_AGEMA_signal_1126, AddRoundKeyOutput[45]}), .clk (clk_gated), .Q ({Output_s1[45], Output_s0[45]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_44 ( .D ({new_AGEMA_signal_1162, AddRoundKeyOutput[44]}), .clk (clk_gated), .Q ({Output_s1[44], Output_s0[44]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_43 ( .D ({new_AGEMA_signal_1144, AddRoundKeyOutput[43]}), .clk (clk_gated), .Q ({Output_s1[43], Output_s0[43]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_42 ( .D ({new_AGEMA_signal_1163, AddRoundKeyOutput[42]}), .clk (clk_gated), .Q ({Output_s1[42], Output_s0[42]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_41 ( .D ({new_AGEMA_signal_1164, AddRoundKeyOutput[41]}), .clk (clk_gated), .Q ({Output_s1[41], Output_s0[41]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_40 ( .D ({new_AGEMA_signal_1165, AddRoundKeyOutput[40]}), .clk (clk_gated), .Q ({Output_s1[40], Output_s0[40]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_39 ( .D ({new_AGEMA_signal_1142, AddRoundKeyOutput[39]}), .clk (clk_gated), .Q ({Output_s1[39], Output_s0[39]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_38 ( .D ({new_AGEMA_signal_1140, AddRoundKeyOutput[38]}), .clk (clk_gated), .Q ({Output_s1[38], Output_s0[38]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_37 ( .D ({new_AGEMA_signal_1138, AddRoundKeyOutput[37]}), .clk (clk_gated), .Q ({Output_s1[37], Output_s0[37]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_36 ( .D ({new_AGEMA_signal_1136, AddRoundKeyOutput[36]}), .clk (clk_gated), .Q ({Output_s1[36], Output_s0[36]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_35 ( .D ({new_AGEMA_signal_1134, AddRoundKeyOutput[35]}), .clk (clk_gated), .Q ({Output_s1[35], Output_s0[35]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_34 ( .D ({new_AGEMA_signal_1132, AddRoundKeyOutput[34]}), .clk (clk_gated), .Q ({Output_s1[34], Output_s0[34]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_33 ( .D ({new_AGEMA_signal_1130, AddRoundKeyOutput[33]}), .clk (clk_gated), .Q ({Output_s1[33], Output_s0[33]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_32 ( .D ({new_AGEMA_signal_1128, AddRoundKeyOutput[32]}), .clk (clk_gated), .Q ({Output_s1[32], Output_s0[32]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_31 ( .D ({new_AGEMA_signal_1103, AddRoundKeyOutput[31]}), .clk (clk_gated), .Q ({Output_s1[31], Output_s0[31]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_30 ( .D ({new_AGEMA_signal_1100, AddRoundKeyOutput[30]}), .clk (clk_gated), .Q ({Output_s1[30], Output_s0[30]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_29 ( .D ({new_AGEMA_signal_1094, AddRoundKeyOutput[29]}), .clk (clk_gated), .Q ({Output_s1[29], Output_s0[29]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_28 ( .D ({new_AGEMA_signal_1091, AddRoundKeyOutput[28]}), .clk (clk_gated), .Q ({Output_s1[28], Output_s0[28]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_27 ( .D ({new_AGEMA_signal_1088, AddRoundKeyOutput[27]}), .clk (clk_gated), .Q ({Output_s1[27], Output_s0[27]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_26 ( .D ({new_AGEMA_signal_1085, AddRoundKeyOutput[26]}), .clk (clk_gated), .Q ({Output_s1[26], Output_s0[26]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_25 ( .D ({new_AGEMA_signal_1082, AddRoundKeyOutput[25]}), .clk (clk_gated), .Q ({Output_s1[25], Output_s0[25]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_24 ( .D ({new_AGEMA_signal_1079, AddRoundKeyOutput[24]}), .clk (clk_gated), .Q ({Output_s1[24], Output_s0[24]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_23 ( .D ({new_AGEMA_signal_1076, AddRoundKeyOutput[23]}), .clk (clk_gated), .Q ({Output_s1[23], Output_s0[23]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_22 ( .D ({new_AGEMA_signal_1073, AddRoundKeyOutput[22]}), .clk (clk_gated), .Q ({Output_s1[22], Output_s0[22]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_21 ( .D ({new_AGEMA_signal_1070, AddRoundKeyOutput[21]}), .clk (clk_gated), .Q ({Output_s1[21], Output_s0[21]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_20 ( .D ({new_AGEMA_signal_1067, AddRoundKeyOutput[20]}), .clk (clk_gated), .Q ({Output_s1[20], Output_s0[20]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_19 ( .D ({new_AGEMA_signal_1061, AddRoundKeyOutput[19]}), .clk (clk_gated), .Q ({Output_s1[19], Output_s0[19]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_18 ( .D ({new_AGEMA_signal_1058, AddRoundKeyOutput[18]}), .clk (clk_gated), .Q ({Output_s1[18], Output_s0[18]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_17 ( .D ({new_AGEMA_signal_1055, AddRoundKeyOutput[17]}), .clk (clk_gated), .Q ({Output_s1[17], Output_s0[17]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_16 ( .D ({new_AGEMA_signal_1052, AddRoundKeyOutput[16]}), .clk (clk_gated), .Q ({Output_s1[16], Output_s0[16]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_15 ( .D ({new_AGEMA_signal_1049, AddRoundKeyOutput[15]}), .clk (clk_gated), .Q ({Output_s1[15], Output_s0[15]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_14 ( .D ({new_AGEMA_signal_1046, AddRoundKeyOutput[14]}), .clk (clk_gated), .Q ({Output_s1[14], Output_s0[14]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_13 ( .D ({new_AGEMA_signal_1043, AddRoundKeyOutput[13]}), .clk (clk_gated), .Q ({Output_s1[13], Output_s0[13]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_12 ( .D ({new_AGEMA_signal_1040, AddRoundKeyOutput[12]}), .clk (clk_gated), .Q ({Output_s1[12], Output_s0[12]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_11 ( .D ({new_AGEMA_signal_1037, AddRoundKeyOutput[11]}), .clk (clk_gated), .Q ({Output_s1[11], Output_s0[11]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_10 ( .D ({new_AGEMA_signal_1034, AddRoundKeyOutput[10]}), .clk (clk_gated), .Q ({Output_s1[10], Output_s0[10]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_9 ( .D ({new_AGEMA_signal_1124, AddRoundKeyOutput[9]}), .clk (clk_gated), .Q ({Output_s1[9], Output_s0[9]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_8 ( .D ({new_AGEMA_signal_1121, AddRoundKeyOutput[8]}), .clk (clk_gated), .Q ({Output_s1[8], Output_s0[8]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_7 ( .D ({new_AGEMA_signal_1118, AddRoundKeyOutput[7]}), .clk (clk_gated), .Q ({Output_s1[7], Output_s0[7]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_6 ( .D ({new_AGEMA_signal_1115, AddRoundKeyOutput[6]}), .clk (clk_gated), .Q ({Output_s1[6], Output_s0[6]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_5 ( .D ({new_AGEMA_signal_1112, AddRoundKeyOutput[5]}), .clk (clk_gated), .Q ({Output_s1[5], Output_s0[5]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_4 ( .D ({new_AGEMA_signal_1109, AddRoundKeyOutput[4]}), .clk (clk_gated), .Q ({Output_s1[4], Output_s0[4]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_3 ( .D ({new_AGEMA_signal_1106, AddRoundKeyOutput[3]}), .clk (clk_gated), .Q ({Output_s1[3], Output_s0[3]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_2 ( .D ({new_AGEMA_signal_1097, AddRoundKeyOutput[2]}), .clk (clk_gated), .Q ({Output_s1[2], Output_s0[2]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_1 ( .D ({new_AGEMA_signal_1064, AddRoundKeyOutput[1]}), .clk (clk_gated), .Q ({Output_s1[1], Output_s0[1]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_0 ( .D ({new_AGEMA_signal_1031, AddRoundKeyOutput[0]}), .clk (clk_gated), .Q ({Output_s1[0], Output_s0[0]}) ) ;
endmodule
