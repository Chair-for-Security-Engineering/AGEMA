/* modified netlist. Source: module AES in file AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_AIG_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [135:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_416 ;
    wire signal_418 ;
    wire signal_420 ;
    wire signal_422 ;
    wire signal_424 ;
    wire signal_426 ;
    wire signal_428 ;
    wire signal_430 ;
    wire signal_432 ;
    wire signal_434 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_440 ;
    wire signal_442 ;
    wire signal_444 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_450 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_456 ;
    wire signal_458 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_588 ;
    wire signal_590 ;
    wire signal_592 ;
    wire signal_594 ;
    wire signal_596 ;
    wire signal_598 ;
    wire signal_600 ;
    wire signal_602 ;
    wire signal_604 ;
    wire signal_606 ;
    wire signal_608 ;
    wire signal_610 ;
    wire signal_612 ;
    wire signal_614 ;
    wire signal_616 ;
    wire signal_618 ;
    wire signal_620 ;
    wire signal_622 ;
    wire signal_624 ;
    wire signal_626 ;
    wire signal_628 ;
    wire signal_630 ;
    wire signal_632 ;
    wire signal_634 ;
    wire signal_636 ;
    wire signal_638 ;
    wire signal_640 ;
    wire signal_642 ;
    wire signal_644 ;
    wire signal_646 ;
    wire signal_648 ;
    wire signal_650 ;
    wire signal_652 ;
    wire signal_654 ;
    wire signal_656 ;
    wire signal_658 ;
    wire signal_660 ;
    wire signal_662 ;
    wire signal_664 ;
    wire signal_666 ;
    wire signal_668 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_788 ;
    wire signal_908 ;
    wire signal_1028 ;
    wire signal_1148 ;
    wire signal_1153 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1297 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1303 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1309 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1315 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1321 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1327 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1333 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1339 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1345 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1351 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1357 ;
    wire signal_1359 ;
    wire signal_1361 ;
    wire signal_1363 ;
    wire signal_1365 ;
    wire signal_1367 ;
    wire signal_1369 ;
    wire signal_1371 ;
    wire signal_1373 ;
    wire signal_1375 ;
    wire signal_1377 ;
    wire signal_1379 ;
    wire signal_1381 ;
    wire signal_1383 ;
    wire signal_1385 ;
    wire signal_1387 ;
    wire signal_1389 ;
    wire signal_1391 ;
    wire signal_1393 ;
    wire signal_1395 ;
    wire signal_1397 ;
    wire signal_1399 ;
    wire signal_1401 ;
    wire signal_1403 ;
    wire signal_1405 ;
    wire signal_1407 ;
    wire signal_1409 ;
    wire signal_1411 ;
    wire signal_1413 ;
    wire signal_1415 ;
    wire signal_1417 ;
    wire signal_1419 ;
    wire signal_1421 ;
    wire signal_1423 ;
    wire signal_1425 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1431 ;
    wire signal_1433 ;
    wire signal_1435 ;
    wire signal_1437 ;
    wire signal_1439 ;
    wire signal_1441 ;
    wire signal_1443 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1449 ;
    wire signal_1451 ;
    wire signal_1453 ;
    wire signal_1455 ;
    wire signal_1457 ;
    wire signal_1459 ;
    wire signal_1461 ;
    wire signal_1463 ;
    wire signal_1465 ;
    wire signal_1467 ;
    wire signal_1469 ;
    wire signal_1471 ;
    wire signal_1473 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1479 ;
    wire signal_1481 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2303 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3433 ;
    wire signal_3435 ;
    wire signal_3437 ;
    wire signal_3439 ;
    wire signal_3441 ;
    wire signal_3443 ;
    wire signal_3445 ;
    wire signal_3447 ;
    wire signal_3449 ;
    wire signal_3451 ;
    wire signal_3453 ;
    wire signal_3455 ;
    wire signal_3457 ;
    wire signal_3459 ;
    wire signal_3461 ;
    wire signal_3463 ;
    wire signal_3465 ;
    wire signal_3467 ;
    wire signal_3469 ;
    wire signal_3471 ;
    wire signal_3473 ;
    wire signal_3475 ;
    wire signal_3477 ;
    wire signal_3479 ;
    wire signal_3481 ;
    wire signal_3483 ;
    wire signal_3485 ;
    wire signal_3487 ;
    wire signal_3489 ;
    wire signal_3491 ;
    wire signal_3493 ;
    wire signal_3495 ;
    wire signal_3497 ;
    wire signal_3499 ;
    wire signal_3501 ;
    wire signal_3503 ;
    wire signal_3505 ;
    wire signal_3507 ;
    wire signal_3509 ;
    wire signal_3511 ;
    wire signal_3513 ;
    wire signal_3515 ;
    wire signal_3517 ;
    wire signal_3519 ;
    wire signal_3521 ;
    wire signal_3523 ;
    wire signal_3525 ;
    wire signal_3527 ;
    wire signal_3529 ;
    wire signal_3531 ;
    wire signal_3533 ;
    wire signal_3535 ;
    wire signal_3537 ;
    wire signal_3539 ;
    wire signal_3541 ;
    wire signal_3543 ;
    wire signal_3545 ;
    wire signal_3547 ;
    wire signal_3549 ;
    wire signal_3551 ;
    wire signal_3553 ;
    wire signal_3555 ;
    wire signal_3557 ;
    wire signal_3559 ;
    wire signal_3561 ;
    wire signal_3563 ;
    wire signal_3565 ;
    wire signal_3567 ;
    wire signal_3569 ;
    wire signal_3571 ;
    wire signal_3573 ;
    wire signal_3575 ;
    wire signal_3577 ;
    wire signal_3579 ;
    wire signal_3581 ;
    wire signal_3583 ;
    wire signal_3585 ;
    wire signal_3587 ;
    wire signal_3589 ;
    wire signal_3591 ;
    wire signal_3593 ;
    wire signal_3595 ;
    wire signal_3597 ;
    wire signal_3599 ;
    wire signal_3601 ;
    wire signal_3603 ;
    wire signal_3605 ;
    wire signal_3607 ;
    wire signal_3609 ;
    wire signal_3611 ;
    wire signal_3613 ;
    wire signal_3615 ;
    wire signal_3617 ;
    wire signal_3619 ;
    wire signal_3621 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4284 ;
    wire signal_4286 ;
    wire signal_4288 ;
    wire signal_4290 ;
    wire signal_4292 ;
    wire signal_4294 ;
    wire signal_4296 ;
    wire signal_4298 ;
    wire signal_4300 ;
    wire signal_4302 ;
    wire signal_4304 ;
    wire signal_4306 ;
    wire signal_4308 ;
    wire signal_4310 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4416 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4422 ;
    wire signal_4424 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4430 ;
    wire signal_4432 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4438 ;
    wire signal_4440 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4446 ;
    wire signal_4448 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4454 ;
    wire signal_4456 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4462 ;
    wire signal_4464 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4470 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4590 ;
    wire signal_4592 ;
    wire signal_4594 ;
    wire signal_4596 ;
    wire signal_4598 ;
    wire signal_4600 ;
    wire signal_4602 ;
    wire signal_4604 ;
    wire signal_4606 ;
    wire signal_4608 ;
    wire signal_4610 ;
    wire signal_4612 ;
    wire signal_4614 ;
    wire signal_4616 ;
    wire signal_4618 ;
    wire signal_4620 ;
    wire signal_4622 ;
    wire signal_4624 ;
    wire signal_4626 ;
    wire signal_4628 ;
    wire signal_4630 ;
    wire signal_4632 ;
    wire signal_4634 ;
    wire signal_4636 ;
    wire signal_4638 ;
    wire signal_4640 ;
    wire signal_4642 ;
    wire signal_4644 ;
    wire signal_4646 ;
    wire signal_4648 ;
    wire signal_4650 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4706 ;
    wire signal_4708 ;
    wire signal_4710 ;
    wire signal_4712 ;
    wire signal_4714 ;
    wire signal_4716 ;
    wire signal_4718 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4746 ;
    wire signal_4748 ;
    wire signal_4750 ;
    wire signal_4752 ;
    wire signal_4754 ;
    wire signal_4756 ;
    wire signal_4758 ;
    wire signal_4760 ;
    wire signal_4762 ;
    wire signal_4764 ;
    wire signal_4766 ;
    wire signal_4768 ;
    wire signal_4770 ;
    wire signal_4772 ;
    wire signal_4774 ;
    wire signal_4776 ;
    wire signal_4778 ;
    wire signal_4780 ;
    wire signal_4782 ;
    wire signal_4784 ;
    wire signal_4786 ;
    wire signal_4788 ;
    wire signal_4790 ;
    wire signal_4792 ;
    wire signal_4794 ;
    wire signal_4796 ;
    wire signal_4798 ;
    wire signal_4800 ;
    wire signal_4802 ;
    wire signal_4804 ;
    wire signal_4806 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4830 ;
    wire signal_4832 ;
    wire signal_4834 ;
    wire signal_4836 ;
    wire signal_4838 ;
    wire signal_4840 ;
    wire signal_4842 ;
    wire signal_4844 ;
    wire signal_4846 ;
    wire signal_4848 ;
    wire signal_4850 ;
    wire signal_4852 ;
    wire signal_4854 ;
    wire signal_4856 ;
    wire signal_4858 ;
    wire signal_4860 ;
    wire signal_4862 ;
    wire signal_4864 ;
    wire signal_4866 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4874 ;
    wire signal_4876 ;
    wire signal_4878 ;
    wire signal_4880 ;
    wire signal_4882 ;
    wire signal_4884 ;
    wire signal_4886 ;
    wire signal_4888 ;
    wire signal_4890 ;
    wire signal_4892 ;
    wire signal_4894 ;
    wire signal_4896 ;
    wire signal_4898 ;
    wire signal_4900 ;
    wire signal_4902 ;
    wire signal_4904 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4911 ;
    wire signal_4913 ;
    wire signal_4915 ;
    wire signal_4917 ;
    wire signal_4919 ;
    wire signal_4921 ;
    wire signal_4923 ;
    wire signal_5060 ;

    /* cells in depth 0 */
    AND2_X1 cell_0 ( .A1 (signal_396), .A2 (signal_395), .ZN (signal_393) ) ;
    NOR2_X1 cell_1 ( .A1 (signal_411), .A2 (signal_400), .ZN (signal_394) ) ;
    AND2_X1 cell_2 ( .A1 (signal_2273), .A2 (signal_394), .ZN (done) ) ;
    INV_X1 cell_3 ( .A (signal_2270), .ZN (signal_411) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_396) ) ;
    INV_X1 cell_5 ( .A (signal_2271), .ZN (signal_397) ) ;
    NAND2_X1 cell_6 ( .A1 (signal_2272), .A2 (signal_397), .ZN (signal_400) ) ;
    NOR2_X1 cell_7 ( .A1 (done), .A2 (signal_2274), .ZN (signal_395) ) ;
    INV_X1 cell_8 ( .A (signal_2272), .ZN (signal_406) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_406), .A2 (signal_397), .ZN (signal_398) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_2273), .A2 (signal_398), .ZN (signal_2141) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_2273), .A2 (signal_2270), .ZN (signal_409) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_409), .A2 (signal_398), .ZN (signal_2140) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_2270), .A2 (signal_400), .ZN (signal_399) ) ;
    NOR2_X1 cell_14 ( .A1 (signal_411), .A2 (signal_398), .ZN (signal_405) ) ;
    MUX2_X1 cell_15 ( .S (signal_2273), .A (signal_399), .B (signal_405), .Z (signal_2139) ) ;
    INV_X1 cell_16 ( .A (signal_2273), .ZN (signal_401) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_401), .A2 (signal_400), .ZN (signal_402) ) ;
    MUX2_X1 cell_18 ( .S (signal_2270), .A (signal_402), .B (signal_2141), .Z (signal_2138) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_2271), .A2 (signal_409), .ZN (signal_403) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_2272), .A2 (signal_403), .ZN (signal_404) ) ;
    OR2_X1 cell_21 ( .A1 (signal_405), .A2 (signal_404), .ZN (signal_2137) ) ;
    XNOR2_X1 cell_22 ( .A (signal_2271), .B (signal_2270), .ZN (signal_408) ) ;
    NAND2_X1 cell_23 ( .A1 (signal_2273), .A2 (signal_406), .ZN (signal_407) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_2136) ) ;
    INV_X1 cell_25 ( .A (signal_409), .ZN (signal_410) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_2272), .A2 (signal_2271), .ZN (signal_412) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_410), .A2 (signal_412), .ZN (signal_2135) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_2273), .A2 (signal_411), .ZN (signal_413) ) ;
    NOR2_X1 cell_29 ( .A1 (signal_413), .A2 (signal_412), .ZN (signal_2134) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_30 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_2921, signal_1793}), .c ({signal_2922, signal_1681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_31 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_2924, signal_2065}), .c ({signal_2925, signal_1709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_32 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_2927, signal_2064}), .c ({signal_2928, signal_1708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_33 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_2930, signal_2063}), .c ({signal_2931, signal_1707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_34 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({signal_2933, signal_2062}), .c ({signal_2934, signal_1706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_35 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_2936, signal_2061}), .c ({signal_2937, signal_1737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_36 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_2939, signal_2060}), .c ({signal_2940, signal_1736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_37 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_2942, signal_2059}), .c ({signal_2943, signal_1735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_38 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({signal_2945, signal_2058}), .c ({signal_2946, signal_1734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_39 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_2948, signal_2057}), .c ({signal_2949, signal_1733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_40 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_2951, signal_2056}), .c ({signal_2952, signal_1732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_41 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({signal_2954, signal_1799}), .c ({signal_2955, signal_1703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_42 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_2957, signal_2055}), .c ({signal_2958, signal_1731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_43 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({signal_2960, signal_2054}), .c ({signal_2961, signal_1730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_44 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_2963, signal_2053}), .c ({signal_2964, signal_1761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_45 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({signal_2966, signal_2052}), .c ({signal_2967, signal_1760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_46 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({signal_2969, signal_2051}), .c ({signal_2970, signal_1759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_47 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({signal_2972, signal_2050}), .c ({signal_2973, signal_1758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_48 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({signal_2975, signal_2049}), .c ({signal_2976, signal_1757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_49 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({signal_2978, signal_2048}), .c ({signal_2979, signal_1756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_50 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({signal_2981, signal_2047}), .c ({signal_2982, signal_1755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_51 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({signal_2984, signal_2046}), .c ({signal_2985, signal_1754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_52 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({signal_2987, signal_1798}), .c ({signal_2988, signal_1702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_53 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2990, signal_2045}), .c ({signal_2991, signal_1657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_54 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2993, signal_2044}), .c ({signal_2994, signal_1656}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_55 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2996, signal_2043}), .c ({signal_2997, signal_1655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_56 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2999, signal_2042}), .c ({signal_3000, signal_1654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_57 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_3002, signal_2041}), .c ({signal_3003, signal_1653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_58 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_3005, signal_2040}), .c ({signal_3006, signal_1652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_59 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_3008, signal_2039}), .c ({signal_3009, signal_1651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_60 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_3011, signal_2038}), .c ({signal_3012, signal_1650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_61 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({signal_3014, signal_1797}), .c ({signal_3015, signal_1701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_62 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({signal_3017, signal_1796}), .c ({signal_3018, signal_1700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_63 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({signal_3020, signal_1795}), .c ({signal_3021, signal_1699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_64 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({signal_3023, signal_1794}), .c ({signal_3024, signal_1698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_65 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_3026, signal_1809}), .c ({signal_3027, signal_1729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_66 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({signal_3029, signal_1808}), .c ({signal_3030, signal_1728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_67 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({signal_3032, signal_1807}), .c ({signal_3033, signal_1727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_68 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({signal_3035, signal_1806}), .c ({signal_3036, signal_1726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_69 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_3038, signal_1792}), .c ({signal_3039, signal_1680}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_70 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({signal_3041, signal_1805}), .c ({signal_3042, signal_1725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_71 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({signal_3044, signal_1804}), .c ({signal_3045, signal_1724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_72 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({signal_3047, signal_1803}), .c ({signal_3048, signal_1723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_73 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({signal_3050, signal_1802}), .c ({signal_3051, signal_1722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_74 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_3053, signal_1785}), .c ({signal_3054, signal_1753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_75 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_3056, signal_1784}), .c ({signal_3057, signal_1752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_76 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_3059, signal_1783}), .c ({signal_3060, signal_1751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_77 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_3062, signal_1782}), .c ({signal_3063, signal_1750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_78 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_3065, signal_1781}), .c ({signal_3066, signal_1749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_79 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_3068, signal_1780}), .c ({signal_3069, signal_1748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_80 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_3071, signal_1791}), .c ({signal_3072, signal_1679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_81 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_3074, signal_1779}), .c ({signal_3075, signal_1747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_82 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_3077, signal_1778}), .c ({signal_3078, signal_1746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_83 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_3080, signal_2133}), .c ({signal_3081, signal_1777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_84 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({signal_3083, signal_2132}), .c ({signal_3084, signal_1776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_85 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({signal_3086, signal_2131}), .c ({signal_3087, signal_1775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_86 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({signal_3089, signal_2130}), .c ({signal_3090, signal_1774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_87 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({signal_3092, signal_2129}), .c ({signal_3093, signal_1773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_88 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({signal_3095, signal_2128}), .c ({signal_3096, signal_1772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_89 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({signal_3098, signal_2127}), .c ({signal_3099, signal_1771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_90 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({signal_3101, signal_2126}), .c ({signal_3102, signal_1770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_91 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({signal_3104, signal_1790}), .c ({signal_3105, signal_1678}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_92 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_3107, signal_2125}), .c ({signal_3108, signal_1673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_93 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({signal_3110, signal_2124}), .c ({signal_3111, signal_1672}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_94 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({signal_3113, signal_2123}), .c ({signal_3114, signal_1671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_95 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({signal_3116, signal_2122}), .c ({signal_3117, signal_1670}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_96 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({signal_3119, signal_2121}), .c ({signal_3120, signal_1669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_97 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({signal_3122, signal_2120}), .c ({signal_3123, signal_1668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_98 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({signal_3125, signal_2119}), .c ({signal_3126, signal_1667}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_99 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({signal_3128, signal_2118}), .c ({signal_3129, signal_1666}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_100 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_3131, signal_2117}), .c ({signal_3132, signal_1697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_101 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_3134, signal_2116}), .c ({signal_3135, signal_1696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_102 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_3137, signal_1789}), .c ({signal_3138, signal_1677}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_103 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_3140, signal_2115}), .c ({signal_3141, signal_1695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_104 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({signal_3143, signal_2114}), .c ({signal_3144, signal_1694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_105 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_3146, signal_2113}), .c ({signal_3147, signal_1693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_106 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_3149, signal_2112}), .c ({signal_3150, signal_1692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_107 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_3152, signal_2111}), .c ({signal_3153, signal_1691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_108 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({signal_3155, signal_2110}), .c ({signal_3156, signal_1690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_109 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_3158, signal_2109}), .c ({signal_3159, signal_1721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_110 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_3161, signal_2108}), .c ({signal_3162, signal_1720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_111 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_3164, signal_2107}), .c ({signal_3165, signal_1719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_112 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_3167, signal_2106}), .c ({signal_3168, signal_1718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_113 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_3170, signal_1788}), .c ({signal_3171, signal_1676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_114 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_3173, signal_2105}), .c ({signal_3174, signal_1717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_115 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_3176, signal_2104}), .c ({signal_3177, signal_1716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_116 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_3179, signal_2103}), .c ({signal_3180, signal_1715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_117 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_3182, signal_2102}), .c ({signal_3183, signal_1714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_118 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_3185, signal_2101}), .c ({signal_3186, signal_1745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_119 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({signal_3188, signal_2100}), .c ({signal_3189, signal_1744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_120 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({signal_3191, signal_2099}), .c ({signal_3192, signal_1743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_121 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({signal_3194, signal_2098}), .c ({signal_3195, signal_1742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_122 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({signal_3197, signal_2097}), .c ({signal_3198, signal_1741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_123 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({signal_3200, signal_2096}), .c ({signal_3201, signal_1740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_124 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_3203, signal_1787}), .c ({signal_3204, signal_1675}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_125 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({signal_3206, signal_2095}), .c ({signal_3207, signal_1739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_126 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({signal_3209, signal_2094}), .c ({signal_3210, signal_1738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_127 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_3212, signal_2093}), .c ({signal_3213, signal_1769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_128 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_3215, signal_2092}), .c ({signal_3216, signal_1768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_129 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_3218, signal_2091}), .c ({signal_3219, signal_1767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_130 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({signal_3221, signal_2090}), .c ({signal_3222, signal_1766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_131 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_3224, signal_2089}), .c ({signal_3225, signal_1765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_132 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_3227, signal_2088}), .c ({signal_3228, signal_1764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_133 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_3230, signal_2087}), .c ({signal_3231, signal_1763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_134 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({signal_3233, signal_2086}), .c ({signal_3234, signal_1762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_135 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({signal_3236, signal_1786}), .c ({signal_3237, signal_1674}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_136 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_3239, signal_2085}), .c ({signal_3240, signal_1665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_137 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_3242, signal_2084}), .c ({signal_3243, signal_1664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_138 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_3245, signal_2083}), .c ({signal_3246, signal_1663}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_139 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({signal_3248, signal_2082}), .c ({signal_3249, signal_1662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_140 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_3251, signal_2081}), .c ({signal_3252, signal_1661}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_141 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_3254, signal_2080}), .c ({signal_3255, signal_1660}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_142 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_3257, signal_2079}), .c ({signal_3258, signal_1659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_143 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({signal_3260, signal_2078}), .c ({signal_3261, signal_1658}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_144 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_3263, signal_2077}), .c ({signal_3264, signal_1689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_145 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_3266, signal_2076}), .c ({signal_3267, signal_1688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_146 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_3269, signal_1801}), .c ({signal_3270, signal_1705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_147 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({signal_3272, signal_2075}), .c ({signal_3273, signal_1687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_148 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_3275, signal_2074}), .c ({signal_3276, signal_1686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_149 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_3278, signal_2073}), .c ({signal_3279, signal_1685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_150 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_3281, signal_2072}), .c ({signal_3282, signal_1684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_151 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_3284, signal_2071}), .c ({signal_3285, signal_1683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_152 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_3287, signal_2070}), .c ({signal_3288, signal_1682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_153 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_3290, signal_2069}), .c ({signal_3291, signal_1713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_154 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_3293, signal_2068}), .c ({signal_3294, signal_1712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_155 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_3296, signal_2067}), .c ({signal_3297, signal_1711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_156 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({signal_3299, signal_2066}), .c ({signal_3300, signal_1710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_157 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({signal_3302, signal_1800}), .c ({signal_3303, signal_1704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_256 ( .s (reset), .b ({signal_3336, signal_1617}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_3433, signal_478}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_259 ( .s (reset), .b ({signal_3337, signal_1616}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_3435, signal_480}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_262 ( .s (reset), .b ({signal_3338, signal_1615}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_3437, signal_482}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_265 ( .s (reset), .b ({signal_3339, signal_1614}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_3439, signal_484}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_268 ( .s (reset), .b ({signal_3340, signal_1613}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_3441, signal_486}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_271 ( .s (reset), .b ({signal_3341, signal_1612}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_3443, signal_488}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_274 ( .s (reset), .b ({signal_3342, signal_1611}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_3445, signal_490}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_277 ( .s (reset), .b ({signal_3343, signal_1610}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_3447, signal_492}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_280 ( .s (reset), .b ({signal_3344, signal_1609}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_3449, signal_494}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_283 ( .s (reset), .b ({signal_3345, signal_1608}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_3451, signal_496}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_286 ( .s (reset), .b ({signal_3346, signal_1607}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_3453, signal_498}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_289 ( .s (reset), .b ({signal_3347, signal_1606}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_3455, signal_500}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_292 ( .s (reset), .b ({signal_3348, signal_1605}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_3457, signal_502}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_295 ( .s (reset), .b ({signal_3349, signal_1604}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_3459, signal_504}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_298 ( .s (reset), .b ({signal_3350, signal_1603}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_3461, signal_506}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_301 ( .s (reset), .b ({signal_3351, signal_1602}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_3463, signal_508}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_304 ( .s (reset), .b ({signal_3352, signal_1601}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_3465, signal_510}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_307 ( .s (reset), .b ({signal_3353, signal_1600}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_3467, signal_512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_310 ( .s (reset), .b ({signal_3354, signal_1599}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_3469, signal_514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_313 ( .s (reset), .b ({signal_3355, signal_1598}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_3471, signal_516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_316 ( .s (reset), .b ({signal_3356, signal_1597}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_3473, signal_518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_319 ( .s (reset), .b ({signal_3357, signal_1596}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_3475, signal_520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_322 ( .s (reset), .b ({signal_3358, signal_1595}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_3477, signal_522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_325 ( .s (reset), .b ({signal_3359, signal_1594}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_3479, signal_524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_328 ( .s (reset), .b ({signal_3360, signal_1593}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_3481, signal_526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_331 ( .s (reset), .b ({signal_3361, signal_1592}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_3483, signal_528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_334 ( .s (reset), .b ({signal_3362, signal_1591}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_3485, signal_530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_337 ( .s (reset), .b ({signal_3363, signal_1590}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_3487, signal_532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_340 ( .s (reset), .b ({signal_3364, signal_1589}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_3489, signal_534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_343 ( .s (reset), .b ({signal_3365, signal_1588}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_3491, signal_536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_346 ( .s (reset), .b ({signal_3366, signal_1587}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_3493, signal_538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_349 ( .s (reset), .b ({signal_3367, signal_1586}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_3495, signal_540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_352 ( .s (reset), .b ({signal_3368, signal_1585}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_3497, signal_542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_355 ( .s (reset), .b ({signal_3369, signal_1584}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_3499, signal_544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_358 ( .s (reset), .b ({signal_3370, signal_1583}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_3501, signal_546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_361 ( .s (reset), .b ({signal_3371, signal_1582}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_3503, signal_548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_364 ( .s (reset), .b ({signal_3372, signal_1581}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_3505, signal_550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_367 ( .s (reset), .b ({signal_3373, signal_1580}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_3507, signal_552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_370 ( .s (reset), .b ({signal_3374, signal_1579}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_3509, signal_554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_373 ( .s (reset), .b ({signal_3375, signal_1578}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_3511, signal_556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_376 ( .s (reset), .b ({signal_3376, signal_1577}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_3513, signal_558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_379 ( .s (reset), .b ({signal_3377, signal_1576}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_3515, signal_560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_382 ( .s (reset), .b ({signal_3378, signal_1575}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_3517, signal_562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_385 ( .s (reset), .b ({signal_3379, signal_1574}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_3519, signal_564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_388 ( .s (reset), .b ({signal_3380, signal_1573}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_3521, signal_566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_391 ( .s (reset), .b ({signal_3381, signal_1572}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_3523, signal_568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_394 ( .s (reset), .b ({signal_3382, signal_1571}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_3525, signal_570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_397 ( .s (reset), .b ({signal_3383, signal_1570}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_3527, signal_572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_400 ( .s (reset), .b ({signal_3384, signal_1569}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_3529, signal_574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_403 ( .s (reset), .b ({signal_3385, signal_1568}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_3531, signal_576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_406 ( .s (reset), .b ({signal_3386, signal_1567}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_3533, signal_578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_409 ( .s (reset), .b ({signal_3387, signal_1566}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_3535, signal_580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_412 ( .s (reset), .b ({signal_3388, signal_1565}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_3537, signal_582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_415 ( .s (reset), .b ({signal_3389, signal_1564}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_3539, signal_584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_418 ( .s (reset), .b ({signal_3390, signal_1563}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_3541, signal_586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_421 ( .s (reset), .b ({signal_3391, signal_1562}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_3543, signal_588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_424 ( .s (reset), .b ({signal_3392, signal_1561}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_3545, signal_590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_427 ( .s (reset), .b ({signal_3393, signal_1560}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_3547, signal_592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_430 ( .s (reset), .b ({signal_3394, signal_1559}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_3549, signal_594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_433 ( .s (reset), .b ({signal_3395, signal_1558}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_3551, signal_596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_436 ( .s (reset), .b ({signal_3396, signal_1557}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_3553, signal_598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_439 ( .s (reset), .b ({signal_3397, signal_1556}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_3555, signal_600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_442 ( .s (reset), .b ({signal_3398, signal_1555}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_3557, signal_602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_445 ( .s (reset), .b ({signal_3399, signal_1554}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_3559, signal_604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_448 ( .s (reset), .b ({signal_3400, signal_1553}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_3561, signal_606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_451 ( .s (reset), .b ({signal_3401, signal_1552}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_3563, signal_608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_454 ( .s (reset), .b ({signal_3402, signal_1551}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_3565, signal_610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_457 ( .s (reset), .b ({signal_3403, signal_1550}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_3567, signal_612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_460 ( .s (reset), .b ({signal_3404, signal_1549}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_3569, signal_614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_463 ( .s (reset), .b ({signal_3405, signal_1548}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_3571, signal_616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_466 ( .s (reset), .b ({signal_3406, signal_1547}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_3573, signal_618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_469 ( .s (reset), .b ({signal_3407, signal_1546}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_3575, signal_620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_472 ( .s (reset), .b ({signal_3408, signal_1545}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_3577, signal_622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_475 ( .s (reset), .b ({signal_3409, signal_1544}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_3579, signal_624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_478 ( .s (reset), .b ({signal_3410, signal_1543}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_3581, signal_626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_481 ( .s (reset), .b ({signal_3411, signal_1542}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_3583, signal_628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_484 ( .s (reset), .b ({signal_3412, signal_1541}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_3585, signal_630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_487 ( .s (reset), .b ({signal_3413, signal_1540}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_3587, signal_632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_490 ( .s (reset), .b ({signal_3414, signal_1539}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_3589, signal_634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_493 ( .s (reset), .b ({signal_3415, signal_1538}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_3591, signal_636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_496 ( .s (reset), .b ({signal_3416, signal_1537}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_3593, signal_638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_499 ( .s (reset), .b ({signal_3417, signal_1536}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_3595, signal_640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_502 ( .s (reset), .b ({signal_3418, signal_1535}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_3597, signal_642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_505 ( .s (reset), .b ({signal_3419, signal_1534}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_3599, signal_644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_508 ( .s (reset), .b ({signal_3420, signal_1533}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_3601, signal_646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_511 ( .s (reset), .b ({signal_3421, signal_1532}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_3603, signal_648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_514 ( .s (reset), .b ({signal_3422, signal_1531}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_3605, signal_650}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_517 ( .s (reset), .b ({signal_3423, signal_1530}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_3607, signal_652}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_520 ( .s (reset), .b ({signal_3424, signal_1529}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_3609, signal_654}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_523 ( .s (reset), .b ({signal_3425, signal_1528}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_3611, signal_656}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_526 ( .s (reset), .b ({signal_3426, signal_1527}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_3613, signal_658}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_529 ( .s (reset), .b ({signal_3427, signal_1526}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_3615, signal_660}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_532 ( .s (reset), .b ({signal_3428, signal_1525}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_3617, signal_662}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_535 ( .s (reset), .b ({signal_3429, signal_1524}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_3619, signal_664}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_538 ( .s (reset), .b ({signal_3430, signal_1523}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_3621, signal_666}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_541 ( .s (reset), .b ({signal_3431, signal_1522}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_3623, signal_668}) ) ;
    INV_X1 cell_542 ( .A (signal_393), .ZN (signal_670) ) ;
    INV_X1 cell_543 ( .A (signal_670), .ZN (signal_672) ) ;
    INV_X1 cell_544 ( .A (signal_670), .ZN (signal_671) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_545 ( .s (signal_671), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({signal_3026, signal_1809}), .c ({signal_3305, signal_1841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_546 ( .s (signal_671), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({signal_3029, signal_1808}), .c ({signal_3306, signal_1840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_547 ( .s (signal_671), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({signal_3032, signal_1807}), .c ({signal_3307, signal_1839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_548 ( .s (signal_671), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({signal_3035, signal_1806}), .c ({signal_3308, signal_1838}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_549 ( .s (signal_671), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({signal_3041, signal_1805}), .c ({signal_3309, signal_1837}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_550 ( .s (signal_671), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({signal_3044, signal_1804}), .c ({signal_3310, signal_1836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_551 ( .s (signal_671), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({signal_3047, signal_1803}), .c ({signal_3311, signal_1835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_552 ( .s (signal_671), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({signal_3050, signal_1802}), .c ({signal_3312, signal_1834}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_553 ( .s (signal_393), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({signal_3269, signal_1801}), .c ({signal_3304, signal_1833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_554 ( .s (signal_672), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({signal_3302, signal_1800}), .c ({signal_3313, signal_1832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_555 ( .s (signal_672), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({signal_2954, signal_1799}), .c ({signal_3314, signal_1831}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_556 ( .s (signal_672), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({signal_2987, signal_1798}), .c ({signal_3315, signal_1830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_557 ( .s (signal_672), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({signal_3014, signal_1797}), .c ({signal_3316, signal_1829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_558 ( .s (signal_671), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({signal_3017, signal_1796}), .c ({signal_3317, signal_1828}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_559 ( .s (signal_671), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({signal_3020, signal_1795}), .c ({signal_3318, signal_1827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_560 ( .s (signal_672), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({signal_3023, signal_1794}), .c ({signal_3319, signal_1826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_561 ( .s (signal_671), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({signal_2921, signal_1793}), .c ({signal_3320, signal_1825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_562 ( .s (signal_672), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({signal_3038, signal_1792}), .c ({signal_3321, signal_1824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_563 ( .s (signal_672), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({signal_3071, signal_1791}), .c ({signal_3322, signal_1823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_564 ( .s (signal_672), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({signal_3104, signal_1790}), .c ({signal_3323, signal_1822}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_565 ( .s (signal_672), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({signal_3137, signal_1789}), .c ({signal_3324, signal_1821}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_566 ( .s (signal_672), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({signal_3170, signal_1788}), .c ({signal_3325, signal_1820}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_567 ( .s (signal_672), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({signal_3203, signal_1787}), .c ({signal_3326, signal_1819}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_568 ( .s (signal_672), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({signal_3236, signal_1786}), .c ({signal_3327, signal_1818}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_569 ( .s (signal_672), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({signal_3053, signal_1785}), .c ({signal_3328, signal_1817}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_570 ( .s (signal_672), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({signal_3056, signal_1784}), .c ({signal_3329, signal_1816}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_571 ( .s (signal_672), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({signal_3059, signal_1783}), .c ({signal_3330, signal_1815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_572 ( .s (signal_672), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({signal_3062, signal_1782}), .c ({signal_3331, signal_1814}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_573 ( .s (signal_672), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({signal_3065, signal_1781}), .c ({signal_3332, signal_1813}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_574 ( .s (signal_672), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({signal_3068, signal_1780}), .c ({signal_3333, signal_1812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_575 ( .s (signal_672), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({signal_3074, signal_1779}), .c ({signal_3334, signal_1811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_576 ( .s (signal_672), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({signal_3077, signal_1778}), .c ({signal_3335, signal_1810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_581 ( .a ({signal_3308, signal_1838}), .b ({signal_3306, signal_1840}), .c ({signal_3624, signal_788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_709 ( .a ({signal_3315, signal_1830}), .b ({signal_3313, signal_1832}), .c ({signal_3625, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_837 ( .a ({signal_3323, signal_1822}), .b ({signal_3321, signal_1824}), .c ({signal_3626, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_965 ( .a ({signal_3331, signal_1814}), .b ({signal_3329, signal_1816}), .c ({signal_3627, signal_1148}) ) ;
    INV_X1 cell_1197 ( .A (signal_394), .ZN (signal_1217) ) ;
    INV_X1 cell_1198 ( .A (signal_1217), .ZN (signal_1218) ) ;
    INV_X1 cell_1199 ( .A (signal_1217), .ZN (signal_1219) ) ;
    INV_X1 cell_1232 ( .A (signal_393), .ZN (signal_1220) ) ;
    INV_X1 cell_1233 ( .A (signal_1220), .ZN (signal_1223) ) ;
    INV_X1 cell_1234 ( .A (signal_1220), .ZN (signal_1225) ) ;
    INV_X1 cell_1235 ( .A (signal_1220), .ZN (signal_1226) ) ;
    INV_X1 cell_1236 ( .A (signal_1220), .ZN (signal_1224) ) ;
    INV_X1 cell_1237 ( .A (signal_1220), .ZN (signal_1221) ) ;
    INV_X1 cell_1238 ( .A (signal_1220), .ZN (signal_1222) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1271 ( .s (signal_1221), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({signal_3186, signal_1745}), .c ({signal_3336, signal_1617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1272 ( .s (signal_1222), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({signal_3189, signal_1744}), .c ({signal_3337, signal_1616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1273 ( .s (signal_1226), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({signal_3192, signal_1743}), .c ({signal_3338, signal_1615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1274 ( .s (signal_1225), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({signal_3195, signal_1742}), .c ({signal_3339, signal_1614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1275 ( .s (signal_1224), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({signal_3198, signal_1741}), .c ({signal_3340, signal_1613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1276 ( .s (signal_1223), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({signal_3201, signal_1740}), .c ({signal_3341, signal_1612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1277 ( .s (signal_1222), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({signal_3207, signal_1739}), .c ({signal_3342, signal_1611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1278 ( .s (signal_1221), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({signal_3210, signal_1738}), .c ({signal_3343, signal_1610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1279 ( .s (signal_1221), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({signal_2937, signal_1737}), .c ({signal_3344, signal_1609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1280 ( .s (signal_1226), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({signal_2940, signal_1736}), .c ({signal_3345, signal_1608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1281 ( .s (signal_1225), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({signal_2943, signal_1735}), .c ({signal_3346, signal_1607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1282 ( .s (signal_1224), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({signal_2946, signal_1734}), .c ({signal_3347, signal_1606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1283 ( .s (signal_1226), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({signal_2949, signal_1733}), .c ({signal_3348, signal_1605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1284 ( .s (signal_1225), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({signal_2952, signal_1732}), .c ({signal_3349, signal_1604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1285 ( .s (signal_1224), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({signal_2958, signal_1731}), .c ({signal_3350, signal_1603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1286 ( .s (signal_1223), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({signal_2961, signal_1730}), .c ({signal_3351, signal_1602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1287 ( .s (signal_1222), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({signal_3027, signal_1729}), .c ({signal_3352, signal_1601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1288 ( .s (signal_1221), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({signal_3030, signal_1728}), .c ({signal_3353, signal_1600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1289 ( .s (signal_1226), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({signal_3033, signal_1727}), .c ({signal_3354, signal_1599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1290 ( .s (signal_1225), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({signal_3036, signal_1726}), .c ({signal_3355, signal_1598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1291 ( .s (signal_1224), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({signal_3042, signal_1725}), .c ({signal_3356, signal_1597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1292 ( .s (signal_1223), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({signal_3045, signal_1724}), .c ({signal_3357, signal_1596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1293 ( .s (signal_1222), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({signal_3048, signal_1723}), .c ({signal_3358, signal_1595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1294 ( .s (signal_1221), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({signal_3051, signal_1722}), .c ({signal_3359, signal_1594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1295 ( .s (signal_1221), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_3159, signal_1721}), .c ({signal_3360, signal_1593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1296 ( .s (signal_1221), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_3162, signal_1720}), .c ({signal_3361, signal_1592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1297 ( .s (signal_1221), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_3165, signal_1719}), .c ({signal_3362, signal_1591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1298 ( .s (signal_1221), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_3168, signal_1718}), .c ({signal_3363, signal_1590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1299 ( .s (signal_1221), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_3174, signal_1717}), .c ({signal_3364, signal_1589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1300 ( .s (signal_1221), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_3177, signal_1716}), .c ({signal_3365, signal_1588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1301 ( .s (signal_1221), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_3180, signal_1715}), .c ({signal_3366, signal_1587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1302 ( .s (signal_1221), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_3183, signal_1714}), .c ({signal_3367, signal_1586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1303 ( .s (signal_1221), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({signal_3291, signal_1713}), .c ({signal_3368, signal_1585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1304 ( .s (signal_1221), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({signal_3294, signal_1712}), .c ({signal_3369, signal_1584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1305 ( .s (signal_1221), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({signal_3297, signal_1711}), .c ({signal_3370, signal_1583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1306 ( .s (signal_1221), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({signal_3300, signal_1710}), .c ({signal_3371, signal_1582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1307 ( .s (signal_1222), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({signal_2925, signal_1709}), .c ({signal_3372, signal_1581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1308 ( .s (signal_1222), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({signal_2928, signal_1708}), .c ({signal_3373, signal_1580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1309 ( .s (signal_1222), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({signal_2931, signal_1707}), .c ({signal_3374, signal_1579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1310 ( .s (signal_1222), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({signal_2934, signal_1706}), .c ({signal_3375, signal_1578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1311 ( .s (signal_1222), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({signal_3270, signal_1705}), .c ({signal_3376, signal_1577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1312 ( .s (signal_1222), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({signal_3303, signal_1704}), .c ({signal_3377, signal_1576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1313 ( .s (signal_1222), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({signal_2955, signal_1703}), .c ({signal_3378, signal_1575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1314 ( .s (signal_1222), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({signal_2988, signal_1702}), .c ({signal_3379, signal_1574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1315 ( .s (signal_1222), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({signal_3015, signal_1701}), .c ({signal_3380, signal_1573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1316 ( .s (signal_1222), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({signal_3018, signal_1700}), .c ({signal_3381, signal_1572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1317 ( .s (signal_1222), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({signal_3021, signal_1699}), .c ({signal_3382, signal_1571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1318 ( .s (signal_1222), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({signal_3024, signal_1698}), .c ({signal_3383, signal_1570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1319 ( .s (signal_1223), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({signal_3132, signal_1697}), .c ({signal_3384, signal_1569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1320 ( .s (signal_1223), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({signal_3135, signal_1696}), .c ({signal_3385, signal_1568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1321 ( .s (signal_1223), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({signal_3141, signal_1695}), .c ({signal_3386, signal_1567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1322 ( .s (signal_1223), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({signal_3144, signal_1694}), .c ({signal_3387, signal_1566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1323 ( .s (signal_1223), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({signal_3147, signal_1693}), .c ({signal_3388, signal_1565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1324 ( .s (signal_1223), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({signal_3150, signal_1692}), .c ({signal_3389, signal_1564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1325 ( .s (signal_1223), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({signal_3153, signal_1691}), .c ({signal_3390, signal_1563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1326 ( .s (signal_1223), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({signal_3156, signal_1690}), .c ({signal_3391, signal_1562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1327 ( .s (signal_1223), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_3264, signal_1689}), .c ({signal_3392, signal_1561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1328 ( .s (signal_1223), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_3267, signal_1688}), .c ({signal_3393, signal_1560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1329 ( .s (signal_1223), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_3273, signal_1687}), .c ({signal_3394, signal_1559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1330 ( .s (signal_1223), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_3276, signal_1686}), .c ({signal_3395, signal_1558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1331 ( .s (signal_1224), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_3279, signal_1685}), .c ({signal_3396, signal_1557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1332 ( .s (signal_1224), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_3282, signal_1684}), .c ({signal_3397, signal_1556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1333 ( .s (signal_1224), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_3285, signal_1683}), .c ({signal_3398, signal_1555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1334 ( .s (signal_1224), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_3288, signal_1682}), .c ({signal_3399, signal_1554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1335 ( .s (signal_1224), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({signal_2922, signal_1681}), .c ({signal_3400, signal_1553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1336 ( .s (signal_1224), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({signal_3039, signal_1680}), .c ({signal_3401, signal_1552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1337 ( .s (signal_1224), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({signal_3072, signal_1679}), .c ({signal_3402, signal_1551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1338 ( .s (signal_1224), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({signal_3105, signal_1678}), .c ({signal_3403, signal_1550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1339 ( .s (signal_1224), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({signal_3138, signal_1677}), .c ({signal_3404, signal_1549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1340 ( .s (signal_1224), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({signal_3171, signal_1676}), .c ({signal_3405, signal_1548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1341 ( .s (signal_1224), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({signal_3204, signal_1675}), .c ({signal_3406, signal_1547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1342 ( .s (signal_1224), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({signal_3237, signal_1674}), .c ({signal_3407, signal_1546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1343 ( .s (signal_1225), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({signal_3108, signal_1673}), .c ({signal_3408, signal_1545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1344 ( .s (signal_1225), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({signal_3111, signal_1672}), .c ({signal_3409, signal_1544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1345 ( .s (signal_1225), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({signal_3114, signal_1671}), .c ({signal_3410, signal_1543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1346 ( .s (signal_1225), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({signal_3117, signal_1670}), .c ({signal_3411, signal_1542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1347 ( .s (signal_1225), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({signal_3120, signal_1669}), .c ({signal_3412, signal_1541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1348 ( .s (signal_1225), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({signal_3123, signal_1668}), .c ({signal_3413, signal_1540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1349 ( .s (signal_1225), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({signal_3126, signal_1667}), .c ({signal_3414, signal_1539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1350 ( .s (signal_1225), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({signal_3129, signal_1666}), .c ({signal_3415, signal_1538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1351 ( .s (signal_1225), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({signal_3240, signal_1665}), .c ({signal_3416, signal_1537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1352 ( .s (signal_1225), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({signal_3243, signal_1664}), .c ({signal_3417, signal_1536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1353 ( .s (signal_1225), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({signal_3246, signal_1663}), .c ({signal_3418, signal_1535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1354 ( .s (signal_1225), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({signal_3249, signal_1662}), .c ({signal_3419, signal_1534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1355 ( .s (signal_1226), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({signal_3252, signal_1661}), .c ({signal_3420, signal_1533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1356 ( .s (signal_1226), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({signal_3255, signal_1660}), .c ({signal_3421, signal_1532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1357 ( .s (signal_1226), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({signal_3258, signal_1659}), .c ({signal_3422, signal_1531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1358 ( .s (signal_1226), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({signal_3261, signal_1658}), .c ({signal_3423, signal_1530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1359 ( .s (signal_1226), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_2991, signal_1657}), .c ({signal_3424, signal_1529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1360 ( .s (signal_1226), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_2994, signal_1656}), .c ({signal_3425, signal_1528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1361 ( .s (signal_1226), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_2997, signal_1655}), .c ({signal_3426, signal_1527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1362 ( .s (signal_1226), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_3000, signal_1654}), .c ({signal_3427, signal_1526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1363 ( .s (signal_1226), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_3003, signal_1653}), .c ({signal_3428, signal_1525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1364 ( .s (signal_1226), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_3006, signal_1652}), .c ({signal_3429, signal_1524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1365 ( .s (signal_1226), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_3009, signal_1651}), .c ({signal_3430, signal_1523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1366 ( .s (signal_1226), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_3012, signal_1650}), .c ({signal_3431, signal_1522}) ) ;
    INV_X1 cell_1887 ( .A (signal_1483), .ZN (signal_1490) ) ;
    INV_X1 cell_1888 ( .A (signal_393), .ZN (signal_1483) ) ;
    INV_X1 cell_1889 ( .A (signal_1483), .ZN (signal_1488) ) ;
    INV_X1 cell_1890 ( .A (signal_1483), .ZN (signal_1487) ) ;
    INV_X1 cell_1891 ( .A (signal_1483), .ZN (signal_1486) ) ;
    INV_X1 cell_1892 ( .A (signal_1483), .ZN (signal_1485) ) ;
    INV_X1 cell_1893 ( .A (signal_1483), .ZN (signal_1484) ) ;
    INV_X1 cell_1894 ( .A (signal_1483), .ZN (signal_1489) ) ;
    NOR2_X1 cell_2023 ( .A1 (reset), .A2 (signal_1491), .ZN (signal_1502) ) ;
    XNOR2_X1 cell_2024 ( .A (signal_2273), .B (signal_393), .ZN (signal_1491) ) ;
    NOR2_X1 cell_2025 ( .A1 (reset), .A2 (signal_1492), .ZN (signal_1501) ) ;
    XOR2_X1 cell_2026 ( .A (signal_2272), .B (signal_1493), .Z (signal_1492) ) ;
    NOR2_X1 cell_2027 ( .A1 (reset), .A2 (signal_1494), .ZN (signal_1498) ) ;
    XOR2_X1 cell_2028 ( .A (signal_2270), .B (signal_1495), .Z (signal_1494) ) ;
    NAND2_X1 cell_2029 ( .A1 (signal_1496), .A2 (signal_2271), .ZN (signal_1495) ) ;
    NOR2_X1 cell_2030 ( .A1 (reset), .A2 (signal_1497), .ZN (signal_1499) ) ;
    XNOR2_X1 cell_2031 ( .A (signal_2271), .B (signal_1496), .ZN (signal_1497) ) ;
    NOR2_X1 cell_2032 ( .A1 (signal_1500), .A2 (signal_1493), .ZN (signal_1496) ) ;
    NAND2_X1 cell_2033 ( .A1 (signal_393), .A2 (signal_2273), .ZN (signal_1493) ) ;
    INV_X1 cell_2036 ( .A (signal_2272), .ZN (signal_1500) ) ;
    NOR2_X1 cell_2042 ( .A1 (reset), .A2 (signal_1506), .ZN (signal_1520) ) ;
    XOR2_X1 cell_2043 ( .A (signal_2276), .B (signal_1507), .Z (signal_1506) ) ;
    NAND2_X1 cell_2044 ( .A1 (signal_1508), .A2 (1'b1), .ZN (signal_1507) ) ;
    NAND2_X1 cell_2045 ( .A1 (signal_1509), .A2 (signal_2274), .ZN (signal_1508) ) ;
    NAND2_X1 cell_2046 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_1509) ) ;
    NOR2_X1 cell_2047 ( .A1 (reset), .A2 (signal_1510), .ZN (signal_1519) ) ;
    MUX2_X1 cell_2048 ( .S (signal_2275), .A (signal_1511), .B (signal_1512), .Z (signal_1510) ) ;
    NOR2_X1 cell_2049 ( .A1 (reset), .A2 (signal_1513), .ZN (signal_1518) ) ;
    NOR2_X1 cell_2050 ( .A1 (signal_1514), .A2 (signal_1515), .ZN (signal_1513) ) ;
    NOR2_X1 cell_2051 ( .A1 (signal_1516), .A2 (signal_1511), .ZN (signal_1515) ) ;
    NAND2_X1 cell_2052 ( .A1 (signal_1512), .A2 (signal_1517), .ZN (signal_1511) ) ;
    AND2_X1 cell_2053 ( .A1 (signal_2276), .A2 (1'b1), .ZN (signal_1512) ) ;
    NOR2_X1 cell_2054 ( .A1 (1'b1), .A2 (signal_1517), .ZN (signal_1514) ) ;
    INV_X1 cell_2057 ( .A (signal_2275), .ZN (signal_1516) ) ;
    INV_X1 cell_2059 ( .A (signal_2274), .ZN (signal_1517) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2061 ( .a ({signal_3309, signal_1837}), .b ({signal_3312, signal_1834}), .c ({signal_3628, signal_2338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2062 ( .a ({signal_3307, signal_1839}), .b ({signal_3312, signal_1834}), .c ({signal_3629, signal_2339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2063 ( .a ({signal_3306, signal_1840}), .b ({signal_3312, signal_1834}), .c ({signal_3630, signal_2340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2064 ( .a ({signal_3307, signal_1839}), .b ({signal_3309, signal_1837}), .c ({signal_3631, signal_2341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2065 ( .a ({signal_3310, signal_1836}), .b ({signal_3311, signal_1835}), .c ({signal_3632, signal_2342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2066 ( .a ({signal_3307, signal_1839}), .b ({signal_3311, signal_1835}), .c ({signal_3633, signal_2343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2067 ( .a ({signal_3307, signal_1839}), .b ({signal_3310, signal_1836}), .c ({signal_3634, signal_2344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2068 ( .a ({signal_3305, signal_1841}), .b ({signal_3309, signal_1837}), .c ({signal_3635, signal_2345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2069 ( .a ({signal_3305, signal_1841}), .b ({signal_3306, signal_1840}), .c ({signal_3636, signal_2346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2070 ( .a ({signal_3316, signal_1829}), .b ({signal_3319, signal_1826}), .c ({signal_3637, signal_2347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2071 ( .a ({signal_3314, signal_1831}), .b ({signal_3319, signal_1826}), .c ({signal_3638, signal_2348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2072 ( .a ({signal_3313, signal_1832}), .b ({signal_3319, signal_1826}), .c ({signal_3639, signal_2349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2073 ( .a ({signal_3314, signal_1831}), .b ({signal_3316, signal_1829}), .c ({signal_3640, signal_2350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2074 ( .a ({signal_3317, signal_1828}), .b ({signal_3318, signal_1827}), .c ({signal_3641, signal_2351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2075 ( .a ({signal_3314, signal_1831}), .b ({signal_3318, signal_1827}), .c ({signal_3642, signal_2352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2076 ( .a ({signal_3314, signal_1831}), .b ({signal_3317, signal_1828}), .c ({signal_3643, signal_2353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2077 ( .a ({signal_3304, signal_1833}), .b ({signal_3316, signal_1829}), .c ({signal_3644, signal_2354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2078 ( .a ({signal_3304, signal_1833}), .b ({signal_3313, signal_1832}), .c ({signal_3645, signal_2355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2079 ( .a ({signal_3324, signal_1821}), .b ({signal_3327, signal_1818}), .c ({signal_3646, signal_2356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2080 ( .a ({signal_3322, signal_1823}), .b ({signal_3327, signal_1818}), .c ({signal_3647, signal_2357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2081 ( .a ({signal_3321, signal_1824}), .b ({signal_3327, signal_1818}), .c ({signal_3648, signal_2358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2082 ( .a ({signal_3322, signal_1823}), .b ({signal_3324, signal_1821}), .c ({signal_3649, signal_2359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2083 ( .a ({signal_3325, signal_1820}), .b ({signal_3326, signal_1819}), .c ({signal_3650, signal_2360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2084 ( .a ({signal_3322, signal_1823}), .b ({signal_3326, signal_1819}), .c ({signal_3651, signal_2361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2085 ( .a ({signal_3322, signal_1823}), .b ({signal_3325, signal_1820}), .c ({signal_3652, signal_2362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2086 ( .a ({signal_3320, signal_1825}), .b ({signal_3324, signal_1821}), .c ({signal_3653, signal_2363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2087 ( .a ({signal_3320, signal_1825}), .b ({signal_3321, signal_1824}), .c ({signal_3654, signal_2364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2088 ( .a ({signal_3332, signal_1813}), .b ({signal_3335, signal_1810}), .c ({signal_3655, signal_2365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2089 ( .a ({signal_3330, signal_1815}), .b ({signal_3335, signal_1810}), .c ({signal_3656, signal_2366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2090 ( .a ({signal_3329, signal_1816}), .b ({signal_3335, signal_1810}), .c ({signal_3657, signal_2367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2091 ( .a ({signal_3330, signal_1815}), .b ({signal_3332, signal_1813}), .c ({signal_3658, signal_2368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2092 ( .a ({signal_3333, signal_1812}), .b ({signal_3334, signal_1811}), .c ({signal_3659, signal_2369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2093 ( .a ({signal_3330, signal_1815}), .b ({signal_3334, signal_1811}), .c ({signal_3660, signal_2370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2094 ( .a ({signal_3330, signal_1815}), .b ({signal_3333, signal_1812}), .c ({signal_3661, signal_2371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2095 ( .a ({signal_3328, signal_1817}), .b ({signal_3332, signal_1813}), .c ({signal_3662, signal_2372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2096 ( .a ({signal_3328, signal_1817}), .b ({signal_3329, signal_1816}), .c ({signal_3663, signal_2373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2097 ( .a ({signal_3624, signal_788}), .b ({signal_3628, signal_2338}), .c ({signal_3664, signal_2374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2098 ( .a ({signal_3305, signal_1841}), .b ({signal_3632, signal_2342}), .c ({signal_3665, signal_2375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2099 ( .a ({signal_3630, signal_2340}), .b ({signal_3631, signal_2341}), .c ({signal_3666, signal_2376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2100 ( .a ({signal_3624, signal_788}), .b ({signal_3633, signal_2343}), .c ({signal_3667, signal_2377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2101 ( .a ({signal_3624, signal_788}), .b ({signal_3634, signal_2344}), .c ({signal_3668, signal_2378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2102 ( .a ({signal_3632, signal_2342}), .b ({signal_3635, signal_2345}), .c ({signal_3669, signal_2379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2103 ( .a ({signal_3632, signal_2342}), .b ({signal_3636, signal_2346}), .c ({signal_3670, signal_2380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2104 ( .a ({signal_3628, signal_2338}), .b ({signal_3634, signal_2344}), .c ({signal_3671, signal_2381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2105 ( .a ({signal_3625, signal_908}), .b ({signal_3637, signal_2347}), .c ({signal_3672, signal_2382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2106 ( .a ({signal_3304, signal_1833}), .b ({signal_3641, signal_2351}), .c ({signal_3673, signal_2383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2107 ( .a ({signal_3639, signal_2349}), .b ({signal_3640, signal_2350}), .c ({signal_3674, signal_2384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2108 ( .a ({signal_3625, signal_908}), .b ({signal_3642, signal_2352}), .c ({signal_3675, signal_2385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2109 ( .a ({signal_3625, signal_908}), .b ({signal_3643, signal_2353}), .c ({signal_3676, signal_2386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2110 ( .a ({signal_3641, signal_2351}), .b ({signal_3644, signal_2354}), .c ({signal_3677, signal_2387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2111 ( .a ({signal_3641, signal_2351}), .b ({signal_3645, signal_2355}), .c ({signal_3678, signal_2388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2112 ( .a ({signal_3637, signal_2347}), .b ({signal_3643, signal_2353}), .c ({signal_3679, signal_2389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2113 ( .a ({signal_3626, signal_1028}), .b ({signal_3646, signal_2356}), .c ({signal_3680, signal_2390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2114 ( .a ({signal_3320, signal_1825}), .b ({signal_3650, signal_2360}), .c ({signal_3681, signal_2391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2115 ( .a ({signal_3648, signal_2358}), .b ({signal_3649, signal_2359}), .c ({signal_3682, signal_2392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2116 ( .a ({signal_3626, signal_1028}), .b ({signal_3651, signal_2361}), .c ({signal_3683, signal_2393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2117 ( .a ({signal_3626, signal_1028}), .b ({signal_3652, signal_2362}), .c ({signal_3684, signal_2394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2118 ( .a ({signal_3650, signal_2360}), .b ({signal_3653, signal_2363}), .c ({signal_3685, signal_2395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2119 ( .a ({signal_3650, signal_2360}), .b ({signal_3654, signal_2364}), .c ({signal_3686, signal_2396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2120 ( .a ({signal_3646, signal_2356}), .b ({signal_3652, signal_2362}), .c ({signal_3687, signal_2397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2121 ( .a ({signal_3627, signal_1148}), .b ({signal_3655, signal_2365}), .c ({signal_3688, signal_2398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2122 ( .a ({signal_3328, signal_1817}), .b ({signal_3659, signal_2369}), .c ({signal_3689, signal_2399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2123 ( .a ({signal_3657, signal_2367}), .b ({signal_3658, signal_2368}), .c ({signal_3690, signal_2400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2124 ( .a ({signal_3627, signal_1148}), .b ({signal_3660, signal_2370}), .c ({signal_3691, signal_2401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2125 ( .a ({signal_3627, signal_1148}), .b ({signal_3661, signal_2371}), .c ({signal_3692, signal_2402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2126 ( .a ({signal_3659, signal_2369}), .b ({signal_3662, signal_2372}), .c ({signal_3693, signal_2403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2127 ( .a ({signal_3659, signal_2369}), .b ({signal_3663, signal_2373}), .c ({signal_3694, signal_2404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2128 ( .a ({signal_3655, signal_2365}), .b ({signal_3661, signal_2371}), .c ({signal_3695, signal_2405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2153 ( .a ({signal_3305, signal_1841}), .b ({signal_3664, signal_2374}), .c ({signal_3720, signal_2430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2154 ( .a ({signal_3632, signal_2342}), .b ({signal_3664, signal_2374}), .c ({signal_3721, signal_2431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2155 ( .a ({signal_3633, signal_2343}), .b ({signal_3664, signal_2374}), .c ({signal_3722, signal_2432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2156 ( .a ({signal_3665, signal_2375}), .b ({signal_3668, signal_2378}), .c ({signal_3723, signal_2433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2157 ( .a ({signal_3628, signal_2338}), .b ({signal_3669, signal_2379}), .c ({signal_3724, signal_2434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2158 ( .a ({signal_3629, signal_2339}), .b ({signal_3670, signal_2380}), .c ({signal_3725, signal_2435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2159 ( .a ({signal_3630, signal_2340}), .b ({signal_3668, signal_2378}), .c ({signal_3726, signal_2436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2160 ( .a ({signal_3304, signal_1833}), .b ({signal_3672, signal_2382}), .c ({signal_3727, signal_2437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2161 ( .a ({signal_3641, signal_2351}), .b ({signal_3672, signal_2382}), .c ({signal_3728, signal_2438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2162 ( .a ({signal_3642, signal_2352}), .b ({signal_3672, signal_2382}), .c ({signal_3729, signal_2439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2163 ( .a ({signal_3673, signal_2383}), .b ({signal_3676, signal_2386}), .c ({signal_3730, signal_2440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2164 ( .a ({signal_3637, signal_2347}), .b ({signal_3677, signal_2387}), .c ({signal_3731, signal_2441}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2165 ( .a ({signal_3638, signal_2348}), .b ({signal_3678, signal_2388}), .c ({signal_3732, signal_2442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2166 ( .a ({signal_3639, signal_2349}), .b ({signal_3676, signal_2386}), .c ({signal_3733, signal_2443}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2167 ( .a ({signal_3320, signal_1825}), .b ({signal_3680, signal_2390}), .c ({signal_3734, signal_2444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2168 ( .a ({signal_3650, signal_2360}), .b ({signal_3680, signal_2390}), .c ({signal_3735, signal_2445}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2169 ( .a ({signal_3651, signal_2361}), .b ({signal_3680, signal_2390}), .c ({signal_3736, signal_2446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2170 ( .a ({signal_3681, signal_2391}), .b ({signal_3684, signal_2394}), .c ({signal_3737, signal_2447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2171 ( .a ({signal_3646, signal_2356}), .b ({signal_3685, signal_2395}), .c ({signal_3738, signal_2448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2172 ( .a ({signal_3647, signal_2357}), .b ({signal_3686, signal_2396}), .c ({signal_3739, signal_2449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2173 ( .a ({signal_3648, signal_2358}), .b ({signal_3684, signal_2394}), .c ({signal_3740, signal_2450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2174 ( .a ({signal_3328, signal_1817}), .b ({signal_3688, signal_2398}), .c ({signal_3741, signal_2451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2175 ( .a ({signal_3659, signal_2369}), .b ({signal_3688, signal_2398}), .c ({signal_3742, signal_2452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2176 ( .a ({signal_3660, signal_2370}), .b ({signal_3688, signal_2398}), .c ({signal_3743, signal_2453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2177 ( .a ({signal_3689, signal_2399}), .b ({signal_3692, signal_2402}), .c ({signal_3744, signal_2454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2178 ( .a ({signal_3655, signal_2365}), .b ({signal_3693, signal_2403}), .c ({signal_3745, signal_2455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2179 ( .a ({signal_3656, signal_2366}), .b ({signal_3694, signal_2404}), .c ({signal_3746, signal_2456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2180 ( .a ({signal_3657, signal_2367}), .b ({signal_3692, signal_2402}), .c ({signal_3747, signal_2457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2193 ( .a ({signal_3629, signal_2339}), .b ({signal_3721, signal_2431}), .c ({signal_3760, signal_2470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2194 ( .a ({signal_3723, signal_2433}), .b ({signal_3724, signal_2434}), .c ({signal_3761, signal_2471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2199 ( .a ({signal_3638, signal_2348}), .b ({signal_3728, signal_2438}), .c ({signal_3766, signal_2476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2200 ( .a ({signal_3730, signal_2440}), .b ({signal_3731, signal_2441}), .c ({signal_3767, signal_2477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2205 ( .a ({signal_3647, signal_2357}), .b ({signal_3735, signal_2445}), .c ({signal_3772, signal_2482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2206 ( .a ({signal_3737, signal_2447}), .b ({signal_3738, signal_2448}), .c ({signal_3773, signal_2483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2211 ( .a ({signal_3656, signal_2366}), .b ({signal_3742, signal_2452}), .c ({signal_3778, signal_2488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2212 ( .a ({signal_3744, signal_2454}), .b ({signal_3745, signal_2455}), .c ({signal_3779, signal_2489}) ) ;
    ClockGatingController #(9) cell_2707 ( .clk (clk), .rst (reset), .GatedClk (signal_5060), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2129 ( .a ({signal_3664, signal_2374}), .b ({signal_3666, signal_2376}), .clk (clk), .r (Fresh[0]), .c ({signal_3696, signal_2406}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2130 ( .a ({signal_3305, signal_1841}), .b ({signal_3669, signal_2379}), .clk (clk), .r (Fresh[1]), .c ({signal_3697, signal_2407}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2131 ( .a ({signal_3630, signal_2340}), .b ({signal_3668, signal_2378}), .clk (clk), .r (Fresh[2]), .c ({signal_3698, signal_2408}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2132 ( .a ({signal_3665, signal_2375}), .b ({signal_3670, signal_2380}), .clk (clk), .r (Fresh[3]), .c ({signal_3699, signal_2409}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2133 ( .a ({signal_3628, signal_2338}), .b ({signal_3667, signal_2377}), .clk (clk), .r (Fresh[4]), .c ({signal_3700, signal_2410}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2134 ( .a ({signal_3631, signal_2341}), .b ({signal_3671, signal_2381}), .clk (clk), .r (Fresh[5]), .c ({signal_3701, signal_2411}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2135 ( .a ({signal_3672, signal_2382}), .b ({signal_3674, signal_2384}), .clk (clk), .r (Fresh[6]), .c ({signal_3702, signal_2412}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2136 ( .a ({signal_3304, signal_1833}), .b ({signal_3677, signal_2387}), .clk (clk), .r (Fresh[7]), .c ({signal_3703, signal_2413}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2137 ( .a ({signal_3639, signal_2349}), .b ({signal_3676, signal_2386}), .clk (clk), .r (Fresh[8]), .c ({signal_3704, signal_2414}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2138 ( .a ({signal_3673, signal_2383}), .b ({signal_3678, signal_2388}), .clk (clk), .r (Fresh[9]), .c ({signal_3705, signal_2415}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2139 ( .a ({signal_3637, signal_2347}), .b ({signal_3675, signal_2385}), .clk (clk), .r (Fresh[10]), .c ({signal_3706, signal_2416}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2140 ( .a ({signal_3640, signal_2350}), .b ({signal_3679, signal_2389}), .clk (clk), .r (Fresh[11]), .c ({signal_3707, signal_2417}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2141 ( .a ({signal_3680, signal_2390}), .b ({signal_3682, signal_2392}), .clk (clk), .r (Fresh[12]), .c ({signal_3708, signal_2418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2142 ( .a ({signal_3320, signal_1825}), .b ({signal_3685, signal_2395}), .clk (clk), .r (Fresh[13]), .c ({signal_3709, signal_2419}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2143 ( .a ({signal_3648, signal_2358}), .b ({signal_3684, signal_2394}), .clk (clk), .r (Fresh[14]), .c ({signal_3710, signal_2420}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2144 ( .a ({signal_3681, signal_2391}), .b ({signal_3686, signal_2396}), .clk (clk), .r (Fresh[15]), .c ({signal_3711, signal_2421}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2145 ( .a ({signal_3646, signal_2356}), .b ({signal_3683, signal_2393}), .clk (clk), .r (Fresh[16]), .c ({signal_3712, signal_2422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2146 ( .a ({signal_3649, signal_2359}), .b ({signal_3687, signal_2397}), .clk (clk), .r (Fresh[17]), .c ({signal_3713, signal_2423}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2147 ( .a ({signal_3688, signal_2398}), .b ({signal_3690, signal_2400}), .clk (clk), .r (Fresh[18]), .c ({signal_3714, signal_2424}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2148 ( .a ({signal_3328, signal_1817}), .b ({signal_3693, signal_2403}), .clk (clk), .r (Fresh[19]), .c ({signal_3715, signal_2425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2149 ( .a ({signal_3657, signal_2367}), .b ({signal_3692, signal_2402}), .clk (clk), .r (Fresh[20]), .c ({signal_3716, signal_2426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2150 ( .a ({signal_3689, signal_2399}), .b ({signal_3694, signal_2404}), .clk (clk), .r (Fresh[21]), .c ({signal_3717, signal_2427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2151 ( .a ({signal_3655, signal_2365}), .b ({signal_3691, signal_2401}), .clk (clk), .r (Fresh[22]), .c ({signal_3718, signal_2428}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2152 ( .a ({signal_3658, signal_2368}), .b ({signal_3695, signal_2405}), .clk (clk), .r (Fresh[23]), .c ({signal_3719, signal_2429}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2181 ( .a ({signal_3720, signal_2430}), .b ({signal_3725, signal_2435}), .clk (clk), .r (Fresh[24]), .c ({signal_3748, signal_2458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2182 ( .a ({signal_3723, signal_2433}), .b ({signal_3724, signal_2434}), .clk (clk), .r (Fresh[25]), .c ({signal_3749, signal_2459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2183 ( .a ({signal_3629, signal_2339}), .b ({signal_3721, signal_2431}), .clk (clk), .r (Fresh[26]), .c ({signal_3750, signal_2460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2184 ( .a ({signal_3727, signal_2437}), .b ({signal_3732, signal_2442}), .clk (clk), .r (Fresh[27]), .c ({signal_3751, signal_2461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2185 ( .a ({signal_3730, signal_2440}), .b ({signal_3731, signal_2441}), .clk (clk), .r (Fresh[28]), .c ({signal_3752, signal_2462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2186 ( .a ({signal_3638, signal_2348}), .b ({signal_3728, signal_2438}), .clk (clk), .r (Fresh[29]), .c ({signal_3753, signal_2463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2187 ( .a ({signal_3734, signal_2444}), .b ({signal_3739, signal_2449}), .clk (clk), .r (Fresh[30]), .c ({signal_3754, signal_2464}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2188 ( .a ({signal_3737, signal_2447}), .b ({signal_3738, signal_2448}), .clk (clk), .r (Fresh[31]), .c ({signal_3755, signal_2465}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2189 ( .a ({signal_3647, signal_2357}), .b ({signal_3735, signal_2445}), .clk (clk), .r (Fresh[32]), .c ({signal_3756, signal_2466}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2190 ( .a ({signal_3741, signal_2451}), .b ({signal_3746, signal_2456}), .clk (clk), .r (Fresh[33]), .c ({signal_3757, signal_2467}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2191 ( .a ({signal_3744, signal_2454}), .b ({signal_3745, signal_2455}), .clk (clk), .r (Fresh[34]), .c ({signal_3758, signal_2468}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2192 ( .a ({signal_3656, signal_2366}), .b ({signal_3742, signal_2452}), .clk (clk), .r (Fresh[35]), .c ({signal_3759, signal_2469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2195 ( .a ({signal_3722, signal_2432}), .b ({signal_3696, signal_2406}), .c ({signal_3762, signal_2472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2196 ( .a ({signal_3696, signal_2406}), .b ({signal_3697, signal_2407}), .c ({signal_3763, signal_2473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2197 ( .a ({signal_3726, signal_2436}), .b ({signal_3698, signal_2408}), .c ({signal_3764, signal_2474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2198 ( .a ({signal_3700, signal_2410}), .b ({signal_3701, signal_2411}), .c ({signal_3765, signal_2475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2201 ( .a ({signal_3729, signal_2439}), .b ({signal_3702, signal_2412}), .c ({signal_3768, signal_2478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2202 ( .a ({signal_3702, signal_2412}), .b ({signal_3703, signal_2413}), .c ({signal_3769, signal_2479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2203 ( .a ({signal_3733, signal_2443}), .b ({signal_3704, signal_2414}), .c ({signal_3770, signal_2480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2204 ( .a ({signal_3706, signal_2416}), .b ({signal_3707, signal_2417}), .c ({signal_3771, signal_2481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2207 ( .a ({signal_3736, signal_2446}), .b ({signal_3708, signal_2418}), .c ({signal_3774, signal_2484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2208 ( .a ({signal_3708, signal_2418}), .b ({signal_3709, signal_2419}), .c ({signal_3775, signal_2485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2209 ( .a ({signal_3740, signal_2450}), .b ({signal_3710, signal_2420}), .c ({signal_3776, signal_2486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2210 ( .a ({signal_3712, signal_2422}), .b ({signal_3713, signal_2423}), .c ({signal_3777, signal_2487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2213 ( .a ({signal_3743, signal_2453}), .b ({signal_3714, signal_2424}), .c ({signal_3780, signal_2490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2214 ( .a ({signal_3714, signal_2424}), .b ({signal_3715, signal_2425}), .c ({signal_3781, signal_2491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2215 ( .a ({signal_3747, signal_2457}), .b ({signal_3716, signal_2426}), .c ({signal_3782, signal_2492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2216 ( .a ({signal_3718, signal_2428}), .b ({signal_3719, signal_2429}), .c ({signal_3783, signal_2493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2217 ( .a ({signal_3698, signal_2408}), .b ({signal_3749, signal_2459}), .c ({signal_3784, signal_2494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2218 ( .a ({signal_3700, signal_2410}), .b ({signal_3750, signal_2460}), .c ({signal_3785, signal_2495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2219 ( .a ({signal_3748, signal_2458}), .b ({signal_3762, signal_2472}), .c ({signal_3786, signal_2496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2220 ( .a ({signal_3760, signal_2470}), .b ({signal_3763, signal_2473}), .c ({signal_3787, signal_2497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2221 ( .a ({signal_3699, signal_2409}), .b ({signal_3764, signal_2474}), .c ({signal_3788, signal_2498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2222 ( .a ({signal_3704, signal_2414}), .b ({signal_3752, signal_2462}), .c ({signal_3789, signal_2499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2223 ( .a ({signal_3706, signal_2416}), .b ({signal_3753, signal_2463}), .c ({signal_3790, signal_2500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2224 ( .a ({signal_3751, signal_2461}), .b ({signal_3768, signal_2478}), .c ({signal_3791, signal_2501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2225 ( .a ({signal_3766, signal_2476}), .b ({signal_3769, signal_2479}), .c ({signal_3792, signal_2502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2226 ( .a ({signal_3705, signal_2415}), .b ({signal_3770, signal_2480}), .c ({signal_3793, signal_2503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2227 ( .a ({signal_3710, signal_2420}), .b ({signal_3755, signal_2465}), .c ({signal_3794, signal_2504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2228 ( .a ({signal_3712, signal_2422}), .b ({signal_3756, signal_2466}), .c ({signal_3795, signal_2505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2229 ( .a ({signal_3754, signal_2464}), .b ({signal_3774, signal_2484}), .c ({signal_3796, signal_2506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2230 ( .a ({signal_3772, signal_2482}), .b ({signal_3775, signal_2485}), .c ({signal_3797, signal_2507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2231 ( .a ({signal_3711, signal_2421}), .b ({signal_3776, signal_2486}), .c ({signal_3798, signal_2508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2232 ( .a ({signal_3716, signal_2426}), .b ({signal_3758, signal_2468}), .c ({signal_3799, signal_2509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2233 ( .a ({signal_3718, signal_2428}), .b ({signal_3759, signal_2469}), .c ({signal_3800, signal_2510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2234 ( .a ({signal_3757, signal_2467}), .b ({signal_3780, signal_2490}), .c ({signal_3801, signal_2511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2235 ( .a ({signal_3778, signal_2488}), .b ({signal_3781, signal_2491}), .c ({signal_3802, signal_2512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2236 ( .a ({signal_3717, signal_2427}), .b ({signal_3782, signal_2492}), .c ({signal_3803, signal_2513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2237 ( .a ({signal_3784, signal_2494}), .b ({signal_3785, signal_2495}), .c ({signal_3804, signal_2514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2238 ( .a ({signal_3765, signal_2475}), .b ({signal_3786, signal_2496}), .c ({signal_3805, signal_2515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2239 ( .a ({signal_3785, signal_2495}), .b ({signal_3787, signal_2497}), .c ({signal_3806, signal_2516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2240 ( .a ({signal_3765, signal_2475}), .b ({signal_3788, signal_2498}), .c ({signal_3807, signal_2517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2241 ( .a ({signal_3789, signal_2499}), .b ({signal_3790, signal_2500}), .c ({signal_3808, signal_2518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2242 ( .a ({signal_3771, signal_2481}), .b ({signal_3791, signal_2501}), .c ({signal_3809, signal_2519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2243 ( .a ({signal_3790, signal_2500}), .b ({signal_3792, signal_2502}), .c ({signal_3810, signal_2520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2244 ( .a ({signal_3771, signal_2481}), .b ({signal_3793, signal_2503}), .c ({signal_3811, signal_2521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2245 ( .a ({signal_3794, signal_2504}), .b ({signal_3795, signal_2505}), .c ({signal_3812, signal_2522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2246 ( .a ({signal_3777, signal_2487}), .b ({signal_3796, signal_2506}), .c ({signal_3813, signal_2523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2247 ( .a ({signal_3795, signal_2505}), .b ({signal_3797, signal_2507}), .c ({signal_3814, signal_2524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2248 ( .a ({signal_3777, signal_2487}), .b ({signal_3798, signal_2508}), .c ({signal_3815, signal_2525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2249 ( .a ({signal_3799, signal_2509}), .b ({signal_3800, signal_2510}), .c ({signal_3816, signal_2526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2250 ( .a ({signal_3783, signal_2493}), .b ({signal_3801, signal_2511}), .c ({signal_3817, signal_2527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2251 ( .a ({signal_3800, signal_2510}), .b ({signal_3802, signal_2512}), .c ({signal_3818, signal_2528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2252 ( .a ({signal_3783, signal_2493}), .b ({signal_3803, signal_2513}), .c ({signal_3819, signal_2529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2261 ( .a ({signal_3761, signal_2471}), .b ({signal_3804, signal_2514}), .c ({signal_3828, signal_2538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2262 ( .a ({signal_3805, signal_2515}), .b ({signal_3806, signal_2516}), .c ({signal_3829, signal_2539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2263 ( .a ({signal_3767, signal_2477}), .b ({signal_3808, signal_2518}), .c ({signal_3830, signal_2540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2264 ( .a ({signal_3809, signal_2519}), .b ({signal_3810, signal_2520}), .c ({signal_3831, signal_2541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2265 ( .a ({signal_3773, signal_2483}), .b ({signal_3812, signal_2522}), .c ({signal_3832, signal_2542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2266 ( .a ({signal_3813, signal_2523}), .b ({signal_3814, signal_2524}), .c ({signal_3833, signal_2543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2267 ( .a ({signal_3779, signal_2489}), .b ({signal_3816, signal_2526}), .c ({signal_3834, signal_2544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2268 ( .a ({signal_3817, signal_2527}), .b ({signal_3818, signal_2528}), .c ({signal_3835, signal_2545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2273 ( .a ({signal_3807, signal_2517}), .b ({signal_3828, signal_2538}), .c ({signal_3840, signal_2550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2277 ( .a ({signal_3811, signal_2521}), .b ({signal_3830, signal_2540}), .c ({signal_3844, signal_2554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2281 ( .a ({signal_3815, signal_2525}), .b ({signal_3832, signal_2542}), .c ({signal_3848, signal_2558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2285 ( .a ({signal_3819, signal_2529}), .b ({signal_3834, signal_2544}), .c ({signal_3852, signal_2562}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2253 ( .a ({signal_3805, signal_2515}), .b ({signal_3807, signal_2517}), .clk (clk), .r (Fresh[36]), .c ({signal_3820, signal_2530}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2254 ( .a ({signal_3806, signal_2516}), .b ({signal_3807, signal_2517}), .clk (clk), .r (Fresh[37]), .c ({signal_3821, signal_2531}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2255 ( .a ({signal_3809, signal_2519}), .b ({signal_3811, signal_2521}), .clk (clk), .r (Fresh[38]), .c ({signal_3822, signal_2532}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2256 ( .a ({signal_3810, signal_2520}), .b ({signal_3811, signal_2521}), .clk (clk), .r (Fresh[39]), .c ({signal_3823, signal_2533}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2257 ( .a ({signal_3813, signal_2523}), .b ({signal_3815, signal_2525}), .clk (clk), .r (Fresh[40]), .c ({signal_3824, signal_2534}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2258 ( .a ({signal_3814, signal_2524}), .b ({signal_3815, signal_2525}), .clk (clk), .r (Fresh[41]), .c ({signal_3825, signal_2535}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2259 ( .a ({signal_3817, signal_2527}), .b ({signal_3819, signal_2529}), .clk (clk), .r (Fresh[42]), .c ({signal_3826, signal_2536}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2260 ( .a ({signal_3818, signal_2528}), .b ({signal_3819, signal_2529}), .clk (clk), .r (Fresh[43]), .c ({signal_3827, signal_2537}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2269 ( .a ({signal_3805, signal_2515}), .b ({signal_3828, signal_2538}), .clk (clk), .r (Fresh[44]), .c ({signal_3836, signal_2546}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2270 ( .a ({signal_3809, signal_2519}), .b ({signal_3830, signal_2540}), .clk (clk), .r (Fresh[45]), .c ({signal_3837, signal_2547}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2271 ( .a ({signal_3813, signal_2523}), .b ({signal_3832, signal_2542}), .clk (clk), .r (Fresh[46]), .c ({signal_3838, signal_2548}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2272 ( .a ({signal_3817, signal_2527}), .b ({signal_3834, signal_2544}), .clk (clk), .r (Fresh[47]), .c ({signal_3839, signal_2549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2274 ( .a ({signal_3806, signal_2516}), .b ({signal_3820, signal_2530}), .c ({signal_3841, signal_2551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2275 ( .a ({signal_3828, signal_2538}), .b ({signal_3820, signal_2530}), .c ({signal_3842, signal_2552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2276 ( .a ({signal_3820, signal_2530}), .b ({signal_3829, signal_2539}), .c ({signal_3843, signal_2553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2278 ( .a ({signal_3810, signal_2520}), .b ({signal_3822, signal_2532}), .c ({signal_3845, signal_2555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2279 ( .a ({signal_3830, signal_2540}), .b ({signal_3822, signal_2532}), .c ({signal_3846, signal_2556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2280 ( .a ({signal_3822, signal_2532}), .b ({signal_3831, signal_2541}), .c ({signal_3847, signal_2557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2282 ( .a ({signal_3814, signal_2524}), .b ({signal_3824, signal_2534}), .c ({signal_3849, signal_2559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2283 ( .a ({signal_3832, signal_2542}), .b ({signal_3824, signal_2534}), .c ({signal_3850, signal_2560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2284 ( .a ({signal_3824, signal_2534}), .b ({signal_3833, signal_2543}), .c ({signal_3851, signal_2561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2286 ( .a ({signal_3818, signal_2528}), .b ({signal_3826, signal_2536}), .c ({signal_3853, signal_2563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2287 ( .a ({signal_3834, signal_2544}), .b ({signal_3826, signal_2536}), .c ({signal_3854, signal_2564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2288 ( .a ({signal_3826, signal_2536}), .b ({signal_3835, signal_2545}), .c ({signal_3855, signal_2565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2305 ( .a ({signal_3820, signal_2530}), .b ({signal_3840, signal_2550}), .c ({signal_3872, signal_2582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2306 ( .a ({signal_3822, signal_2532}), .b ({signal_3844, signal_2554}), .c ({signal_3873, signal_2583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2307 ( .a ({signal_3824, signal_2534}), .b ({signal_3848, signal_2558}), .c ({signal_3874, signal_2584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2308 ( .a ({signal_3826, signal_2536}), .b ({signal_3852, signal_2562}), .c ({signal_3875, signal_2585}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2289 ( .a ({signal_3829, signal_2539}), .b ({signal_3842, signal_2552}), .clk (clk), .r (Fresh[48]), .c ({signal_3856, signal_2566}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2290 ( .a ({signal_3840, signal_2550}), .b ({signal_3841, signal_2551}), .clk (clk), .r (Fresh[49]), .c ({signal_3857, signal_2567}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2291 ( .a ({signal_3829, signal_2539}), .b ({signal_3836, signal_2546}), .clk (clk), .r (Fresh[50]), .c ({signal_3858, signal_2568}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2292 ( .a ({signal_3821, signal_2531}), .b ({signal_3840, signal_2550}), .clk (clk), .r (Fresh[51]), .c ({signal_3859, signal_2569}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2293 ( .a ({signal_3831, signal_2541}), .b ({signal_3846, signal_2556}), .clk (clk), .r (Fresh[52]), .c ({signal_3860, signal_2570}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2294 ( .a ({signal_3844, signal_2554}), .b ({signal_3845, signal_2555}), .clk (clk), .r (Fresh[53]), .c ({signal_3861, signal_2571}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2295 ( .a ({signal_3831, signal_2541}), .b ({signal_3837, signal_2547}), .clk (clk), .r (Fresh[54]), .c ({signal_3862, signal_2572}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2296 ( .a ({signal_3823, signal_2533}), .b ({signal_3844, signal_2554}), .clk (clk), .r (Fresh[55]), .c ({signal_3863, signal_2573}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2297 ( .a ({signal_3833, signal_2543}), .b ({signal_3850, signal_2560}), .clk (clk), .r (Fresh[56]), .c ({signal_3864, signal_2574}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2298 ( .a ({signal_3848, signal_2558}), .b ({signal_3849, signal_2559}), .clk (clk), .r (Fresh[57]), .c ({signal_3865, signal_2575}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2299 ( .a ({signal_3833, signal_2543}), .b ({signal_3838, signal_2548}), .clk (clk), .r (Fresh[58]), .c ({signal_3866, signal_2576}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2300 ( .a ({signal_3825, signal_2535}), .b ({signal_3848, signal_2558}), .clk (clk), .r (Fresh[59]), .c ({signal_3867, signal_2577}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2301 ( .a ({signal_3835, signal_2545}), .b ({signal_3854, signal_2564}), .clk (clk), .r (Fresh[60]), .c ({signal_3868, signal_2578}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2302 ( .a ({signal_3852, signal_2562}), .b ({signal_3853, signal_2563}), .clk (clk), .r (Fresh[61]), .c ({signal_3869, signal_2579}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2303 ( .a ({signal_3835, signal_2545}), .b ({signal_3839, signal_2549}), .clk (clk), .r (Fresh[62]), .c ({signal_3870, signal_2580}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2304 ( .a ({signal_3827, signal_2537}), .b ({signal_3852, signal_2562}), .clk (clk), .r (Fresh[63]), .c ({signal_3871, signal_2581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2309 ( .a ({signal_3806, signal_2516}), .b ({signal_3856, signal_2566}), .c ({signal_3876, signal_2586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2310 ( .a ({signal_3843, signal_2553}), .b ({signal_3858, signal_2568}), .c ({signal_3877, signal_2587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2311 ( .a ({signal_3828, signal_2538}), .b ({signal_3857, signal_2567}), .c ({signal_3878, signal_2588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2312 ( .a ({signal_3859, signal_2569}), .b ({signal_3872, signal_2582}), .c ({signal_3879, signal_2589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2313 ( .a ({signal_3810, signal_2520}), .b ({signal_3860, signal_2570}), .c ({signal_3880, signal_2590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2314 ( .a ({signal_3847, signal_2557}), .b ({signal_3862, signal_2572}), .c ({signal_3881, signal_2591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2315 ( .a ({signal_3830, signal_2540}), .b ({signal_3861, signal_2571}), .c ({signal_3882, signal_2592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2316 ( .a ({signal_3863, signal_2573}), .b ({signal_3873, signal_2583}), .c ({signal_3883, signal_2593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2317 ( .a ({signal_3814, signal_2524}), .b ({signal_3864, signal_2574}), .c ({signal_3884, signal_2594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2318 ( .a ({signal_3851, signal_2561}), .b ({signal_3866, signal_2576}), .c ({signal_3885, signal_2595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2319 ( .a ({signal_3832, signal_2542}), .b ({signal_3865, signal_2575}), .c ({signal_3886, signal_2596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2320 ( .a ({signal_3867, signal_2577}), .b ({signal_3874, signal_2584}), .c ({signal_3887, signal_2597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2321 ( .a ({signal_3818, signal_2528}), .b ({signal_3868, signal_2578}), .c ({signal_3888, signal_2598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2322 ( .a ({signal_3855, signal_2565}), .b ({signal_3870, signal_2580}), .c ({signal_3889, signal_2599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2323 ( .a ({signal_3834, signal_2544}), .b ({signal_3869, signal_2579}), .c ({signal_3890, signal_2600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2324 ( .a ({signal_3871, signal_2581}), .b ({signal_3875, signal_2585}), .c ({signal_3891, signal_2601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2357 ( .a ({signal_3877, signal_2587}), .b ({signal_3879, signal_2589}), .c ({signal_3924, signal_2634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2358 ( .a ({signal_3876, signal_2586}), .b ({signal_3878, signal_2588}), .c ({signal_3925, signal_2635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2359 ( .a ({signal_3876, signal_2586}), .b ({signal_3877, signal_2587}), .c ({signal_3926, signal_2636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2360 ( .a ({signal_3878, signal_2588}), .b ({signal_3879, signal_2589}), .c ({signal_3927, signal_2637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2361 ( .a ({signal_3881, signal_2591}), .b ({signal_3883, signal_2593}), .c ({signal_3928, signal_2638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2362 ( .a ({signal_3880, signal_2590}), .b ({signal_3882, signal_2592}), .c ({signal_3929, signal_2639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2363 ( .a ({signal_3880, signal_2590}), .b ({signal_3881, signal_2591}), .c ({signal_3930, signal_2640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2364 ( .a ({signal_3882, signal_2592}), .b ({signal_3883, signal_2593}), .c ({signal_3931, signal_2641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2365 ( .a ({signal_3885, signal_2595}), .b ({signal_3887, signal_2597}), .c ({signal_3932, signal_2642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2366 ( .a ({signal_3884, signal_2594}), .b ({signal_3886, signal_2596}), .c ({signal_3933, signal_2643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2367 ( .a ({signal_3884, signal_2594}), .b ({signal_3885, signal_2595}), .c ({signal_3934, signal_2644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2368 ( .a ({signal_3886, signal_2596}), .b ({signal_3887, signal_2597}), .c ({signal_3935, signal_2645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2369 ( .a ({signal_3889, signal_2599}), .b ({signal_3891, signal_2601}), .c ({signal_3936, signal_2646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2370 ( .a ({signal_3888, signal_2598}), .b ({signal_3890, signal_2600}), .c ({signal_3937, signal_2647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2371 ( .a ({signal_3888, signal_2598}), .b ({signal_3889, signal_2599}), .c ({signal_3938, signal_2648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2372 ( .a ({signal_3890, signal_2600}), .b ({signal_3891, signal_2601}), .c ({signal_3939, signal_2649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2405 ( .a ({signal_3924, signal_2634}), .b ({signal_3925, signal_2635}), .c ({signal_3972, signal_2682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2409 ( .a ({signal_3928, signal_2638}), .b ({signal_3929, signal_2639}), .c ({signal_3976, signal_2686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2413 ( .a ({signal_3932, signal_2642}), .b ({signal_3933, signal_2643}), .c ({signal_3980, signal_2690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2417 ( .a ({signal_3936, signal_2646}), .b ({signal_3937, signal_2647}), .c ({signal_3984, signal_2694}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_160 ( .s (reset), .b ({signal_4725, signal_1649}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_4830, signal_414}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_163 ( .s (reset), .b ({signal_4869, signal_1648}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_4911, signal_416}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_166 ( .s (reset), .b ({signal_4581, signal_1647}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_4706, signal_418}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_169 ( .s (reset), .b ({signal_4726, signal_1646}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_4832, signal_420}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_172 ( .s (reset), .b ({signal_4727, signal_1645}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_4834, signal_422}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_175 ( .s (reset), .b ({signal_4728, signal_1644}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_4836, signal_424}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_178 ( .s (reset), .b ({signal_4729, signal_1643}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_4838, signal_426}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_181 ( .s (reset), .b ({signal_4582, signal_1642}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_4708, signal_428}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_184 ( .s (reset), .b ({signal_4730, signal_1641}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_4840, signal_430}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_187 ( .s (reset), .b ({signal_4870, signal_1640}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_4913, signal_432}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_190 ( .s (reset), .b ({signal_4583, signal_1639}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_4710, signal_434}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_193 ( .s (reset), .b ({signal_4731, signal_1638}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_4842, signal_436}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_196 ( .s (reset), .b ({signal_4732, signal_1637}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_4844, signal_438}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_199 ( .s (reset), .b ({signal_4733, signal_1636}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_4846, signal_440}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_202 ( .s (reset), .b ({signal_4734, signal_1635}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_4848, signal_442}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_205 ( .s (reset), .b ({signal_4584, signal_1634}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_4712, signal_444}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_208 ( .s (reset), .b ({signal_4735, signal_1633}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_4850, signal_446}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_211 ( .s (reset), .b ({signal_4871, signal_1632}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_4915, signal_448}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_214 ( .s (reset), .b ({signal_4585, signal_1631}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_4714, signal_450}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_217 ( .s (reset), .b ({signal_4736, signal_1630}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_4852, signal_452}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_220 ( .s (reset), .b ({signal_4737, signal_1629}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_4854, signal_454}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_223 ( .s (reset), .b ({signal_4738, signal_1628}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_4856, signal_456}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_226 ( .s (reset), .b ({signal_4739, signal_1627}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_4858, signal_458}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_229 ( .s (reset), .b ({signal_4586, signal_1626}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_4716, signal_460}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_232 ( .s (reset), .b ({signal_4740, signal_1625}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_4860, signal_462}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_235 ( .s (reset), .b ({signal_4872, signal_1624}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_4917, signal_464}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_238 ( .s (reset), .b ({signal_4587, signal_1623}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_4718, signal_466}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_241 ( .s (reset), .b ({signal_4741, signal_1622}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_4862, signal_468}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_244 ( .s (reset), .b ({signal_4742, signal_1621}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_4864, signal_470}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_247 ( .s (reset), .b ({signal_4743, signal_1620}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_4866, signal_472}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_250 ( .s (reset), .b ({signal_4744, signal_1619}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_4868, signal_474}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_253 ( .s (reset), .b ({signal_4588, signal_1618}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_4720, signal_476}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .a ({signal_4537, signal_1153}), .b ({signal_4168, signal_2328}), .c ({signal_4560, signal_1868}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_4374, signal_1216}), .b ({signal_4109, signal_2321}), .c ({signal_4406, signal_1877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1200 ( .s (signal_1218), .b ({signal_4406, signal_1877}), .a ({signal_4108, signal_1845}), .c ({signal_4561, signal_1909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1201 ( .s (signal_394), .b ({signal_4703, signal_1876}), .a ({signal_4162, signal_2303}), .c ({signal_4721, signal_1908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1202 ( .s (signal_394), .b ({signal_4384, signal_1875}), .a ({signal_4117, signal_1843}), .c ({signal_4407, signal_1907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1203 ( .s (signal_394), .b ({signal_4550, signal_1874}), .a ({signal_4116, signal_1842}), .c ({signal_4562, signal_1906}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1204 ( .s (signal_394), .b ({signal_4549, signal_1873}), .a ({signal_4115, signal_2300}), .c ({signal_4563, signal_1905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1205 ( .s (signal_394), .b ({signal_4540, signal_1872}), .a ({signal_4161, signal_2299}), .c ({signal_4564, signal_1904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1206 ( .s (signal_394), .b ({signal_4539, signal_1871}), .a ({signal_4160, signal_2298}), .c ({signal_4565, signal_1903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1207 ( .s (signal_1219), .b ({signal_4377, signal_1870}), .a ({signal_4112, signal_2305}), .c ({signal_4408, signal_1902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1208 ( .s (signal_1218), .b ({signal_4538, signal_1869}), .a ({signal_4109, signal_2321}), .c ({signal_4566, signal_1901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1209 ( .s (signal_1218), .b ({signal_4560, signal_1868}), .a ({signal_4165, signal_2320}), .c ({signal_4722, signal_1900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1210 ( .s (signal_1218), .b ({signal_4405, signal_1867}), .a ({signal_4124, signal_2319}), .c ({signal_4409, signal_1899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1211 ( .s (signal_1218), .b ({signal_4559, signal_1866}), .a ({signal_4123, signal_2318}), .c ({signal_4567, signal_1898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1212 ( .s (signal_1218), .b ({signal_4558, signal_1865}), .a ({signal_4122, signal_2317}), .c ({signal_4568, signal_1897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1213 ( .s (signal_1218), .b ({signal_4548, signal_1864}), .a ({signal_4164, signal_2316}), .c ({signal_4569, signal_1896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1214 ( .s (signal_1218), .b ({signal_4547, signal_1863}), .a ({signal_4163, signal_2315}), .c ({signal_4570, signal_1895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1215 ( .s (signal_1218), .b ({signal_4400, signal_1862}), .a ({signal_4119, signal_2314}), .c ({signal_4410, signal_1894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1216 ( .s (signal_1218), .b ({signal_4546, signal_1861}), .a ({signal_4110, signal_2329}), .c ({signal_4571, signal_1893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1217 ( .s (signal_1218), .b ({signal_4704, signal_1860}), .a ({signal_4168, signal_2328}), .c ({signal_4723, signal_1892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1218 ( .s (signal_1218), .b ({signal_4397, signal_1859}), .a ({signal_4131, signal_2327}), .c ({signal_4411, signal_1891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1219 ( .s (signal_1218), .b ({signal_4556, signal_1858}), .a ({signal_4130, signal_2326}), .c ({signal_4572, signal_1890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1220 ( .s (signal_1219), .b ({signal_4554, signal_1857}), .a ({signal_4129, signal_2325}), .c ({signal_4573, signal_1889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1221 ( .s (signal_1219), .b ({signal_4545, signal_1856}), .a ({signal_4167, signal_2324}), .c ({signal_4574, signal_1888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1222 ( .s (signal_1219), .b ({signal_4544, signal_1855}), .a ({signal_4166, signal_2323}), .c ({signal_4575, signal_1887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1223 ( .s (signal_1219), .b ({signal_4391, signal_1854}), .a ({signal_4126, signal_2322}), .c ({signal_4412, signal_1886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1224 ( .s (signal_1219), .b ({signal_4543, signal_1853}), .a ({signal_4111, signal_2337}), .c ({signal_4576, signal_1885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1225 ( .s (signal_1219), .b ({signal_4702, signal_1852}), .a ({signal_4171, signal_2336}), .c ({signal_4724, signal_1884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1226 ( .s (signal_1219), .b ({signal_4388, signal_1851}), .a ({signal_4138, signal_2335}), .c ({signal_4413, signal_1883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1227 ( .s (signal_1219), .b ({signal_4552, signal_1850}), .a ({signal_4137, signal_2334}), .c ({signal_4577, signal_1882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1228 ( .s (signal_1219), .b ({signal_4551, signal_1849}), .a ({signal_4136, signal_2333}), .c ({signal_4578, signal_1881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1229 ( .s (signal_1219), .b ({signal_4542, signal_1848}), .a ({signal_4170, signal_2332}), .c ({signal_4579, signal_1880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1230 ( .s (signal_1219), .b ({signal_4541, signal_1847}), .a ({signal_4169, signal_2331}), .c ({signal_4580, signal_1879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1231 ( .s (signal_1219), .b ({signal_4382, signal_1846}), .a ({signal_4133, signal_2330}), .c ({signal_4414, signal_1878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1239 ( .s (signal_393), .b ({signal_4561, signal_1909}), .a ({signal_3081, signal_1777}), .c ({signal_4725, signal_1649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1240 ( .s (signal_1226), .b ({signal_4721, signal_1908}), .a ({signal_3084, signal_1776}), .c ({signal_4869, signal_1648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1241 ( .s (signal_1225), .b ({signal_4407, signal_1907}), .a ({signal_3087, signal_1775}), .c ({signal_4581, signal_1647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1242 ( .s (signal_1224), .b ({signal_4562, signal_1906}), .a ({signal_3090, signal_1774}), .c ({signal_4726, signal_1646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1243 ( .s (signal_1223), .b ({signal_4563, signal_1905}), .a ({signal_3093, signal_1773}), .c ({signal_4727, signal_1645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1244 ( .s (signal_1222), .b ({signal_4564, signal_1904}), .a ({signal_3096, signal_1772}), .c ({signal_4728, signal_1644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1245 ( .s (signal_1221), .b ({signal_4565, signal_1903}), .a ({signal_3099, signal_1771}), .c ({signal_4729, signal_1643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1246 ( .s (signal_1226), .b ({signal_4408, signal_1902}), .a ({signal_3102, signal_1770}), .c ({signal_4582, signal_1642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1247 ( .s (signal_1223), .b ({signal_4566, signal_1901}), .a ({signal_3213, signal_1769}), .c ({signal_4730, signal_1641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1248 ( .s (signal_1226), .b ({signal_4722, signal_1900}), .a ({signal_3216, signal_1768}), .c ({signal_4870, signal_1640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1249 ( .s (signal_393), .b ({signal_4409, signal_1899}), .a ({signal_3219, signal_1767}), .c ({signal_4583, signal_1639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1250 ( .s (signal_393), .b ({signal_4567, signal_1898}), .a ({signal_3222, signal_1766}), .c ({signal_4731, signal_1638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1251 ( .s (signal_393), .b ({signal_4568, signal_1897}), .a ({signal_3225, signal_1765}), .c ({signal_4732, signal_1637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1252 ( .s (signal_393), .b ({signal_4569, signal_1896}), .a ({signal_3228, signal_1764}), .c ({signal_4733, signal_1636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1253 ( .s (signal_393), .b ({signal_4570, signal_1895}), .a ({signal_3231, signal_1763}), .c ({signal_4734, signal_1635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1254 ( .s (signal_393), .b ({signal_4410, signal_1894}), .a ({signal_3234, signal_1762}), .c ({signal_4584, signal_1634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1255 ( .s (signal_393), .b ({signal_4571, signal_1893}), .a ({signal_2964, signal_1761}), .c ({signal_4735, signal_1633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1256 ( .s (signal_393), .b ({signal_4723, signal_1892}), .a ({signal_2967, signal_1760}), .c ({signal_4871, signal_1632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1257 ( .s (signal_393), .b ({signal_4411, signal_1891}), .a ({signal_2970, signal_1759}), .c ({signal_4585, signal_1631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1258 ( .s (signal_393), .b ({signal_4572, signal_1890}), .a ({signal_2973, signal_1758}), .c ({signal_4736, signal_1630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1259 ( .s (signal_1225), .b ({signal_4573, signal_1889}), .a ({signal_2976, signal_1757}), .c ({signal_4737, signal_1629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1260 ( .s (signal_1224), .b ({signal_4574, signal_1888}), .a ({signal_2979, signal_1756}), .c ({signal_4738, signal_1628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1261 ( .s (signal_1223), .b ({signal_4575, signal_1887}), .a ({signal_2982, signal_1755}), .c ({signal_4739, signal_1627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1262 ( .s (signal_1222), .b ({signal_4412, signal_1886}), .a ({signal_2985, signal_1754}), .c ({signal_4586, signal_1626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1263 ( .s (signal_1221), .b ({signal_4576, signal_1885}), .a ({signal_3054, signal_1753}), .c ({signal_4740, signal_1625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1264 ( .s (signal_1223), .b ({signal_4724, signal_1884}), .a ({signal_3057, signal_1752}), .c ({signal_4872, signal_1624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1265 ( .s (signal_1222), .b ({signal_4413, signal_1883}), .a ({signal_3060, signal_1751}), .c ({signal_4587, signal_1623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1266 ( .s (signal_393), .b ({signal_4577, signal_1882}), .a ({signal_3063, signal_1750}), .c ({signal_4741, signal_1622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1267 ( .s (signal_393), .b ({signal_4578, signal_1881}), .a ({signal_3066, signal_1749}), .c ({signal_4742, signal_1621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1268 ( .s (signal_1226), .b ({signal_4579, signal_1880}), .a ({signal_3069, signal_1748}), .c ({signal_4743, signal_1620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1269 ( .s (signal_1225), .b ({signal_4580, signal_1879}), .a ({signal_3075, signal_1747}), .c ({signal_4744, signal_1619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1270 ( .s (signal_1224), .b ({signal_4414, signal_1878}), .a ({signal_3078, signal_1746}), .c ({signal_4588, signal_1618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1369 ( .s (reset), .b ({signal_4670, signal_2037}), .a ({key_s1[0], key_s0[0]}), .c ({signal_4746, signal_1227}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1372 ( .s (reset), .b ({signal_4812, signal_2036}), .a ({key_s1[1], key_s0[1]}), .c ({signal_4874, signal_1229}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1375 ( .s (reset), .b ({signal_4671, signal_2035}), .a ({key_s1[2], key_s0[2]}), .c ({signal_4748, signal_1231}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1378 ( .s (reset), .b ({signal_4672, signal_2034}), .a ({key_s1[3], key_s0[3]}), .c ({signal_4750, signal_1233}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1381 ( .s (reset), .b ({signal_4673, signal_2033}), .a ({key_s1[4], key_s0[4]}), .c ({signal_4752, signal_1235}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1384 ( .s (reset), .b ({signal_4813, signal_2032}), .a ({key_s1[5], key_s0[5]}), .c ({signal_4876, signal_1237}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1387 ( .s (reset), .b ({signal_4814, signal_2031}), .a ({key_s1[6], key_s0[6]}), .c ({signal_4878, signal_1239}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1390 ( .s (reset), .b ({signal_4674, signal_2030}), .a ({key_s1[7], key_s0[7]}), .c ({signal_4754, signal_1241}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1393 ( .s (reset), .b ({signal_4675, signal_2029}), .a ({key_s1[8], key_s0[8]}), .c ({signal_4756, signal_1243}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1396 ( .s (reset), .b ({signal_4815, signal_2028}), .a ({key_s1[9], key_s0[9]}), .c ({signal_4880, signal_1245}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1399 ( .s (reset), .b ({signal_4676, signal_2027}), .a ({key_s1[10], key_s0[10]}), .c ({signal_4758, signal_1247}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1402 ( .s (reset), .b ({signal_4677, signal_2026}), .a ({key_s1[11], key_s0[11]}), .c ({signal_4760, signal_1249}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1405 ( .s (reset), .b ({signal_4678, signal_2025}), .a ({key_s1[12], key_s0[12]}), .c ({signal_4762, signal_1251}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1408 ( .s (reset), .b ({signal_4816, signal_2024}), .a ({key_s1[13], key_s0[13]}), .c ({signal_4882, signal_1253}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1411 ( .s (reset), .b ({signal_4817, signal_2023}), .a ({key_s1[14], key_s0[14]}), .c ({signal_4884, signal_1255}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1414 ( .s (reset), .b ({signal_4679, signal_2022}), .a ({key_s1[15], key_s0[15]}), .c ({signal_4764, signal_1257}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1417 ( .s (reset), .b ({signal_4680, signal_2021}), .a ({key_s1[16], key_s0[16]}), .c ({signal_4766, signal_1259}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1420 ( .s (reset), .b ({signal_4818, signal_2020}), .a ({key_s1[17], key_s0[17]}), .c ({signal_4886, signal_1261}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1423 ( .s (reset), .b ({signal_4681, signal_2019}), .a ({key_s1[18], key_s0[18]}), .c ({signal_4768, signal_1263}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1426 ( .s (reset), .b ({signal_4682, signal_2018}), .a ({key_s1[19], key_s0[19]}), .c ({signal_4770, signal_1265}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1429 ( .s (reset), .b ({signal_4683, signal_2017}), .a ({key_s1[20], key_s0[20]}), .c ({signal_4772, signal_1267}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1432 ( .s (reset), .b ({signal_4819, signal_2016}), .a ({key_s1[21], key_s0[21]}), .c ({signal_4888, signal_1269}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1435 ( .s (reset), .b ({signal_4820, signal_2015}), .a ({key_s1[22], key_s0[22]}), .c ({signal_4890, signal_1271}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1438 ( .s (reset), .b ({signal_4684, signal_2014}), .a ({key_s1[23], key_s0[23]}), .c ({signal_4774, signal_1273}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1441 ( .s (reset), .b ({signal_4821, signal_2013}), .a ({key_s1[24], key_s0[24]}), .c ({signal_4892, signal_1275}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1444 ( .s (reset), .b ({signal_4907, signal_2012}), .a ({key_s1[25], key_s0[25]}), .c ({signal_4919, signal_1277}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1447 ( .s (reset), .b ({signal_4822, signal_2011}), .a ({key_s1[26], key_s0[26]}), .c ({signal_4894, signal_1279}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1450 ( .s (reset), .b ({signal_4823, signal_2010}), .a ({key_s1[27], key_s0[27]}), .c ({signal_4896, signal_1281}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1453 ( .s (reset), .b ({signal_4824, signal_2009}), .a ({key_s1[28], key_s0[28]}), .c ({signal_4898, signal_1283}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1456 ( .s (reset), .b ({signal_4908, signal_2008}), .a ({key_s1[29], key_s0[29]}), .c ({signal_4921, signal_1285}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1459 ( .s (reset), .b ({signal_4909, signal_2007}), .a ({key_s1[30], key_s0[30]}), .c ({signal_4923, signal_1287}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1462 ( .s (reset), .b ({signal_4825, signal_2006}), .a ({key_s1[31], key_s0[31]}), .c ({signal_4900, signal_1289}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1465 ( .s (reset), .b ({signal_4505, signal_2005}), .a ({key_s1[32], key_s0[32]}), .c ({signal_4590, signal_1291}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1468 ( .s (reset), .b ({signal_4685, signal_2004}), .a ({key_s1[33], key_s0[33]}), .c ({signal_4776, signal_1293}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1471 ( .s (reset), .b ({signal_4506, signal_2003}), .a ({key_s1[34], key_s0[34]}), .c ({signal_4592, signal_1295}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1474 ( .s (reset), .b ({signal_4507, signal_2002}), .a ({key_s1[35], key_s0[35]}), .c ({signal_4594, signal_1297}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1477 ( .s (reset), .b ({signal_4508, signal_2001}), .a ({key_s1[36], key_s0[36]}), .c ({signal_4596, signal_1299}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1480 ( .s (reset), .b ({signal_4686, signal_2000}), .a ({key_s1[37], key_s0[37]}), .c ({signal_4778, signal_1301}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1483 ( .s (reset), .b ({signal_4687, signal_1999}), .a ({key_s1[38], key_s0[38]}), .c ({signal_4780, signal_1303}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1486 ( .s (reset), .b ({signal_4509, signal_1998}), .a ({key_s1[39], key_s0[39]}), .c ({signal_4598, signal_1305}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1489 ( .s (reset), .b ({signal_4510, signal_1997}), .a ({key_s1[40], key_s0[40]}), .c ({signal_4600, signal_1307}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1492 ( .s (reset), .b ({signal_4688, signal_1996}), .a ({key_s1[41], key_s0[41]}), .c ({signal_4782, signal_1309}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1495 ( .s (reset), .b ({signal_4511, signal_1995}), .a ({key_s1[42], key_s0[42]}), .c ({signal_4602, signal_1311}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1498 ( .s (reset), .b ({signal_4512, signal_1994}), .a ({key_s1[43], key_s0[43]}), .c ({signal_4604, signal_1313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1501 ( .s (reset), .b ({signal_4513, signal_1993}), .a ({key_s1[44], key_s0[44]}), .c ({signal_4606, signal_1315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1504 ( .s (reset), .b ({signal_4689, signal_1992}), .a ({key_s1[45], key_s0[45]}), .c ({signal_4784, signal_1317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1507 ( .s (reset), .b ({signal_4690, signal_1991}), .a ({key_s1[46], key_s0[46]}), .c ({signal_4786, signal_1319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1510 ( .s (reset), .b ({signal_4514, signal_1990}), .a ({key_s1[47], key_s0[47]}), .c ({signal_4608, signal_1321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1513 ( .s (reset), .b ({signal_4515, signal_1989}), .a ({key_s1[48], key_s0[48]}), .c ({signal_4610, signal_1323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1516 ( .s (reset), .b ({signal_4691, signal_1988}), .a ({key_s1[49], key_s0[49]}), .c ({signal_4788, signal_1325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1519 ( .s (reset), .b ({signal_4516, signal_1987}), .a ({key_s1[50], key_s0[50]}), .c ({signal_4612, signal_1327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1522 ( .s (reset), .b ({signal_4517, signal_1986}), .a ({key_s1[51], key_s0[51]}), .c ({signal_4614, signal_1329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1525 ( .s (reset), .b ({signal_4518, signal_1985}), .a ({key_s1[52], key_s0[52]}), .c ({signal_4616, signal_1331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1528 ( .s (reset), .b ({signal_4692, signal_1984}), .a ({key_s1[53], key_s0[53]}), .c ({signal_4790, signal_1333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1531 ( .s (reset), .b ({signal_4693, signal_1983}), .a ({key_s1[54], key_s0[54]}), .c ({signal_4792, signal_1335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1534 ( .s (reset), .b ({signal_4519, signal_1982}), .a ({key_s1[55], key_s0[55]}), .c ({signal_4618, signal_1337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1537 ( .s (reset), .b ({signal_4694, signal_1981}), .a ({key_s1[56], key_s0[56]}), .c ({signal_4794, signal_1339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1540 ( .s (reset), .b ({signal_4826, signal_1980}), .a ({key_s1[57], key_s0[57]}), .c ({signal_4902, signal_1341}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1543 ( .s (reset), .b ({signal_4695, signal_1979}), .a ({key_s1[58], key_s0[58]}), .c ({signal_4796, signal_1343}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1546 ( .s (reset), .b ({signal_4696, signal_1978}), .a ({key_s1[59], key_s0[59]}), .c ({signal_4798, signal_1345}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1549 ( .s (reset), .b ({signal_4697, signal_1977}), .a ({key_s1[60], key_s0[60]}), .c ({signal_4800, signal_1347}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1552 ( .s (reset), .b ({signal_4827, signal_1976}), .a ({key_s1[61], key_s0[61]}), .c ({signal_4904, signal_1349}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1555 ( .s (reset), .b ({signal_4828, signal_1975}), .a ({key_s1[62], key_s0[62]}), .c ({signal_4906, signal_1351}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1558 ( .s (reset), .b ({signal_4698, signal_1974}), .a ({key_s1[63], key_s0[63]}), .c ({signal_4802, signal_1353}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1561 ( .s (reset), .b ({signal_4345, signal_1973}), .a ({key_s1[64], key_s0[64]}), .c ({signal_4416, signal_1355}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1564 ( .s (reset), .b ({signal_4520, signal_1972}), .a ({key_s1[65], key_s0[65]}), .c ({signal_4620, signal_1357}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1567 ( .s (reset), .b ({signal_4346, signal_1971}), .a ({key_s1[66], key_s0[66]}), .c ({signal_4418, signal_1359}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1570 ( .s (reset), .b ({signal_4347, signal_1970}), .a ({key_s1[67], key_s0[67]}), .c ({signal_4420, signal_1361}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1573 ( .s (reset), .b ({signal_4348, signal_1969}), .a ({key_s1[68], key_s0[68]}), .c ({signal_4422, signal_1363}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1576 ( .s (reset), .b ({signal_4521, signal_1968}), .a ({key_s1[69], key_s0[69]}), .c ({signal_4622, signal_1365}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1579 ( .s (reset), .b ({signal_4522, signal_1967}), .a ({key_s1[70], key_s0[70]}), .c ({signal_4624, signal_1367}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1582 ( .s (reset), .b ({signal_4349, signal_1966}), .a ({key_s1[71], key_s0[71]}), .c ({signal_4424, signal_1369}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1585 ( .s (reset), .b ({signal_4350, signal_1965}), .a ({key_s1[72], key_s0[72]}), .c ({signal_4426, signal_1371}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1588 ( .s (reset), .b ({signal_4523, signal_1964}), .a ({key_s1[73], key_s0[73]}), .c ({signal_4626, signal_1373}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1591 ( .s (reset), .b ({signal_4351, signal_1963}), .a ({key_s1[74], key_s0[74]}), .c ({signal_4428, signal_1375}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1594 ( .s (reset), .b ({signal_4352, signal_1962}), .a ({key_s1[75], key_s0[75]}), .c ({signal_4430, signal_1377}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1597 ( .s (reset), .b ({signal_4353, signal_1961}), .a ({key_s1[76], key_s0[76]}), .c ({signal_4432, signal_1379}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1600 ( .s (reset), .b ({signal_4524, signal_1960}), .a ({key_s1[77], key_s0[77]}), .c ({signal_4628, signal_1381}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1603 ( .s (reset), .b ({signal_4525, signal_1959}), .a ({key_s1[78], key_s0[78]}), .c ({signal_4630, signal_1383}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1606 ( .s (reset), .b ({signal_4354, signal_1958}), .a ({key_s1[79], key_s0[79]}), .c ({signal_4434, signal_1385}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1609 ( .s (reset), .b ({signal_4355, signal_1957}), .a ({key_s1[80], key_s0[80]}), .c ({signal_4436, signal_1387}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1612 ( .s (reset), .b ({signal_4526, signal_1956}), .a ({key_s1[81], key_s0[81]}), .c ({signal_4632, signal_1389}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1615 ( .s (reset), .b ({signal_4356, signal_1955}), .a ({key_s1[82], key_s0[82]}), .c ({signal_4438, signal_1391}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1618 ( .s (reset), .b ({signal_4357, signal_1954}), .a ({key_s1[83], key_s0[83]}), .c ({signal_4440, signal_1393}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1621 ( .s (reset), .b ({signal_4358, signal_1953}), .a ({key_s1[84], key_s0[84]}), .c ({signal_4442, signal_1395}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1624 ( .s (reset), .b ({signal_4527, signal_1952}), .a ({key_s1[85], key_s0[85]}), .c ({signal_4634, signal_1397}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1627 ( .s (reset), .b ({signal_4528, signal_1951}), .a ({key_s1[86], key_s0[86]}), .c ({signal_4636, signal_1399}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1630 ( .s (reset), .b ({signal_4359, signal_1950}), .a ({key_s1[87], key_s0[87]}), .c ({signal_4444, signal_1401}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1633 ( .s (reset), .b ({signal_4529, signal_1949}), .a ({key_s1[88], key_s0[88]}), .c ({signal_4638, signal_1403}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1636 ( .s (reset), .b ({signal_4699, signal_1948}), .a ({key_s1[89], key_s0[89]}), .c ({signal_4804, signal_1405}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1639 ( .s (reset), .b ({signal_4530, signal_1947}), .a ({key_s1[90], key_s0[90]}), .c ({signal_4640, signal_1407}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1642 ( .s (reset), .b ({signal_4531, signal_1946}), .a ({key_s1[91], key_s0[91]}), .c ({signal_4642, signal_1409}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1645 ( .s (reset), .b ({signal_4532, signal_1945}), .a ({key_s1[92], key_s0[92]}), .c ({signal_4644, signal_1411}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1648 ( .s (reset), .b ({signal_4700, signal_1944}), .a ({key_s1[93], key_s0[93]}), .c ({signal_4806, signal_1413}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1651 ( .s (reset), .b ({signal_4701, signal_1943}), .a ({key_s1[94], key_s0[94]}), .c ({signal_4808, signal_1415}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1654 ( .s (reset), .b ({signal_4533, signal_1942}), .a ({key_s1[95], key_s0[95]}), .c ({signal_4646, signal_1417}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1657 ( .s (reset), .b ({signal_4236, signal_1941}), .a ({key_s1[96], key_s0[96]}), .c ({signal_4284, signal_1419}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1660 ( .s (reset), .b ({signal_4360, signal_1940}), .a ({key_s1[97], key_s0[97]}), .c ({signal_4446, signal_1421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1663 ( .s (reset), .b ({signal_4237, signal_1939}), .a ({key_s1[98], key_s0[98]}), .c ({signal_4286, signal_1423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1666 ( .s (reset), .b ({signal_4238, signal_1938}), .a ({key_s1[99], key_s0[99]}), .c ({signal_4288, signal_1425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1669 ( .s (reset), .b ({signal_4239, signal_1937}), .a ({key_s1[100], key_s0[100]}), .c ({signal_4290, signal_1427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1672 ( .s (reset), .b ({signal_4361, signal_1936}), .a ({key_s1[101], key_s0[101]}), .c ({signal_4448, signal_1429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1675 ( .s (reset), .b ({signal_4362, signal_1935}), .a ({key_s1[102], key_s0[102]}), .c ({signal_4450, signal_1431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1678 ( .s (reset), .b ({signal_4240, signal_1934}), .a ({key_s1[103], key_s0[103]}), .c ({signal_4292, signal_1433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1681 ( .s (reset), .b ({signal_4241, signal_1933}), .a ({key_s1[104], key_s0[104]}), .c ({signal_4294, signal_1435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1684 ( .s (reset), .b ({signal_4363, signal_1932}), .a ({key_s1[105], key_s0[105]}), .c ({signal_4452, signal_1437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1687 ( .s (reset), .b ({signal_4242, signal_1931}), .a ({key_s1[106], key_s0[106]}), .c ({signal_4296, signal_1439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1690 ( .s (reset), .b ({signal_4243, signal_1930}), .a ({key_s1[107], key_s0[107]}), .c ({signal_4298, signal_1441}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1693 ( .s (reset), .b ({signal_4244, signal_1929}), .a ({key_s1[108], key_s0[108]}), .c ({signal_4300, signal_1443}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1696 ( .s (reset), .b ({signal_4364, signal_1928}), .a ({key_s1[109], key_s0[109]}), .c ({signal_4454, signal_1445}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1699 ( .s (reset), .b ({signal_4365, signal_1927}), .a ({key_s1[110], key_s0[110]}), .c ({signal_4456, signal_1447}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1702 ( .s (reset), .b ({signal_4245, signal_1926}), .a ({key_s1[111], key_s0[111]}), .c ({signal_4302, signal_1449}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1705 ( .s (reset), .b ({signal_4246, signal_1925}), .a ({key_s1[112], key_s0[112]}), .c ({signal_4304, signal_1451}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1708 ( .s (reset), .b ({signal_4366, signal_1924}), .a ({key_s1[113], key_s0[113]}), .c ({signal_4458, signal_1453}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1711 ( .s (reset), .b ({signal_4247, signal_1923}), .a ({key_s1[114], key_s0[114]}), .c ({signal_4306, signal_1455}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1714 ( .s (reset), .b ({signal_4248, signal_1922}), .a ({key_s1[115], key_s0[115]}), .c ({signal_4308, signal_1457}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1717 ( .s (reset), .b ({signal_4249, signal_1921}), .a ({key_s1[116], key_s0[116]}), .c ({signal_4310, signal_1459}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1720 ( .s (reset), .b ({signal_4367, signal_1920}), .a ({key_s1[117], key_s0[117]}), .c ({signal_4460, signal_1461}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1723 ( .s (reset), .b ({signal_4368, signal_1919}), .a ({key_s1[118], key_s0[118]}), .c ({signal_4462, signal_1463}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1726 ( .s (reset), .b ({signal_4250, signal_1918}), .a ({key_s1[119], key_s0[119]}), .c ({signal_4312, signal_1465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1729 ( .s (reset), .b ({signal_4369, signal_1917}), .a ({key_s1[120], key_s0[120]}), .c ({signal_4464, signal_1467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1732 ( .s (reset), .b ({signal_4534, signal_1916}), .a ({key_s1[121], key_s0[121]}), .c ({signal_4648, signal_1469}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1735 ( .s (reset), .b ({signal_4370, signal_1915}), .a ({key_s1[122], key_s0[122]}), .c ({signal_4466, signal_1471}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1738 ( .s (reset), .b ({signal_4371, signal_1914}), .a ({key_s1[123], key_s0[123]}), .c ({signal_4468, signal_1473}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1741 ( .s (reset), .b ({signal_4372, signal_1913}), .a ({key_s1[124], key_s0[124]}), .c ({signal_4470, signal_1475}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1744 ( .s (reset), .b ({signal_4535, signal_1912}), .a ({key_s1[125], key_s0[125]}), .c ({signal_4650, signal_1477}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1747 ( .s (reset), .b ({signal_4536, signal_1911}), .a ({key_s1[126], key_s0[126]}), .c ({signal_4652, signal_1479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1750 ( .s (reset), .b ({signal_4373, signal_1910}), .a ({key_s1[127], key_s0[127]}), .c ({signal_4472, signal_1481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1751 ( .a ({signal_3302, signal_1800}), .b ({signal_4476, signal_2228}), .c ({signal_4653, signal_2260}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1752 ( .a ({signal_3269, signal_1801}), .b ({signal_4314, signal_2229}), .c ({signal_4473, signal_2261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1753 ( .a ({signal_3236, signal_1786}), .b ({signal_4315, signal_2230}), .c ({signal_4474, signal_2262}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1754 ( .a ({signal_3203, signal_1787}), .b ({signal_4478, signal_2231}), .c ({signal_4654, signal_2263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1755 ( .a ({signal_3170, signal_1788}), .b ({signal_4479, signal_2232}), .c ({signal_4655, signal_2264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1756 ( .a ({signal_3137, signal_1789}), .b ({signal_4318, signal_2233}), .c ({signal_4475, signal_2265}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1757 ( .a ({signal_3110, signal_2124}), .b ({signal_4313, signal_2196}), .c ({signal_4476, signal_2228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1758 ( .a ({signal_3215, signal_2092}), .b ({signal_4229, signal_2164}), .c ({signal_4313, signal_2196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1759 ( .a ({signal_3107, signal_2125}), .b ({signal_4204, signal_2197}), .c ({signal_4314, signal_2229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1760 ( .a ({signal_3212, signal_2093}), .b ({signal_4151, signal_2165}), .c ({signal_4204, signal_2197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1761 ( .a ({signal_3104, signal_1790}), .b ({signal_4319, signal_2234}), .c ({signal_4477, signal_2266}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1762 ( .a ({signal_3101, signal_2126}), .b ({signal_4205, signal_2198}), .c ({signal_4315, signal_2230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1763 ( .a ({signal_3209, signal_2094}), .b ({signal_4152, signal_2166}), .c ({signal_4205, signal_2198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1764 ( .a ({signal_3098, signal_2127}), .b ({signal_4316, signal_2199}), .c ({signal_4478, signal_2231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1765 ( .a ({signal_3206, signal_2095}), .b ({signal_4230, signal_2167}), .c ({signal_4316, signal_2199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1766 ( .a ({signal_3095, signal_2128}), .b ({signal_4317, signal_2200}), .c ({signal_4479, signal_2232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1767 ( .a ({signal_3200, signal_2096}), .b ({signal_4231, signal_2168}), .c ({signal_4317, signal_2200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1768 ( .a ({signal_3092, signal_2129}), .b ({signal_4206, signal_2201}), .c ({signal_4318, signal_2233}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1769 ( .a ({signal_3197, signal_2097}), .b ({signal_4153, signal_2169}), .c ({signal_4206, signal_2201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1770 ( .a ({signal_3089, signal_2130}), .b ({signal_4207, signal_2202}), .c ({signal_4319, signal_2234}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1771 ( .a ({signal_3194, signal_2098}), .b ({signal_4140, signal_2170}), .c ({signal_4207, signal_2202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1772 ( .a ({signal_3299, signal_2066}), .b ({signal_4137, signal_2334}), .c ({signal_4140, signal_2170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1773 ( .a ({signal_3077, signal_1778}), .b ({signal_4480, signal_2206}), .c ({signal_4656, signal_2238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1774 ( .a ({signal_3182, signal_2102}), .b ({signal_4320, signal_2174}), .c ({signal_4480, signal_2206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1775 ( .a ({signal_3287, signal_2070}), .b ({signal_4217, signal_2142}), .c ({signal_4320, signal_2174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1776 ( .a ({signal_3074, signal_1779}), .b ({signal_4657, signal_2207}), .c ({signal_4809, signal_2239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1777 ( .a ({signal_3179, signal_2103}), .b ({signal_4481, signal_2175}), .c ({signal_4657, signal_2207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1778 ( .a ({signal_3284, signal_2071}), .b ({signal_4339, signal_2143}), .c ({signal_4481, signal_2175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1779 ( .a ({signal_3071, signal_1791}), .b ({signal_4321, signal_2235}), .c ({signal_4482, signal_2267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1780 ( .a ({signal_3086, signal_2131}), .b ({signal_4208, signal_2203}), .c ({signal_4321, signal_2235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1781 ( .a ({signal_3191, signal_2099}), .b ({signal_4141, signal_2171}), .c ({signal_4208, signal_2203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1782 ( .a ({signal_3296, signal_2067}), .b ({signal_4138, signal_2335}), .c ({signal_4141, signal_2171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1783 ( .a ({signal_3068, signal_1780}), .b ({signal_4658, signal_2208}), .c ({signal_4810, signal_2240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1784 ( .a ({signal_3176, signal_2104}), .b ({signal_4483, signal_2176}), .c ({signal_4658, signal_2208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1785 ( .a ({signal_3281, signal_2072}), .b ({signal_4340, signal_2144}), .c ({signal_4483, signal_2176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1786 ( .a ({signal_3065, signal_1781}), .b ({signal_4484, signal_2209}), .c ({signal_4659, signal_2241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1787 ( .a ({signal_3173, signal_2105}), .b ({signal_4322, signal_2177}), .c ({signal_4484, signal_2209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1788 ( .a ({signal_3278, signal_2073}), .b ({signal_4218, signal_2145}), .c ({signal_4322, signal_2177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1789 ( .a ({signal_3062, signal_1782}), .b ({signal_4485, signal_2210}), .c ({signal_4660, signal_2242}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1790 ( .a ({signal_3167, signal_2106}), .b ({signal_4323, signal_2178}), .c ({signal_4485, signal_2210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1791 ( .a ({signal_3275, signal_2074}), .b ({signal_4219, signal_2146}), .c ({signal_4323, signal_2178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1792 ( .a ({signal_3059, signal_1783}), .b ({signal_4486, signal_2211}), .c ({signal_4661, signal_2243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1793 ( .a ({signal_3164, signal_2107}), .b ({signal_4324, signal_2179}), .c ({signal_4486, signal_2211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1794 ( .a ({signal_3272, signal_2075}), .b ({signal_4220, signal_2147}), .c ({signal_4324, signal_2179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1795 ( .a ({signal_3056, signal_1784}), .b ({signal_4662, signal_2212}), .c ({signal_4811, signal_2244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1796 ( .a ({signal_3161, signal_2108}), .b ({signal_4487, signal_2180}), .c ({signal_4662, signal_2212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1797 ( .a ({signal_3266, signal_2076}), .b ({signal_4341, signal_2148}), .c ({signal_4487, signal_2180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1798 ( .a ({signal_3053, signal_1785}), .b ({signal_4488, signal_2213}), .c ({signal_4663, signal_2245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1799 ( .a ({signal_3158, signal_2109}), .b ({signal_4325, signal_2181}), .c ({signal_4488, signal_2213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1800 ( .a ({signal_3263, signal_2077}), .b ({signal_4221, signal_2149}), .c ({signal_4325, signal_2181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1801 ( .a ({signal_3050, signal_1802}), .b ({signal_4326, signal_2214}), .c ({signal_4489, signal_2246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1802 ( .a ({signal_3155, signal_2110}), .b ({signal_4209, signal_2182}), .c ({signal_4326, signal_2214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1803 ( .a ({signal_3260, signal_2078}), .b ({signal_4142, signal_2150}), .c ({signal_4209, signal_2182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1804 ( .a ({signal_3047, signal_1803}), .b ({signal_4490, signal_2215}), .c ({signal_4664, signal_2247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1805 ( .a ({signal_3152, signal_2111}), .b ({signal_4327, signal_2183}), .c ({signal_4490, signal_2215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1806 ( .a ({signal_3257, signal_2079}), .b ({signal_4223, signal_2151}), .c ({signal_4327, signal_2183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1807 ( .a ({signal_3044, signal_1804}), .b ({signal_4491, signal_2216}), .c ({signal_4665, signal_2248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1808 ( .a ({signal_3149, signal_2112}), .b ({signal_4328, signal_2184}), .c ({signal_4491, signal_2216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1809 ( .a ({signal_3254, signal_2080}), .b ({signal_4224, signal_2152}), .c ({signal_4328, signal_2184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1810 ( .a ({signal_3041, signal_1805}), .b ({signal_4329, signal_2217}), .c ({signal_4492, signal_2249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1811 ( .a ({signal_3146, signal_2113}), .b ({signal_4210, signal_2185}), .c ({signal_4329, signal_2217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1812 ( .a ({signal_3251, signal_2081}), .b ({signal_4143, signal_2153}), .c ({signal_4210, signal_2185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1813 ( .a ({signal_3038, signal_1792}), .b ({signal_4493, signal_2236}), .c ({signal_4666, signal_2268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1814 ( .a ({signal_3083, signal_2132}), .b ({signal_4330, signal_2204}), .c ({signal_4493, signal_2236}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1815 ( .a ({signal_3188, signal_2100}), .b ({signal_4211, signal_2172}), .c ({signal_4330, signal_2204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1816 ( .a ({signal_3293, signal_2068}), .b ({signal_4171, signal_2336}), .c ({signal_4211, signal_2172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1817 ( .a ({signal_3035, signal_1806}), .b ({signal_4331, signal_2218}), .c ({signal_4494, signal_2250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1818 ( .a ({signal_3143, signal_2114}), .b ({signal_4212, signal_2186}), .c ({signal_4331, signal_2218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1819 ( .a ({signal_3248, signal_2082}), .b ({signal_4144, signal_2154}), .c ({signal_4212, signal_2186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1820 ( .a ({signal_3032, signal_1807}), .b ({signal_4332, signal_2219}), .c ({signal_4495, signal_2251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1821 ( .a ({signal_3140, signal_2115}), .b ({signal_4213, signal_2187}), .c ({signal_4332, signal_2219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1822 ( .a ({signal_3245, signal_2083}), .b ({signal_4145, signal_2155}), .c ({signal_4213, signal_2187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1823 ( .a ({signal_3029, signal_1808}), .b ({signal_4496, signal_2220}), .c ({signal_4667, signal_2252}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1824 ( .a ({signal_3134, signal_2116}), .b ({signal_4333, signal_2188}), .c ({signal_4496, signal_2220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1825 ( .a ({signal_3242, signal_2084}), .b ({signal_4225, signal_2156}), .c ({signal_4333, signal_2188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1826 ( .a ({signal_3026, signal_1809}), .b ({signal_4334, signal_2221}), .c ({signal_4497, signal_2253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1827 ( .a ({signal_3131, signal_2117}), .b ({signal_4214, signal_2189}), .c ({signal_4334, signal_2221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1828 ( .a ({signal_3239, signal_2085}), .b ({signal_4146, signal_2157}), .c ({signal_4214, signal_2189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1829 ( .a ({signal_3023, signal_1794}), .b ({signal_4335, signal_2222}), .c ({signal_4498, signal_2254}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1830 ( .a ({signal_3128, signal_2118}), .b ({signal_4215, signal_2190}), .c ({signal_4335, signal_2222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1831 ( .a ({signal_3233, signal_2086}), .b ({signal_4147, signal_2158}), .c ({signal_4215, signal_2190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1832 ( .a ({signal_3020, signal_1795}), .b ({signal_4499, signal_2223}), .c ({signal_4668, signal_2255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1833 ( .a ({signal_3125, signal_2119}), .b ({signal_4336, signal_2191}), .c ({signal_4499, signal_2223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1834 ( .a ({signal_3230, signal_2087}), .b ({signal_4226, signal_2159}), .c ({signal_4336, signal_2191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1835 ( .a ({signal_3017, signal_1796}), .b ({signal_4500, signal_2224}), .c ({signal_4669, signal_2256}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1836 ( .a ({signal_3122, signal_2120}), .b ({signal_4337, signal_2192}), .c ({signal_4500, signal_2224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1837 ( .a ({signal_3227, signal_2088}), .b ({signal_4228, signal_2160}), .c ({signal_4337, signal_2192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1838 ( .a ({signal_3014, signal_1797}), .b ({signal_4338, signal_2225}), .c ({signal_4501, signal_2257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1839 ( .a ({signal_3119, signal_2121}), .b ({signal_4216, signal_2193}), .c ({signal_4338, signal_2225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1840 ( .a ({signal_3224, signal_2089}), .b ({signal_4148, signal_2161}), .c ({signal_4216, signal_2193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1841 ( .a ({signal_3011, signal_2038}), .b ({signal_4155, signal_2306}), .c ({signal_4217, signal_2142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1842 ( .a ({signal_3008, signal_2039}), .b ({signal_4233, signal_2307}), .c ({signal_4339, signal_2143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1843 ( .a ({signal_3005, signal_2040}), .b ({signal_4234, signal_2308}), .c ({signal_4340, signal_2144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1844 ( .a ({signal_3002, signal_2041}), .b ({signal_4156, signal_2309}), .c ({signal_4218, signal_2145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1845 ( .a ({signal_2999, signal_2042}), .b ({signal_4157, signal_2310}), .c ({signal_4219, signal_2146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1846 ( .a ({signal_2996, signal_2043}), .b ({signal_4158, signal_2311}), .c ({signal_4220, signal_2147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1847 ( .a ({signal_2993, signal_2044}), .b ({signal_4235, signal_2312}), .c ({signal_4341, signal_2148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1848 ( .a ({signal_2990, signal_2045}), .b ({signal_4159, signal_2313}), .c ({signal_4221, signal_2149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1849 ( .a ({signal_2987, signal_1798}), .b ({signal_4342, signal_2226}), .c ({signal_4502, signal_2258}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1850 ( .a ({signal_3116, signal_2122}), .b ({signal_4222, signal_2194}), .c ({signal_4342, signal_2226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1851 ( .a ({signal_3221, signal_2090}), .b ({signal_4149, signal_2162}), .c ({signal_4222, signal_2194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1852 ( .a ({signal_2984, signal_2046}), .b ({signal_4119, signal_2314}), .c ({signal_4142, signal_2150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1853 ( .a ({signal_2981, signal_2047}), .b ({signal_4163, signal_2315}), .c ({signal_4223, signal_2151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1854 ( .a ({signal_2978, signal_2048}), .b ({signal_4164, signal_2316}), .c ({signal_4224, signal_2152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1855 ( .a ({signal_2975, signal_2049}), .b ({signal_4122, signal_2317}), .c ({signal_4143, signal_2153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1856 ( .a ({signal_2972, signal_2050}), .b ({signal_4123, signal_2318}), .c ({signal_4144, signal_2154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1857 ( .a ({signal_2969, signal_2051}), .b ({signal_4124, signal_2319}), .c ({signal_4145, signal_2155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1858 ( .a ({signal_2966, signal_2052}), .b ({signal_4165, signal_2320}), .c ({signal_4225, signal_2156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1859 ( .a ({signal_2963, signal_2053}), .b ({signal_4109, signal_2321}), .c ({signal_4146, signal_2157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1860 ( .a ({signal_2960, signal_2054}), .b ({signal_4126, signal_2322}), .c ({signal_4147, signal_2158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1861 ( .a ({signal_2957, signal_2055}), .b ({signal_4166, signal_2323}), .c ({signal_4226, signal_2159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1862 ( .a ({signal_2954, signal_1799}), .b ({signal_4343, signal_2227}), .c ({signal_4503, signal_2259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1863 ( .a ({signal_3113, signal_2123}), .b ({signal_4227, signal_2195}), .c ({signal_4343, signal_2227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1864 ( .a ({signal_3218, signal_2091}), .b ({signal_4150, signal_2163}), .c ({signal_4227, signal_2195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1865 ( .a ({signal_2951, signal_2056}), .b ({signal_4167, signal_2324}), .c ({signal_4228, signal_2160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1866 ( .a ({signal_2948, signal_2057}), .b ({signal_4129, signal_2325}), .c ({signal_4148, signal_2161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1867 ( .a ({signal_2945, signal_2058}), .b ({signal_4130, signal_2326}), .c ({signal_4149, signal_2162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1868 ( .a ({signal_2942, signal_2059}), .b ({signal_4131, signal_2327}), .c ({signal_4150, signal_2163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1869 ( .a ({signal_2939, signal_2060}), .b ({signal_4168, signal_2328}), .c ({signal_4229, signal_2164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1870 ( .a ({signal_2936, signal_2061}), .b ({signal_4110, signal_2329}), .c ({signal_4151, signal_2165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1871 ( .a ({signal_2933, signal_2062}), .b ({signal_4133, signal_2330}), .c ({signal_4152, signal_2166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1872 ( .a ({signal_2930, signal_2063}), .b ({signal_4169, signal_2331}), .c ({signal_4230, signal_2167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1873 ( .a ({signal_2927, signal_2064}), .b ({signal_4170, signal_2332}), .c ({signal_4231, signal_2168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1874 ( .a ({signal_2924, signal_2065}), .b ({signal_4136, signal_2333}), .c ({signal_4153, signal_2169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1875 ( .a ({signal_2921, signal_1793}), .b ({signal_4344, signal_2237}), .c ({signal_4504, signal_2269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1876 ( .a ({signal_3080, signal_2133}), .b ({signal_4232, signal_2205}), .c ({signal_4344, signal_2237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1877 ( .a ({signal_3185, signal_2101}), .b ({signal_4154, signal_2173}), .c ({signal_4232, signal_2205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1878 ( .a ({signal_3290, signal_2069}), .b ({signal_4111, signal_2337}), .c ({signal_4154, signal_2173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1879 ( .a ({1'b0, signal_2134}), .b ({signal_4112, signal_2305}), .c ({signal_4155, signal_2306}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1880 ( .a ({1'b0, signal_2135}), .b ({signal_4160, signal_2298}), .c ({signal_4233, signal_2307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1881 ( .a ({1'b0, signal_2136}), .b ({signal_4161, signal_2299}), .c ({signal_4234, signal_2308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1882 ( .a ({1'b0, signal_2137}), .b ({signal_4115, signal_2300}), .c ({signal_4156, signal_2309}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1883 ( .a ({1'b0, signal_2138}), .b ({signal_4116, signal_1842}), .c ({signal_4157, signal_2310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1884 ( .a ({1'b0, signal_2139}), .b ({signal_4117, signal_1843}), .c ({signal_4158, signal_2311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1885 ( .a ({1'b0, signal_2140}), .b ({signal_4162, signal_2303}), .c ({signal_4235, signal_2312}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1886 ( .a ({1'b0, signal_2141}), .b ({signal_4108, signal_1845}), .c ({signal_4159, signal_2313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1895 ( .s (signal_1489), .b ({signal_2921, signal_1793}), .a ({signal_4504, signal_2269}), .c ({signal_4670, signal_2037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1896 ( .s (signal_1488), .b ({signal_3038, signal_1792}), .a ({signal_4666, signal_2268}), .c ({signal_4812, signal_2036}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1897 ( .s (signal_1487), .b ({signal_3071, signal_1791}), .a ({signal_4482, signal_2267}), .c ({signal_4671, signal_2035}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1898 ( .s (signal_1486), .b ({signal_3104, signal_1790}), .a ({signal_4477, signal_2266}), .c ({signal_4672, signal_2034}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1899 ( .s (signal_1485), .b ({signal_3137, signal_1789}), .a ({signal_4475, signal_2265}), .c ({signal_4673, signal_2033}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1900 ( .s (signal_1484), .b ({signal_3170, signal_1788}), .a ({signal_4655, signal_2264}), .c ({signal_4813, signal_2032}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1901 ( .s (signal_1488), .b ({signal_3203, signal_1787}), .a ({signal_4654, signal_2263}), .c ({signal_4814, signal_2031}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1902 ( .s (signal_1486), .b ({signal_3236, signal_1786}), .a ({signal_4474, signal_2262}), .c ({signal_4674, signal_2030}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1903 ( .s (signal_1489), .b ({signal_3269, signal_1801}), .a ({signal_4473, signal_2261}), .c ({signal_4675, signal_2029}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1904 ( .s (signal_1488), .b ({signal_3302, signal_1800}), .a ({signal_4653, signal_2260}), .c ({signal_4815, signal_2028}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1905 ( .s (signal_1487), .b ({signal_2954, signal_1799}), .a ({signal_4503, signal_2259}), .c ({signal_4676, signal_2027}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1906 ( .s (signal_1486), .b ({signal_2987, signal_1798}), .a ({signal_4502, signal_2258}), .c ({signal_4677, signal_2026}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1907 ( .s (signal_1485), .b ({signal_3014, signal_1797}), .a ({signal_4501, signal_2257}), .c ({signal_4678, signal_2025}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1908 ( .s (signal_1484), .b ({signal_3017, signal_1796}), .a ({signal_4669, signal_2256}), .c ({signal_4816, signal_2024}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1909 ( .s (signal_1485), .b ({signal_3020, signal_1795}), .a ({signal_4668, signal_2255}), .c ({signal_4817, signal_2023}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1910 ( .s (signal_1485), .b ({signal_3023, signal_1794}), .a ({signal_4498, signal_2254}), .c ({signal_4679, signal_2022}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1911 ( .s (signal_1489), .b ({signal_3026, signal_1809}), .a ({signal_4497, signal_2253}), .c ({signal_4680, signal_2021}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1912 ( .s (signal_1488), .b ({signal_3029, signal_1808}), .a ({signal_4667, signal_2252}), .c ({signal_4818, signal_2020}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1913 ( .s (signal_1487), .b ({signal_3032, signal_1807}), .a ({signal_4495, signal_2251}), .c ({signal_4681, signal_2019}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1914 ( .s (signal_1486), .b ({signal_3035, signal_1806}), .a ({signal_4494, signal_2250}), .c ({signal_4682, signal_2018}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1915 ( .s (signal_1484), .b ({signal_3041, signal_1805}), .a ({signal_4492, signal_2249}), .c ({signal_4683, signal_2017}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1916 ( .s (signal_1484), .b ({signal_3044, signal_1804}), .a ({signal_4665, signal_2248}), .c ({signal_4819, signal_2016}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1917 ( .s (signal_1489), .b ({signal_3047, signal_1803}), .a ({signal_4664, signal_2247}), .c ({signal_4820, signal_2015}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1918 ( .s (signal_1488), .b ({signal_3050, signal_1802}), .a ({signal_4489, signal_2246}), .c ({signal_4684, signal_2014}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1919 ( .s (signal_1487), .b ({signal_3053, signal_1785}), .a ({signal_4663, signal_2245}), .c ({signal_4821, signal_2013}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1920 ( .s (signal_1486), .b ({signal_3056, signal_1784}), .a ({signal_4811, signal_2244}), .c ({signal_4907, signal_2012}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1921 ( .s (signal_1485), .b ({signal_3059, signal_1783}), .a ({signal_4661, signal_2243}), .c ({signal_4822, signal_2011}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1922 ( .s (signal_1484), .b ({signal_3062, signal_1782}), .a ({signal_4660, signal_2242}), .c ({signal_4823, signal_2010}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1923 ( .s (signal_1489), .b ({signal_3065, signal_1781}), .a ({signal_4659, signal_2241}), .c ({signal_4824, signal_2009}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1924 ( .s (signal_1489), .b ({signal_3068, signal_1780}), .a ({signal_4810, signal_2240}), .c ({signal_4908, signal_2008}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1925 ( .s (signal_1488), .b ({signal_3074, signal_1779}), .a ({signal_4809, signal_2239}), .c ({signal_4909, signal_2007}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1926 ( .s (signal_1487), .b ({signal_3077, signal_1778}), .a ({signal_4656, signal_2238}), .c ({signal_4825, signal_2006}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1927 ( .s (signal_1488), .b ({signal_3080, signal_2133}), .a ({signal_4344, signal_2237}), .c ({signal_4505, signal_2005}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1928 ( .s (signal_1487), .b ({signal_3083, signal_2132}), .a ({signal_4493, signal_2236}), .c ({signal_4685, signal_2004}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1929 ( .s (signal_1486), .b ({signal_3086, signal_2131}), .a ({signal_4321, signal_2235}), .c ({signal_4506, signal_2003}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1930 ( .s (signal_1485), .b ({signal_3089, signal_2130}), .a ({signal_4319, signal_2234}), .c ({signal_4507, signal_2002}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1931 ( .s (signal_1484), .b ({signal_3092, signal_2129}), .a ({signal_4318, signal_2233}), .c ({signal_4508, signal_2001}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1932 ( .s (signal_1489), .b ({signal_3095, signal_2128}), .a ({signal_4479, signal_2232}), .c ({signal_4686, signal_2000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1933 ( .s (signal_1488), .b ({signal_3098, signal_2127}), .a ({signal_4478, signal_2231}), .c ({signal_4687, signal_1999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1934 ( .s (signal_1487), .b ({signal_3101, signal_2126}), .a ({signal_4315, signal_2230}), .c ({signal_4509, signal_1998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1935 ( .s (signal_1486), .b ({signal_3107, signal_2125}), .a ({signal_4314, signal_2229}), .c ({signal_4510, signal_1997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1936 ( .s (signal_1485), .b ({signal_3110, signal_2124}), .a ({signal_4476, signal_2228}), .c ({signal_4688, signal_1996}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1937 ( .s (signal_1484), .b ({signal_3113, signal_2123}), .a ({signal_4343, signal_2227}), .c ({signal_4511, signal_1995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1938 ( .s (signal_1489), .b ({signal_3116, signal_2122}), .a ({signal_4342, signal_2226}), .c ({signal_4512, signal_1994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1939 ( .s (signal_1484), .b ({signal_3119, signal_2121}), .a ({signal_4338, signal_2225}), .c ({signal_4513, signal_1993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1940 ( .s (signal_1484), .b ({signal_3122, signal_2120}), .a ({signal_4500, signal_2224}), .c ({signal_4689, signal_1992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1941 ( .s (signal_1484), .b ({signal_3125, signal_2119}), .a ({signal_4499, signal_2223}), .c ({signal_4690, signal_1991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1942 ( .s (signal_1484), .b ({signal_3128, signal_2118}), .a ({signal_4335, signal_2222}), .c ({signal_4514, signal_1990}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1943 ( .s (signal_1484), .b ({signal_3131, signal_2117}), .a ({signal_4334, signal_2221}), .c ({signal_4515, signal_1989}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1944 ( .s (signal_1484), .b ({signal_3134, signal_2116}), .a ({signal_4496, signal_2220}), .c ({signal_4691, signal_1988}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1945 ( .s (signal_1484), .b ({signal_3140, signal_2115}), .a ({signal_4332, signal_2219}), .c ({signal_4516, signal_1987}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1946 ( .s (signal_1484), .b ({signal_3143, signal_2114}), .a ({signal_4331, signal_2218}), .c ({signal_4517, signal_1986}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1947 ( .s (signal_1484), .b ({signal_3146, signal_2113}), .a ({signal_4329, signal_2217}), .c ({signal_4518, signal_1985}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1948 ( .s (signal_1484), .b ({signal_3149, signal_2112}), .a ({signal_4491, signal_2216}), .c ({signal_4692, signal_1984}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1949 ( .s (signal_1484), .b ({signal_3152, signal_2111}), .a ({signal_4490, signal_2215}), .c ({signal_4693, signal_1983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1950 ( .s (signal_1484), .b ({signal_3155, signal_2110}), .a ({signal_4326, signal_2214}), .c ({signal_4519, signal_1982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1951 ( .s (signal_1485), .b ({signal_3158, signal_2109}), .a ({signal_4488, signal_2213}), .c ({signal_4694, signal_1981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1952 ( .s (signal_1485), .b ({signal_3161, signal_2108}), .a ({signal_4662, signal_2212}), .c ({signal_4826, signal_1980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1953 ( .s (signal_1485), .b ({signal_3164, signal_2107}), .a ({signal_4486, signal_2211}), .c ({signal_4695, signal_1979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1954 ( .s (signal_1485), .b ({signal_3167, signal_2106}), .a ({signal_4485, signal_2210}), .c ({signal_4696, signal_1978}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1955 ( .s (signal_1485), .b ({signal_3173, signal_2105}), .a ({signal_4484, signal_2209}), .c ({signal_4697, signal_1977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1956 ( .s (signal_1485), .b ({signal_3176, signal_2104}), .a ({signal_4658, signal_2208}), .c ({signal_4827, signal_1976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1957 ( .s (signal_1485), .b ({signal_3179, signal_2103}), .a ({signal_4657, signal_2207}), .c ({signal_4828, signal_1975}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1958 ( .s (signal_1485), .b ({signal_3182, signal_2102}), .a ({signal_4480, signal_2206}), .c ({signal_4698, signal_1974}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1959 ( .s (signal_1485), .b ({signal_3185, signal_2101}), .a ({signal_4232, signal_2205}), .c ({signal_4345, signal_1973}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1960 ( .s (signal_1485), .b ({signal_3188, signal_2100}), .a ({signal_4330, signal_2204}), .c ({signal_4520, signal_1972}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1961 ( .s (signal_1485), .b ({signal_3191, signal_2099}), .a ({signal_4208, signal_2203}), .c ({signal_4346, signal_1971}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1962 ( .s (signal_1485), .b ({signal_3194, signal_2098}), .a ({signal_4207, signal_2202}), .c ({signal_4347, signal_1970}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1963 ( .s (signal_1486), .b ({signal_3197, signal_2097}), .a ({signal_4206, signal_2201}), .c ({signal_4348, signal_1969}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1964 ( .s (signal_1486), .b ({signal_3200, signal_2096}), .a ({signal_4317, signal_2200}), .c ({signal_4521, signal_1968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1965 ( .s (signal_1486), .b ({signal_3206, signal_2095}), .a ({signal_4316, signal_2199}), .c ({signal_4522, signal_1967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1966 ( .s (signal_1486), .b ({signal_3209, signal_2094}), .a ({signal_4205, signal_2198}), .c ({signal_4349, signal_1966}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1967 ( .s (signal_1486), .b ({signal_3212, signal_2093}), .a ({signal_4204, signal_2197}), .c ({signal_4350, signal_1965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1968 ( .s (signal_1486), .b ({signal_3215, signal_2092}), .a ({signal_4313, signal_2196}), .c ({signal_4523, signal_1964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1969 ( .s (signal_1486), .b ({signal_3218, signal_2091}), .a ({signal_4227, signal_2195}), .c ({signal_4351, signal_1963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1970 ( .s (signal_1486), .b ({signal_3221, signal_2090}), .a ({signal_4222, signal_2194}), .c ({signal_4352, signal_1962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1971 ( .s (signal_1486), .b ({signal_3224, signal_2089}), .a ({signal_4216, signal_2193}), .c ({signal_4353, signal_1961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1972 ( .s (signal_1486), .b ({signal_3227, signal_2088}), .a ({signal_4337, signal_2192}), .c ({signal_4524, signal_1960}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1973 ( .s (signal_1486), .b ({signal_3230, signal_2087}), .a ({signal_4336, signal_2191}), .c ({signal_4525, signal_1959}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1974 ( .s (signal_1486), .b ({signal_3233, signal_2086}), .a ({signal_4215, signal_2190}), .c ({signal_4354, signal_1958}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1975 ( .s (signal_1487), .b ({signal_3239, signal_2085}), .a ({signal_4214, signal_2189}), .c ({signal_4355, signal_1957}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1976 ( .s (signal_1487), .b ({signal_3242, signal_2084}), .a ({signal_4333, signal_2188}), .c ({signal_4526, signal_1956}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1977 ( .s (signal_1487), .b ({signal_3245, signal_2083}), .a ({signal_4213, signal_2187}), .c ({signal_4356, signal_1955}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1978 ( .s (signal_1487), .b ({signal_3248, signal_2082}), .a ({signal_4212, signal_2186}), .c ({signal_4357, signal_1954}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1979 ( .s (signal_1487), .b ({signal_3251, signal_2081}), .a ({signal_4210, signal_2185}), .c ({signal_4358, signal_1953}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1980 ( .s (signal_1487), .b ({signal_3254, signal_2080}), .a ({signal_4328, signal_2184}), .c ({signal_4527, signal_1952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1981 ( .s (signal_1487), .b ({signal_3257, signal_2079}), .a ({signal_4327, signal_2183}), .c ({signal_4528, signal_1951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1982 ( .s (signal_1487), .b ({signal_3260, signal_2078}), .a ({signal_4209, signal_2182}), .c ({signal_4359, signal_1950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1983 ( .s (signal_1487), .b ({signal_3263, signal_2077}), .a ({signal_4325, signal_2181}), .c ({signal_4529, signal_1949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1984 ( .s (signal_1487), .b ({signal_3266, signal_2076}), .a ({signal_4487, signal_2180}), .c ({signal_4699, signal_1948}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1985 ( .s (signal_1487), .b ({signal_3272, signal_2075}), .a ({signal_4324, signal_2179}), .c ({signal_4530, signal_1947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1986 ( .s (signal_1487), .b ({signal_3275, signal_2074}), .a ({signal_4323, signal_2178}), .c ({signal_4531, signal_1946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1987 ( .s (signal_1488), .b ({signal_3278, signal_2073}), .a ({signal_4322, signal_2177}), .c ({signal_4532, signal_1945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1988 ( .s (signal_1488), .b ({signal_3281, signal_2072}), .a ({signal_4483, signal_2176}), .c ({signal_4700, signal_1944}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1989 ( .s (signal_1488), .b ({signal_3284, signal_2071}), .a ({signal_4481, signal_2175}), .c ({signal_4701, signal_1943}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1990 ( .s (signal_1488), .b ({signal_3287, signal_2070}), .a ({signal_4320, signal_2174}), .c ({signal_4533, signal_1942}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1991 ( .s (signal_1488), .b ({signal_3290, signal_2069}), .a ({signal_4154, signal_2173}), .c ({signal_4236, signal_1941}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1992 ( .s (signal_1488), .b ({signal_3293, signal_2068}), .a ({signal_4211, signal_2172}), .c ({signal_4360, signal_1940}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1993 ( .s (signal_1488), .b ({signal_3296, signal_2067}), .a ({signal_4141, signal_2171}), .c ({signal_4237, signal_1939}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1994 ( .s (signal_1488), .b ({signal_3299, signal_2066}), .a ({signal_4140, signal_2170}), .c ({signal_4238, signal_1938}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1995 ( .s (signal_1488), .b ({signal_2924, signal_2065}), .a ({signal_4153, signal_2169}), .c ({signal_4239, signal_1937}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1996 ( .s (signal_1488), .b ({signal_2927, signal_2064}), .a ({signal_4231, signal_2168}), .c ({signal_4361, signal_1936}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1997 ( .s (signal_1488), .b ({signal_2930, signal_2063}), .a ({signal_4230, signal_2167}), .c ({signal_4362, signal_1935}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1998 ( .s (signal_1488), .b ({signal_2933, signal_2062}), .a ({signal_4152, signal_2166}), .c ({signal_4240, signal_1934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1999 ( .s (signal_1489), .b ({signal_2936, signal_2061}), .a ({signal_4151, signal_2165}), .c ({signal_4241, signal_1933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2000 ( .s (signal_1489), .b ({signal_2939, signal_2060}), .a ({signal_4229, signal_2164}), .c ({signal_4363, signal_1932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2001 ( .s (signal_1489), .b ({signal_2942, signal_2059}), .a ({signal_4150, signal_2163}), .c ({signal_4242, signal_1931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2002 ( .s (signal_1489), .b ({signal_2945, signal_2058}), .a ({signal_4149, signal_2162}), .c ({signal_4243, signal_1930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2003 ( .s (signal_1489), .b ({signal_2948, signal_2057}), .a ({signal_4148, signal_2161}), .c ({signal_4244, signal_1929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2004 ( .s (signal_1489), .b ({signal_2951, signal_2056}), .a ({signal_4228, signal_2160}), .c ({signal_4364, signal_1928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2005 ( .s (signal_1489), .b ({signal_2957, signal_2055}), .a ({signal_4226, signal_2159}), .c ({signal_4365, signal_1927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2006 ( .s (signal_1489), .b ({signal_2960, signal_2054}), .a ({signal_4147, signal_2158}), .c ({signal_4245, signal_1926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2007 ( .s (signal_1489), .b ({signal_2963, signal_2053}), .a ({signal_4146, signal_2157}), .c ({signal_4246, signal_1925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2008 ( .s (signal_1489), .b ({signal_2966, signal_2052}), .a ({signal_4225, signal_2156}), .c ({signal_4366, signal_1924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2009 ( .s (signal_1489), .b ({signal_2969, signal_2051}), .a ({signal_4145, signal_2155}), .c ({signal_4247, signal_1923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2010 ( .s (signal_1489), .b ({signal_2972, signal_2050}), .a ({signal_4144, signal_2154}), .c ({signal_4248, signal_1922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2011 ( .s (signal_1490), .b ({signal_2975, signal_2049}), .a ({signal_4143, signal_2153}), .c ({signal_4249, signal_1921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2012 ( .s (signal_1490), .b ({signal_2978, signal_2048}), .a ({signal_4224, signal_2152}), .c ({signal_4367, signal_1920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2013 ( .s (signal_1490), .b ({signal_2981, signal_2047}), .a ({signal_4223, signal_2151}), .c ({signal_4368, signal_1919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2014 ( .s (signal_1490), .b ({signal_2984, signal_2046}), .a ({signal_4142, signal_2150}), .c ({signal_4250, signal_1918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2015 ( .s (signal_1490), .b ({signal_2990, signal_2045}), .a ({signal_4221, signal_2149}), .c ({signal_4369, signal_1917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2016 ( .s (signal_1490), .b ({signal_2993, signal_2044}), .a ({signal_4341, signal_2148}), .c ({signal_4534, signal_1916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2017 ( .s (signal_1490), .b ({signal_2996, signal_2043}), .a ({signal_4220, signal_2147}), .c ({signal_4370, signal_1915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2018 ( .s (signal_1490), .b ({signal_2999, signal_2042}), .a ({signal_4219, signal_2146}), .c ({signal_4371, signal_1914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2019 ( .s (signal_1490), .b ({signal_3002, signal_2041}), .a ({signal_4218, signal_2145}), .c ({signal_4372, signal_1913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2020 ( .s (signal_1490), .b ({signal_3005, signal_2040}), .a ({signal_4340, signal_2144}), .c ({signal_4535, signal_1912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2021 ( .s (signal_1490), .b ({signal_3008, signal_2039}), .a ({signal_4339, signal_2143}), .c ({signal_4536, signal_1911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2022 ( .s (signal_1490), .b ({signal_3011, signal_2038}), .a ({signal_4217, signal_2142}), .c ({signal_4373, signal_1910}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2325 ( .a ({signal_3720, signal_2430}), .b ({signal_3879, signal_2589}), .clk (clk), .r (Fresh[64]), .c ({signal_3892, signal_2602}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2326 ( .a ({signal_3305, signal_1841}), .b ({signal_3878, signal_2588}), .clk (clk), .r (Fresh[65]), .c ({signal_3893, signal_2603}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2327 ( .a ({signal_3665, signal_2375}), .b ({signal_3877, signal_2587}), .clk (clk), .r (Fresh[66]), .c ({signal_3894, signal_2604}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2328 ( .a ({signal_3723, signal_2433}), .b ({signal_3876, signal_2586}), .clk (clk), .r (Fresh[67]), .c ({signal_3895, signal_2605}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2329 ( .a ({signal_3725, signal_2435}), .b ({signal_3879, signal_2589}), .clk (clk), .r (Fresh[68]), .c ({signal_3896, signal_2606}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2330 ( .a ({signal_3669, signal_2379}), .b ({signal_3878, signal_2588}), .clk (clk), .r (Fresh[69]), .c ({signal_3897, signal_2607}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2331 ( .a ({signal_3670, signal_2380}), .b ({signal_3877, signal_2587}), .clk (clk), .r (Fresh[70]), .c ({signal_3898, signal_2608}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2332 ( .a ({signal_3724, signal_2434}), .b ({signal_3876, signal_2586}), .clk (clk), .r (Fresh[71]), .c ({signal_3899, signal_2609}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2333 ( .a ({signal_3727, signal_2437}), .b ({signal_3883, signal_2593}), .clk (clk), .r (Fresh[72]), .c ({signal_3900, signal_2610}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2334 ( .a ({signal_3304, signal_1833}), .b ({signal_3882, signal_2592}), .clk (clk), .r (Fresh[73]), .c ({signal_3901, signal_2611}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2335 ( .a ({signal_3673, signal_2383}), .b ({signal_3881, signal_2591}), .clk (clk), .r (Fresh[74]), .c ({signal_3902, signal_2612}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2336 ( .a ({signal_3730, signal_2440}), .b ({signal_3880, signal_2590}), .clk (clk), .r (Fresh[75]), .c ({signal_3903, signal_2613}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2337 ( .a ({signal_3732, signal_2442}), .b ({signal_3883, signal_2593}), .clk (clk), .r (Fresh[76]), .c ({signal_3904, signal_2614}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2338 ( .a ({signal_3677, signal_2387}), .b ({signal_3882, signal_2592}), .clk (clk), .r (Fresh[77]), .c ({signal_3905, signal_2615}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2339 ( .a ({signal_3678, signal_2388}), .b ({signal_3881, signal_2591}), .clk (clk), .r (Fresh[78]), .c ({signal_3906, signal_2616}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2340 ( .a ({signal_3731, signal_2441}), .b ({signal_3880, signal_2590}), .clk (clk), .r (Fresh[79]), .c ({signal_3907, signal_2617}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2341 ( .a ({signal_3734, signal_2444}), .b ({signal_3887, signal_2597}), .clk (clk), .r (Fresh[80]), .c ({signal_3908, signal_2618}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2342 ( .a ({signal_3320, signal_1825}), .b ({signal_3886, signal_2596}), .clk (clk), .r (Fresh[81]), .c ({signal_3909, signal_2619}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2343 ( .a ({signal_3681, signal_2391}), .b ({signal_3885, signal_2595}), .clk (clk), .r (Fresh[82]), .c ({signal_3910, signal_2620}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2344 ( .a ({signal_3737, signal_2447}), .b ({signal_3884, signal_2594}), .clk (clk), .r (Fresh[83]), .c ({signal_3911, signal_2621}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2345 ( .a ({signal_3739, signal_2449}), .b ({signal_3887, signal_2597}), .clk (clk), .r (Fresh[84]), .c ({signal_3912, signal_2622}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2346 ( .a ({signal_3685, signal_2395}), .b ({signal_3886, signal_2596}), .clk (clk), .r (Fresh[85]), .c ({signal_3913, signal_2623}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2347 ( .a ({signal_3686, signal_2396}), .b ({signal_3885, signal_2595}), .clk (clk), .r (Fresh[86]), .c ({signal_3914, signal_2624}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2348 ( .a ({signal_3738, signal_2448}), .b ({signal_3884, signal_2594}), .clk (clk), .r (Fresh[87]), .c ({signal_3915, signal_2625}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2349 ( .a ({signal_3741, signal_2451}), .b ({signal_3891, signal_2601}), .clk (clk), .r (Fresh[88]), .c ({signal_3916, signal_2626}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2350 ( .a ({signal_3328, signal_1817}), .b ({signal_3890, signal_2600}), .clk (clk), .r (Fresh[89]), .c ({signal_3917, signal_2627}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2351 ( .a ({signal_3689, signal_2399}), .b ({signal_3889, signal_2599}), .clk (clk), .r (Fresh[90]), .c ({signal_3918, signal_2628}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2352 ( .a ({signal_3744, signal_2454}), .b ({signal_3888, signal_2598}), .clk (clk), .r (Fresh[91]), .c ({signal_3919, signal_2629}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2353 ( .a ({signal_3746, signal_2456}), .b ({signal_3891, signal_2601}), .clk (clk), .r (Fresh[92]), .c ({signal_3920, signal_2630}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2354 ( .a ({signal_3693, signal_2403}), .b ({signal_3890, signal_2600}), .clk (clk), .r (Fresh[93]), .c ({signal_3921, signal_2631}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2355 ( .a ({signal_3694, signal_2404}), .b ({signal_3889, signal_2599}), .clk (clk), .r (Fresh[94]), .c ({signal_3922, signal_2632}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2356 ( .a ({signal_3745, signal_2455}), .b ({signal_3888, signal_2598}), .clk (clk), .r (Fresh[95]), .c ({signal_3923, signal_2633}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2373 ( .a ({signal_3664, signal_2374}), .b ({signal_3927, signal_2637}), .clk (clk), .r (Fresh[96]), .c ({signal_3940, signal_2650}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2374 ( .a ({signal_3668, signal_2378}), .b ({signal_3926, signal_2636}), .clk (clk), .r (Fresh[97]), .c ({signal_3941, signal_2651}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2375 ( .a ({signal_3667, signal_2377}), .b ({signal_3925, signal_2635}), .clk (clk), .r (Fresh[98]), .c ({signal_3942, signal_2652}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2376 ( .a ({signal_3721, signal_2431}), .b ({signal_3924, signal_2634}), .clk (clk), .r (Fresh[99]), .c ({signal_3943, signal_2653}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2377 ( .a ({signal_3666, signal_2376}), .b ({signal_3927, signal_2637}), .clk (clk), .r (Fresh[100]), .c ({signal_3944, signal_2654}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2378 ( .a ({signal_3630, signal_2340}), .b ({signal_3926, signal_2636}), .clk (clk), .r (Fresh[101]), .c ({signal_3945, signal_2655}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2379 ( .a ({signal_3628, signal_2338}), .b ({signal_3925, signal_2635}), .clk (clk), .r (Fresh[102]), .c ({signal_3946, signal_2656}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2380 ( .a ({signal_3629, signal_2339}), .b ({signal_3924, signal_2634}), .clk (clk), .r (Fresh[103]), .c ({signal_3947, signal_2657}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2381 ( .a ({signal_3672, signal_2382}), .b ({signal_3931, signal_2641}), .clk (clk), .r (Fresh[104]), .c ({signal_3948, signal_2658}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2382 ( .a ({signal_3676, signal_2386}), .b ({signal_3930, signal_2640}), .clk (clk), .r (Fresh[105]), .c ({signal_3949, signal_2659}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2383 ( .a ({signal_3675, signal_2385}), .b ({signal_3929, signal_2639}), .clk (clk), .r (Fresh[106]), .c ({signal_3950, signal_2660}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2384 ( .a ({signal_3728, signal_2438}), .b ({signal_3928, signal_2638}), .clk (clk), .r (Fresh[107]), .c ({signal_3951, signal_2661}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2385 ( .a ({signal_3674, signal_2384}), .b ({signal_3931, signal_2641}), .clk (clk), .r (Fresh[108]), .c ({signal_3952, signal_2662}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2386 ( .a ({signal_3639, signal_2349}), .b ({signal_3930, signal_2640}), .clk (clk), .r (Fresh[109]), .c ({signal_3953, signal_2663}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2387 ( .a ({signal_3637, signal_2347}), .b ({signal_3929, signal_2639}), .clk (clk), .r (Fresh[110]), .c ({signal_3954, signal_2664}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2388 ( .a ({signal_3638, signal_2348}), .b ({signal_3928, signal_2638}), .clk (clk), .r (Fresh[111]), .c ({signal_3955, signal_2665}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2389 ( .a ({signal_3680, signal_2390}), .b ({signal_3935, signal_2645}), .clk (clk), .r (Fresh[112]), .c ({signal_3956, signal_2666}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2390 ( .a ({signal_3684, signal_2394}), .b ({signal_3934, signal_2644}), .clk (clk), .r (Fresh[113]), .c ({signal_3957, signal_2667}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2391 ( .a ({signal_3683, signal_2393}), .b ({signal_3933, signal_2643}), .clk (clk), .r (Fresh[114]), .c ({signal_3958, signal_2668}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2392 ( .a ({signal_3735, signal_2445}), .b ({signal_3932, signal_2642}), .clk (clk), .r (Fresh[115]), .c ({signal_3959, signal_2669}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2393 ( .a ({signal_3682, signal_2392}), .b ({signal_3935, signal_2645}), .clk (clk), .r (Fresh[116]), .c ({signal_3960, signal_2670}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2394 ( .a ({signal_3648, signal_2358}), .b ({signal_3934, signal_2644}), .clk (clk), .r (Fresh[117]), .c ({signal_3961, signal_2671}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2395 ( .a ({signal_3646, signal_2356}), .b ({signal_3933, signal_2643}), .clk (clk), .r (Fresh[118]), .c ({signal_3962, signal_2672}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2396 ( .a ({signal_3647, signal_2357}), .b ({signal_3932, signal_2642}), .clk (clk), .r (Fresh[119]), .c ({signal_3963, signal_2673}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2397 ( .a ({signal_3688, signal_2398}), .b ({signal_3939, signal_2649}), .clk (clk), .r (Fresh[120]), .c ({signal_3964, signal_2674}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2398 ( .a ({signal_3692, signal_2402}), .b ({signal_3938, signal_2648}), .clk (clk), .r (Fresh[121]), .c ({signal_3965, signal_2675}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2399 ( .a ({signal_3691, signal_2401}), .b ({signal_3937, signal_2647}), .clk (clk), .r (Fresh[122]), .c ({signal_3966, signal_2676}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2400 ( .a ({signal_3742, signal_2452}), .b ({signal_3936, signal_2646}), .clk (clk), .r (Fresh[123]), .c ({signal_3967, signal_2677}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2401 ( .a ({signal_3690, signal_2400}), .b ({signal_3939, signal_2649}), .clk (clk), .r (Fresh[124]), .c ({signal_3968, signal_2678}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2402 ( .a ({signal_3657, signal_2367}), .b ({signal_3938, signal_2648}), .clk (clk), .r (Fresh[125]), .c ({signal_3969, signal_2679}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2403 ( .a ({signal_3655, signal_2365}), .b ({signal_3937, signal_2647}), .clk (clk), .r (Fresh[126]), .c ({signal_3970, signal_2680}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2404 ( .a ({signal_3656, signal_2366}), .b ({signal_3936, signal_2646}), .clk (clk), .r (Fresh[127]), .c ({signal_3971, signal_2681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2406 ( .a ({signal_3894, signal_2604}), .b ({signal_3896, signal_2606}), .c ({signal_3973, signal_2683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2407 ( .a ({signal_3895, signal_2605}), .b ({signal_3898, signal_2608}), .c ({signal_3974, signal_2684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2408 ( .a ({signal_3893, signal_2603}), .b ({signal_3895, signal_2605}), .c ({signal_3975, signal_2685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2410 ( .a ({signal_3902, signal_2612}), .b ({signal_3904, signal_2614}), .c ({signal_3977, signal_2687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2411 ( .a ({signal_3903, signal_2613}), .b ({signal_3906, signal_2616}), .c ({signal_3978, signal_2688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2412 ( .a ({signal_3901, signal_2611}), .b ({signal_3903, signal_2613}), .c ({signal_3979, signal_2689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2414 ( .a ({signal_3910, signal_2620}), .b ({signal_3912, signal_2622}), .c ({signal_3981, signal_2691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2415 ( .a ({signal_3911, signal_2621}), .b ({signal_3914, signal_2624}), .c ({signal_3982, signal_2692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2416 ( .a ({signal_3909, signal_2619}), .b ({signal_3911, signal_2621}), .c ({signal_3983, signal_2693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2418 ( .a ({signal_3918, signal_2628}), .b ({signal_3920, signal_2630}), .c ({signal_3985, signal_2695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2419 ( .a ({signal_3919, signal_2629}), .b ({signal_3922, signal_2632}), .c ({signal_3986, signal_2696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2420 ( .a ({signal_3917, signal_2627}), .b ({signal_3919, signal_2629}), .c ({signal_3987, signal_2697}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2421 ( .a ({signal_3671, signal_2381}), .b ({signal_3972, signal_2682}), .clk (clk), .r (Fresh[128]), .c ({signal_3988, signal_2698}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2422 ( .a ({signal_3631, signal_2341}), .b ({signal_3972, signal_2682}), .clk (clk), .r (Fresh[129]), .c ({signal_3989, signal_2699}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2423 ( .a ({signal_3679, signal_2389}), .b ({signal_3976, signal_2686}), .clk (clk), .r (Fresh[130]), .c ({signal_3990, signal_2700}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2424 ( .a ({signal_3640, signal_2350}), .b ({signal_3976, signal_2686}), .clk (clk), .r (Fresh[131]), .c ({signal_3991, signal_2701}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2425 ( .a ({signal_3687, signal_2397}), .b ({signal_3980, signal_2690}), .clk (clk), .r (Fresh[132]), .c ({signal_3992, signal_2702}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2426 ( .a ({signal_3649, signal_2359}), .b ({signal_3980, signal_2690}), .clk (clk), .r (Fresh[133]), .c ({signal_3993, signal_2703}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2427 ( .a ({signal_3695, signal_2405}), .b ({signal_3984, signal_2694}), .clk (clk), .r (Fresh[134]), .c ({signal_3994, signal_2704}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2428 ( .a ({signal_3658, signal_2368}), .b ({signal_3984, signal_2694}), .clk (clk), .r (Fresh[135]), .c ({signal_3995, signal_2705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2429 ( .a ({signal_3893, signal_2603}), .b ({signal_3940, signal_2650}), .c ({signal_3996, signal_2706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2430 ( .a ({signal_3892, signal_2602}), .b ({signal_3944, signal_2654}), .c ({signal_3997, signal_2707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2431 ( .a ({signal_3943, signal_2653}), .b ({signal_3945, signal_2655}), .c ({signal_3998, signal_2708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2432 ( .a ({signal_3941, signal_2651}), .b ({signal_3946, signal_2656}), .c ({signal_3999, signal_2709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2433 ( .a ({signal_3942, signal_2652}), .b ({signal_3946, signal_2656}), .c ({signal_4000, signal_2710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2434 ( .a ({signal_3944, signal_2654}), .b ({signal_3973, signal_2683}), .c ({signal_4001, signal_2711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2435 ( .a ({signal_3897, signal_2607}), .b ({signal_3973, signal_2683}), .c ({signal_4002, signal_2712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2436 ( .a ({signal_3945, signal_2655}), .b ({signal_3974, signal_2684}), .c ({signal_4003, signal_2713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2437 ( .a ({signal_3901, signal_2611}), .b ({signal_3948, signal_2658}), .c ({signal_4004, signal_2714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2438 ( .a ({signal_3900, signal_2610}), .b ({signal_3952, signal_2662}), .c ({signal_4005, signal_2715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2439 ( .a ({signal_3951, signal_2661}), .b ({signal_3953, signal_2663}), .c ({signal_4006, signal_2716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2440 ( .a ({signal_3949, signal_2659}), .b ({signal_3954, signal_2664}), .c ({signal_4007, signal_2717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2441 ( .a ({signal_3950, signal_2660}), .b ({signal_3954, signal_2664}), .c ({signal_4008, signal_2718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2442 ( .a ({signal_3952, signal_2662}), .b ({signal_3977, signal_2687}), .c ({signal_4009, signal_2719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2443 ( .a ({signal_3905, signal_2615}), .b ({signal_3977, signal_2687}), .c ({signal_4010, signal_2720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2444 ( .a ({signal_3953, signal_2663}), .b ({signal_3978, signal_2688}), .c ({signal_4011, signal_2721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2445 ( .a ({signal_3909, signal_2619}), .b ({signal_3956, signal_2666}), .c ({signal_4012, signal_2722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2446 ( .a ({signal_3908, signal_2618}), .b ({signal_3960, signal_2670}), .c ({signal_4013, signal_2723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2447 ( .a ({signal_3959, signal_2669}), .b ({signal_3961, signal_2671}), .c ({signal_4014, signal_2724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2448 ( .a ({signal_3957, signal_2667}), .b ({signal_3962, signal_2672}), .c ({signal_4015, signal_2725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2449 ( .a ({signal_3958, signal_2668}), .b ({signal_3962, signal_2672}), .c ({signal_4016, signal_2726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2450 ( .a ({signal_3960, signal_2670}), .b ({signal_3981, signal_2691}), .c ({signal_4017, signal_2727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2451 ( .a ({signal_3913, signal_2623}), .b ({signal_3981, signal_2691}), .c ({signal_4018, signal_2728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2452 ( .a ({signal_3961, signal_2671}), .b ({signal_3982, signal_2692}), .c ({signal_4019, signal_2729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2453 ( .a ({signal_3917, signal_2627}), .b ({signal_3964, signal_2674}), .c ({signal_4020, signal_2730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2454 ( .a ({signal_3916, signal_2626}), .b ({signal_3968, signal_2678}), .c ({signal_4021, signal_2731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2455 ( .a ({signal_3967, signal_2677}), .b ({signal_3969, signal_2679}), .c ({signal_4022, signal_2732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2456 ( .a ({signal_3965, signal_2675}), .b ({signal_3970, signal_2680}), .c ({signal_4023, signal_2733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2457 ( .a ({signal_3966, signal_2676}), .b ({signal_3970, signal_2680}), .c ({signal_4024, signal_2734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2458 ( .a ({signal_3968, signal_2678}), .b ({signal_3985, signal_2695}), .c ({signal_4025, signal_2735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2459 ( .a ({signal_3921, signal_2631}), .b ({signal_3985, signal_2695}), .c ({signal_4026, signal_2736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2460 ( .a ({signal_3969, signal_2679}), .b ({signal_3986, signal_2696}), .c ({signal_4027, signal_2737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2461 ( .a ({signal_3946, signal_2656}), .b ({signal_3989, signal_2699}), .c ({signal_4028, signal_2738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2462 ( .a ({signal_3989, signal_2699}), .b ({signal_3999, signal_2709}), .c ({signal_4029, signal_2739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2463 ( .a ({signal_3940, signal_2650}), .b ({signal_3997, signal_2707}), .c ({signal_4030, signal_2740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2464 ( .a ({signal_3942, signal_2652}), .b ({signal_3988, signal_2698}), .c ({signal_4031, signal_2741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2465 ( .a ({signal_3988, signal_2698}), .b ({signal_3998, signal_2708}), .c ({signal_4032, signal_2742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2466 ( .a ({signal_3899, signal_2609}), .b ({signal_3996, signal_2706}), .c ({signal_4033, signal_2743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2467 ( .a ({signal_3947, signal_2657}), .b ({signal_3998, signal_2708}), .c ({signal_4034, signal_2744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2468 ( .a ({signal_3975, signal_2685}), .b ({signal_3997, signal_2707}), .c ({signal_4035, signal_2745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2469 ( .a ({signal_3996, signal_2706}), .b ({signal_4003, signal_2713}), .c ({signal_4036, signal_2746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2470 ( .a ({signal_3954, signal_2664}), .b ({signal_3991, signal_2701}), .c ({signal_4037, signal_2747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2471 ( .a ({signal_3991, signal_2701}), .b ({signal_4007, signal_2717}), .c ({signal_4038, signal_2748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2472 ( .a ({signal_3948, signal_2658}), .b ({signal_4005, signal_2715}), .c ({signal_4039, signal_2749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2473 ( .a ({signal_3950, signal_2660}), .b ({signal_3990, signal_2700}), .c ({signal_4040, signal_2750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2474 ( .a ({signal_3990, signal_2700}), .b ({signal_4006, signal_2716}), .c ({signal_4041, signal_2751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2475 ( .a ({signal_3907, signal_2617}), .b ({signal_4004, signal_2714}), .c ({signal_4042, signal_2752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2476 ( .a ({signal_3955, signal_2665}), .b ({signal_4006, signal_2716}), .c ({signal_4043, signal_2753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2477 ( .a ({signal_3979, signal_2689}), .b ({signal_4005, signal_2715}), .c ({signal_4044, signal_2754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2478 ( .a ({signal_4004, signal_2714}), .b ({signal_4011, signal_2721}), .c ({signal_4045, signal_2755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2479 ( .a ({signal_3962, signal_2672}), .b ({signal_3993, signal_2703}), .c ({signal_4046, signal_2756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2480 ( .a ({signal_3993, signal_2703}), .b ({signal_4015, signal_2725}), .c ({signal_4047, signal_2757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2481 ( .a ({signal_3956, signal_2666}), .b ({signal_4013, signal_2723}), .c ({signal_4048, signal_2758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2482 ( .a ({signal_3958, signal_2668}), .b ({signal_3992, signal_2702}), .c ({signal_4049, signal_2759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2483 ( .a ({signal_3992, signal_2702}), .b ({signal_4014, signal_2724}), .c ({signal_4050, signal_2760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2484 ( .a ({signal_3915, signal_2625}), .b ({signal_4012, signal_2722}), .c ({signal_4051, signal_2761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2485 ( .a ({signal_3963, signal_2673}), .b ({signal_4014, signal_2724}), .c ({signal_4052, signal_2762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2486 ( .a ({signal_3983, signal_2693}), .b ({signal_4013, signal_2723}), .c ({signal_4053, signal_2763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2487 ( .a ({signal_4012, signal_2722}), .b ({signal_4019, signal_2729}), .c ({signal_4054, signal_2764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2488 ( .a ({signal_3970, signal_2680}), .b ({signal_3995, signal_2705}), .c ({signal_4055, signal_2765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2489 ( .a ({signal_3995, signal_2705}), .b ({signal_4023, signal_2733}), .c ({signal_4056, signal_2766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2490 ( .a ({signal_3964, signal_2674}), .b ({signal_4021, signal_2731}), .c ({signal_4057, signal_2767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2491 ( .a ({signal_3966, signal_2676}), .b ({signal_3994, signal_2704}), .c ({signal_4058, signal_2768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2492 ( .a ({signal_3994, signal_2704}), .b ({signal_4022, signal_2732}), .c ({signal_4059, signal_2769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2493 ( .a ({signal_3923, signal_2633}), .b ({signal_4020, signal_2730}), .c ({signal_4060, signal_2770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2494 ( .a ({signal_3971, signal_2681}), .b ({signal_4022, signal_2732}), .c ({signal_4061, signal_2771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2495 ( .a ({signal_3987, signal_2697}), .b ({signal_4021, signal_2731}), .c ({signal_4062, signal_2772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2496 ( .a ({signal_4020, signal_2730}), .b ({signal_4027, signal_2737}), .c ({signal_4063, signal_2773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2497 ( .a ({signal_3894, signal_2604}), .b ({signal_4028, signal_2738}), .c ({signal_4064, signal_2774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2498 ( .a ({signal_3896, signal_2606}), .b ({signal_4028, signal_2738}), .c ({signal_4065, signal_2775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2499 ( .a ({signal_3973, signal_2683}), .b ({signal_4028, signal_2738}), .c ({signal_4066, signal_2776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2500 ( .a ({signal_3973, signal_2683}), .b ({signal_4030, signal_2740}), .c ({signal_4067, signal_2777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2501 ( .a ({signal_4001, signal_2711}), .b ({signal_4031, signal_2741}), .c ({signal_4068, signal_2778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2502 ( .a ({signal_4029, signal_2739}), .b ({signal_4032, signal_2742}), .c ({signal_4069, signal_2779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2503 ( .a ({signal_4030, signal_2740}), .b ({signal_4031, signal_2741}), .c ({signal_4070, signal_2780}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2504 ( .a ({signal_3974, signal_2684}), .b ({signal_4032, signal_2742}), .c ({signal_4071, signal_2781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2505 ( .a ({signal_4000, signal_2710}), .b ({signal_4033, signal_2743}), .c ({signal_4072, signal_2782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2506 ( .a ({signal_4002, signal_2712}), .b ({signal_4033, signal_2743}), .c ({signal_4073, signal_2783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2507 ( .a ({signal_4029, signal_2739}), .b ({signal_4036, signal_2746}), .c ({signal_4074, signal_2784}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2508 ( .a ({signal_3902, signal_2612}), .b ({signal_4037, signal_2747}), .c ({signal_4075, signal_2785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2509 ( .a ({signal_3904, signal_2614}), .b ({signal_4037, signal_2747}), .c ({signal_4076, signal_2786}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2510 ( .a ({signal_3977, signal_2687}), .b ({signal_4037, signal_2747}), .c ({signal_4077, signal_2787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2511 ( .a ({signal_3977, signal_2687}), .b ({signal_4039, signal_2749}), .c ({signal_4078, signal_2788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2512 ( .a ({signal_4009, signal_2719}), .b ({signal_4040, signal_2750}), .c ({signal_4079, signal_2789}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2513 ( .a ({signal_4038, signal_2748}), .b ({signal_4041, signal_2751}), .c ({signal_4080, signal_2790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2514 ( .a ({signal_4039, signal_2749}), .b ({signal_4040, signal_2750}), .c ({signal_4081, signal_2791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2515 ( .a ({signal_3978, signal_2688}), .b ({signal_4041, signal_2751}), .c ({signal_4082, signal_2792}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2516 ( .a ({signal_4008, signal_2718}), .b ({signal_4042, signal_2752}), .c ({signal_4083, signal_2793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2517 ( .a ({signal_4010, signal_2720}), .b ({signal_4042, signal_2752}), .c ({signal_4084, signal_2794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2518 ( .a ({signal_4038, signal_2748}), .b ({signal_4045, signal_2755}), .c ({signal_4085, signal_2795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2519 ( .a ({signal_3910, signal_2620}), .b ({signal_4046, signal_2756}), .c ({signal_4086, signal_2796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2520 ( .a ({signal_3912, signal_2622}), .b ({signal_4046, signal_2756}), .c ({signal_4087, signal_2797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2521 ( .a ({signal_3981, signal_2691}), .b ({signal_4046, signal_2756}), .c ({signal_4088, signal_2798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2522 ( .a ({signal_3981, signal_2691}), .b ({signal_4048, signal_2758}), .c ({signal_4089, signal_2799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2523 ( .a ({signal_4017, signal_2727}), .b ({signal_4049, signal_2759}), .c ({signal_4090, signal_2800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2524 ( .a ({signal_4047, signal_2757}), .b ({signal_4050, signal_2760}), .c ({signal_4091, signal_2801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2525 ( .a ({signal_4048, signal_2758}), .b ({signal_4049, signal_2759}), .c ({signal_4092, signal_2802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2526 ( .a ({signal_3982, signal_2692}), .b ({signal_4050, signal_2760}), .c ({signal_4093, signal_2803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2527 ( .a ({signal_4016, signal_2726}), .b ({signal_4051, signal_2761}), .c ({signal_4094, signal_2804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2528 ( .a ({signal_4018, signal_2728}), .b ({signal_4051, signal_2761}), .c ({signal_4095, signal_2805}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2529 ( .a ({signal_4047, signal_2757}), .b ({signal_4054, signal_2764}), .c ({signal_4096, signal_2806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2530 ( .a ({signal_3918, signal_2628}), .b ({signal_4055, signal_2765}), .c ({signal_4097, signal_2807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2531 ( .a ({signal_3920, signal_2630}), .b ({signal_4055, signal_2765}), .c ({signal_4098, signal_2808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2532 ( .a ({signal_3985, signal_2695}), .b ({signal_4055, signal_2765}), .c ({signal_4099, signal_2809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2533 ( .a ({signal_3985, signal_2695}), .b ({signal_4057, signal_2767}), .c ({signal_4100, signal_2810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2534 ( .a ({signal_4025, signal_2735}), .b ({signal_4058, signal_2768}), .c ({signal_4101, signal_2811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2535 ( .a ({signal_4056, signal_2766}), .b ({signal_4059, signal_2769}), .c ({signal_4102, signal_2812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2536 ( .a ({signal_4057, signal_2767}), .b ({signal_4058, signal_2768}), .c ({signal_4103, signal_2813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2537 ( .a ({signal_3986, signal_2696}), .b ({signal_4059, signal_2769}), .c ({signal_4104, signal_2814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2538 ( .a ({signal_4024, signal_2734}), .b ({signal_4060, signal_2770}), .c ({signal_4105, signal_2815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2539 ( .a ({signal_4026, signal_2736}), .b ({signal_4060, signal_2770}), .c ({signal_4106, signal_2816}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2540 ( .a ({signal_4056, signal_2766}), .b ({signal_4063, signal_2773}), .c ({signal_4107, signal_2817}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2541 ( .a ({signal_4074, signal_2784}), .b ({signal_4108, signal_1845}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2542 ( .a ({signal_4085, signal_2795}), .b ({signal_4109, signal_2321}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2543 ( .a ({signal_4096, signal_2806}), .b ({signal_4110, signal_2329}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2544 ( .a ({signal_4107, signal_2817}), .b ({signal_4111, signal_2337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2545 ( .a ({signal_4029, signal_2739}), .b ({signal_4068, signal_2778}), .c ({signal_4112, signal_2305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2546 ( .a ({signal_4065, signal_2775}), .b ({signal_4070, signal_2780}), .c ({signal_4113, signal_2818}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2547 ( .a ({signal_4034, signal_2744}), .b ({signal_4072, signal_2782}), .c ({signal_4114, signal_2819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2548 ( .a ({signal_4029, signal_2739}), .b ({signal_4067, signal_2777}), .c ({signal_4115, signal_2300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2549 ( .a ({signal_4035, signal_2745}), .b ({signal_4066, signal_2776}), .c ({signal_4116, signal_1842}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2550 ( .a ({signal_4069, signal_2779}), .b ({signal_4073, signal_2783}), .c ({signal_4117, signal_1843}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2551 ( .a ({signal_4064, signal_2774}), .b ({signal_4071, signal_2781}), .c ({signal_4118, signal_2820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2552 ( .a ({signal_4038, signal_2748}), .b ({signal_4079, signal_2789}), .c ({signal_4119, signal_2314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2553 ( .a ({signal_4076, signal_2786}), .b ({signal_4081, signal_2791}), .c ({signal_4120, signal_2821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2554 ( .a ({signal_4043, signal_2753}), .b ({signal_4083, signal_2793}), .c ({signal_4121, signal_2822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2555 ( .a ({signal_4038, signal_2748}), .b ({signal_4078, signal_2788}), .c ({signal_4122, signal_2317}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2556 ( .a ({signal_4044, signal_2754}), .b ({signal_4077, signal_2787}), .c ({signal_4123, signal_2318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2557 ( .a ({signal_4080, signal_2790}), .b ({signal_4084, signal_2794}), .c ({signal_4124, signal_2319}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2558 ( .a ({signal_4075, signal_2785}), .b ({signal_4082, signal_2792}), .c ({signal_4125, signal_2823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2559 ( .a ({signal_4047, signal_2757}), .b ({signal_4090, signal_2800}), .c ({signal_4126, signal_2322}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2560 ( .a ({signal_4087, signal_2797}), .b ({signal_4092, signal_2802}), .c ({signal_4127, signal_2824}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2561 ( .a ({signal_4052, signal_2762}), .b ({signal_4094, signal_2804}), .c ({signal_4128, signal_2825}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2562 ( .a ({signal_4047, signal_2757}), .b ({signal_4089, signal_2799}), .c ({signal_4129, signal_2325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2563 ( .a ({signal_4053, signal_2763}), .b ({signal_4088, signal_2798}), .c ({signal_4130, signal_2326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2564 ( .a ({signal_4091, signal_2801}), .b ({signal_4095, signal_2805}), .c ({signal_4131, signal_2327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2565 ( .a ({signal_4086, signal_2796}), .b ({signal_4093, signal_2803}), .c ({signal_4132, signal_2826}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2566 ( .a ({signal_4056, signal_2766}), .b ({signal_4101, signal_2811}), .c ({signal_4133, signal_2330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2567 ( .a ({signal_4098, signal_2808}), .b ({signal_4103, signal_2813}), .c ({signal_4134, signal_2827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2568 ( .a ({signal_4061, signal_2771}), .b ({signal_4105, signal_2815}), .c ({signal_4135, signal_2828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2569 ( .a ({signal_4056, signal_2766}), .b ({signal_4100, signal_2810}), .c ({signal_4136, signal_2333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2570 ( .a ({signal_4062, signal_2772}), .b ({signal_4099, signal_2809}), .c ({signal_4137, signal_2334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2571 ( .a ({signal_4102, signal_2812}), .b ({signal_4106, signal_2816}), .c ({signal_4138, signal_2335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2572 ( .a ({signal_4097, signal_2807}), .b ({signal_4104, signal_2814}), .c ({signal_4139, signal_2829}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2573 ( .a ({signal_4113, signal_2818}), .b ({signal_4160, signal_2298}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2574 ( .a ({signal_4114, signal_2819}), .b ({signal_4161, signal_2299}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2575 ( .a ({signal_4118, signal_2820}), .b ({signal_4162, signal_2303}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2576 ( .a ({signal_4120, signal_2821}), .b ({signal_4163, signal_2315}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2577 ( .a ({signal_4121, signal_2822}), .b ({signal_4164, signal_2316}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2578 ( .a ({signal_4125, signal_2823}), .b ({signal_4165, signal_2320}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2579 ( .a ({signal_4127, signal_2824}), .b ({signal_4166, signal_2323}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2580 ( .a ({signal_4128, signal_2825}), .b ({signal_4167, signal_2324}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2581 ( .a ({signal_4132, signal_2826}), .b ({signal_4168, signal_2328}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2582 ( .a ({signal_4134, signal_2827}), .b ({signal_4169, signal_2331}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2583 ( .a ({signal_4135, signal_2828}), .b ({signal_4170, signal_2332}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2584 ( .a ({signal_4139, signal_2829}), .b ({signal_4171, signal_2336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2585 ( .a ({signal_4126, signal_2322}), .b ({signal_4134, signal_2827}), .c ({signal_4172, signal_2830}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2586 ( .a ({signal_4127, signal_2824}), .b ({signal_4135, signal_2828}), .c ({signal_4173, signal_2831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2587 ( .a ({signal_4128, signal_2825}), .b ({signal_4136, signal_2333}), .c ({signal_4174, signal_2832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2588 ( .a ({signal_4131, signal_2327}), .b ({signal_4139, signal_2829}), .c ({signal_4175, signal_2833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2589 ( .a ({signal_4119, signal_2314}), .b ({signal_4127, signal_2824}), .c ({signal_4176, signal_2834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2590 ( .a ({signal_4120, signal_2821}), .b ({signal_4128, signal_2825}), .c ({signal_4177, signal_2835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2591 ( .a ({signal_4121, signal_2822}), .b ({signal_4129, signal_2325}), .c ({signal_4178, signal_2836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2592 ( .a ({signal_4124, signal_2319}), .b ({signal_4132, signal_2826}), .c ({signal_4179, signal_2837}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2593 ( .a ({signal_4085, signal_2795}), .b ({signal_4126, signal_2322}), .c ({signal_4180, signal_2838}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2594 ( .a ({signal_4074, signal_2784}), .b ({signal_4119, signal_2314}), .c ({signal_4181, signal_2839}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2595 ( .a ({signal_4112, signal_2305}), .b ({signal_4120, signal_2821}), .c ({signal_4182, signal_2840}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2596 ( .a ({signal_4113, signal_2818}), .b ({signal_4133, signal_2330}), .c ({signal_4183, signal_2841}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2597 ( .a ({signal_4113, signal_2818}), .b ({signal_4121, signal_2822}), .c ({signal_4184, signal_2842}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2598 ( .a ({signal_4114, signal_2819}), .b ({signal_4134, signal_2827}), .c ({signal_4185, signal_2843}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2599 ( .a ({signal_4114, signal_2819}), .b ({signal_4122, signal_2317}), .c ({signal_4186, signal_2844}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2600 ( .a ({signal_4115, signal_2300}), .b ({signal_4135, signal_2828}), .c ({signal_4187, signal_2845}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2601 ( .a ({signal_4117, signal_1843}), .b ({signal_4125, signal_2823}), .c ({signal_4188, signal_2846}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2602 ( .a ({signal_4118, signal_2820}), .b ({signal_4138, signal_2335}), .c ({signal_4189, signal_2847}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2603 ( .a ({signal_4096, signal_2806}), .b ({signal_4133, signal_2330}), .c ({signal_4190, signal_2848}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2604 ( .a ({signal_4107, signal_2817}), .b ({signal_4112, signal_2305}), .c ({signal_4191, signal_2849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2605 ( .a ({signal_4133, signal_2330}), .b ({signal_4137, signal_2334}), .c ({signal_4192, signal_2850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2606 ( .a ({signal_4133, signal_2330}), .b ({signal_4138, signal_2335}), .c ({signal_4193, signal_2851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2607 ( .a ({signal_4107, signal_2817}), .b ({signal_4133, signal_2330}), .c ({signal_4194, signal_2852}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2608 ( .a ({signal_4126, signal_2322}), .b ({signal_4130, signal_2326}), .c ({signal_4195, signal_2853}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2609 ( .a ({signal_4126, signal_2322}), .b ({signal_4131, signal_2327}), .c ({signal_4196, signal_2854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2610 ( .a ({signal_4096, signal_2806}), .b ({signal_4126, signal_2322}), .c ({signal_4197, signal_2855}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2611 ( .a ({signal_4119, signal_2314}), .b ({signal_4123, signal_2318}), .c ({signal_4198, signal_2856}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2612 ( .a ({signal_4119, signal_2314}), .b ({signal_4124, signal_2319}), .c ({signal_4199, signal_2857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2613 ( .a ({signal_4085, signal_2795}), .b ({signal_4119, signal_2314}), .c ({signal_4200, signal_2858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2614 ( .a ({signal_4112, signal_2305}), .b ({signal_4116, signal_1842}), .c ({signal_4201, signal_2859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2615 ( .a ({signal_4112, signal_2305}), .b ({signal_4117, signal_1843}), .c ({signal_4202, signal_2860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2616 ( .a ({signal_4074, signal_2784}), .b ({signal_4112, signal_2305}), .c ({signal_4203, signal_2861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2617 ( .a ({signal_4096, signal_2806}), .b ({signal_4191, signal_2849}), .c ({signal_4251, signal_2862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2618 ( .a ({signal_4119, signal_2314}), .b ({signal_4183, signal_2841}), .c ({signal_4252, signal_2863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2619 ( .a ({signal_4120, signal_2821}), .b ({signal_4185, signal_2843}), .c ({signal_4253, signal_2864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2620 ( .a ({signal_4121, signal_2822}), .b ({signal_4187, signal_2845}), .c ({signal_4254, signal_2865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2621 ( .a ({signal_4112, signal_2305}), .b ({signal_4176, signal_2834}), .c ({signal_4255, signal_2866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2622 ( .a ({signal_4113, signal_2818}), .b ({signal_4177, signal_2835}), .c ({signal_4256, signal_2867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2623 ( .a ({signal_4124, signal_2319}), .b ({signal_4189, signal_2847}), .c ({signal_4257, signal_2868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2624 ( .a ({signal_4114, signal_2819}), .b ({signal_4178, signal_2836}), .c ({signal_4258, signal_2869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2625 ( .a ({signal_4129, signal_2325}), .b ({signal_4192, signal_2850}), .c ({signal_4259, signal_2870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2626 ( .a ({signal_4130, signal_2326}), .b ({signal_4193, signal_2851}), .c ({signal_4260, signal_2871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2627 ( .a ({signal_4117, signal_1843}), .b ({signal_4179, signal_2837}), .c ({signal_4261, signal_2872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2628 ( .a ({signal_4074, signal_2784}), .b ({signal_4190, signal_2848}), .c ({signal_4262, signal_2873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2629 ( .a ({signal_4133, signal_2330}), .b ({signal_4182, signal_2840}), .c ({signal_4263, signal_2874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2630 ( .a ({signal_4134, signal_2827}), .b ({signal_4184, signal_2842}), .c ({signal_4264, signal_2875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2631 ( .a ({signal_4135, signal_2828}), .b ({signal_4186, signal_2844}), .c ({signal_4265, signal_2876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2632 ( .a ({signal_4122, signal_2317}), .b ({signal_4195, signal_2853}), .c ({signal_4266, signal_2877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2633 ( .a ({signal_4132, signal_2826}), .b ({signal_4194, signal_2852}), .c ({signal_4267, signal_2878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2634 ( .a ({signal_4139, signal_2829}), .b ({signal_4203, signal_2861}), .c ({signal_4268, signal_2879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2635 ( .a ({signal_4123, signal_2318}), .b ({signal_4196, signal_2854}), .c ({signal_4269, signal_2880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2636 ( .a ({signal_4138, signal_2335}), .b ({signal_4188, signal_2846}), .c ({signal_4270, signal_2881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2637 ( .a ({signal_4125, signal_2823}), .b ({signal_4197, signal_2855}), .c ({signal_4271, signal_2882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2638 ( .a ({signal_4118, signal_2820}), .b ({signal_4200, signal_2858}), .c ({signal_4272, signal_2883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2639 ( .a ({signal_4107, signal_2817}), .b ({signal_4181, signal_2839}), .c ({signal_4273, signal_2884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2640 ( .a ({signal_4126, signal_2322}), .b ({signal_4183, signal_2841}), .c ({signal_4274, signal_2885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2641 ( .a ({signal_4127, signal_2824}), .b ({signal_4185, signal_2843}), .c ({signal_4275, signal_2886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2642 ( .a ({signal_4128, signal_2825}), .b ({signal_4187, signal_2845}), .c ({signal_4276, signal_2887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2643 ( .a ({signal_4115, signal_2300}), .b ({signal_4198, signal_2856}), .c ({signal_4277, signal_2888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2644 ( .a ({signal_4136, signal_2333}), .b ({signal_4201, signal_2859}), .c ({signal_4278, signal_2889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2645 ( .a ({signal_4116, signal_1842}), .b ({signal_4199, signal_2857}), .c ({signal_4279, signal_2890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2646 ( .a ({signal_4137, signal_2334}), .b ({signal_4202, signal_2860}), .c ({signal_4280, signal_2891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2647 ( .a ({signal_4131, signal_2327}), .b ({signal_4189, signal_2847}), .c ({signal_4281, signal_2892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2648 ( .a ({signal_4190, signal_2848}), .b ({signal_4191, signal_2849}), .c ({signal_4282, signal_2893}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2649 ( .a ({signal_4282, signal_2893}), .b ({signal_4374, signal_1216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2650 ( .a ({signal_4268, signal_2879}), .b ({signal_4272, signal_2883}), .c ({signal_4375, signal_2894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2651 ( .a ({signal_4181, signal_2839}), .b ({signal_4251, signal_2862}), .c ({signal_4376, signal_2895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2652 ( .a ({signal_4172, signal_2830}), .b ({signal_4252, signal_2863}), .c ({signal_4377, signal_1870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2653 ( .a ({signal_4173, signal_2831}), .b ({signal_4253, signal_2864}), .c ({signal_4378, signal_2896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2654 ( .a ({signal_4174, signal_2832}), .b ({signal_4254, signal_2865}), .c ({signal_4379, signal_2897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2655 ( .a ({signal_4122, signal_2317}), .b ({signal_4278, signal_2889}), .c ({signal_4380, signal_2898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2656 ( .a ({signal_4123, signal_2318}), .b ({signal_4280, signal_2891}), .c ({signal_4381, signal_2899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2657 ( .a ({signal_4172, signal_2830}), .b ({signal_4255, signal_2866}), .c ({signal_4382, signal_1846}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2658 ( .a ({signal_4173, signal_2831}), .b ({signal_4256, signal_2867}), .c ({signal_4383, signal_2900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2659 ( .a ({signal_4175, signal_2833}), .b ({signal_4257, signal_2868}), .c ({signal_4384, signal_1875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2660 ( .a ({signal_4174, signal_2832}), .b ({signal_4258, signal_2869}), .c ({signal_4385, signal_2901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2661 ( .a ({signal_4115, signal_2300}), .b ({signal_4266, signal_2877}), .c ({signal_4386, signal_2902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2662 ( .a ({signal_4116, signal_1842}), .b ({signal_4269, signal_2880}), .c ({signal_4387, signal_2903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2663 ( .a ({signal_4175, signal_2833}), .b ({signal_4261, signal_2872}), .c ({signal_4388, signal_1851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2664 ( .a ({signal_4118, signal_2820}), .b ({signal_4271, signal_2882}), .c ({signal_4389, signal_2904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2665 ( .a ({signal_4180, signal_2838}), .b ({signal_4262, signal_2873}), .c ({signal_4390, signal_2905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2666 ( .a ({signal_4176, signal_2834}), .b ({signal_4263, signal_2874}), .c ({signal_4391, signal_1854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2667 ( .a ({signal_4177, signal_2835}), .b ({signal_4264, signal_2875}), .c ({signal_4392, signal_2906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2668 ( .a ({signal_4178, signal_2836}), .b ({signal_4265, signal_2876}), .c ({signal_4393, signal_2907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2669 ( .a ({signal_4136, signal_2333}), .b ({signal_4277, signal_2888}), .c ({signal_4394, signal_2908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2670 ( .a ({signal_4125, signal_2823}), .b ({signal_4268, signal_2879}), .c ({signal_4395, signal_2909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2671 ( .a ({signal_4137, signal_2334}), .b ({signal_4279, signal_2890}), .c ({signal_4396, signal_2910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2672 ( .a ({signal_4179, signal_2837}), .b ({signal_4270, signal_2881}), .c ({signal_4397, signal_1859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2673 ( .a ({signal_4139, signal_2829}), .b ({signal_4272, signal_2883}), .c ({signal_4398, signal_2911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2674 ( .a ({signal_4180, signal_2838}), .b ({signal_4273, signal_2884}), .c ({signal_4399, signal_2912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2675 ( .a ({signal_4182, signal_2840}), .b ({signal_4274, signal_2885}), .c ({signal_4400, signal_1862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2676 ( .a ({signal_4184, signal_2842}), .b ({signal_4275, signal_2886}), .c ({signal_4401, signal_2913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2677 ( .a ({signal_4186, signal_2844}), .b ({signal_4276, signal_2887}), .c ({signal_4402, signal_2914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2678 ( .a ({signal_4129, signal_2325}), .b ({signal_4278, signal_2889}), .c ({signal_4403, signal_2915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2679 ( .a ({signal_4130, signal_2326}), .b ({signal_4280, signal_2891}), .c ({signal_4404, signal_2916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2680 ( .a ({signal_4188, signal_2846}), .b ({signal_4281, signal_2892}), .c ({signal_4405, signal_1867}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2681 ( .a ({signal_4375, signal_2894}), .b ({signal_4537, signal_1153}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2682 ( .a ({signal_4376, signal_2895}), .b ({signal_4538, signal_1869}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2683 ( .a ({signal_4378, signal_2896}), .b ({signal_4539, signal_1871}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2684 ( .a ({signal_4379, signal_2897}), .b ({signal_4540, signal_1872}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2685 ( .a ({signal_4383, signal_2900}), .b ({signal_4541, signal_1847}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2686 ( .a ({signal_4385, signal_2901}), .b ({signal_4542, signal_1848}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2687 ( .a ({signal_4390, signal_2905}), .b ({signal_4543, signal_1853}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2688 ( .a ({signal_4392, signal_2906}), .b ({signal_4544, signal_1855}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2689 ( .a ({signal_4393, signal_2907}), .b ({signal_4545, signal_1856}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2690 ( .a ({signal_4399, signal_2912}), .b ({signal_4546, signal_1861}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2691 ( .a ({signal_4401, signal_2913}), .b ({signal_4547, signal_1863}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2692 ( .a ({signal_4402, signal_2914}), .b ({signal_4548, signal_1864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2693 ( .a ({signal_4259, signal_2870}), .b ({signal_4380, signal_2898}), .c ({signal_4549, signal_1873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2694 ( .a ({signal_4260, signal_2871}), .b ({signal_4381, signal_2899}), .c ({signal_4550, signal_1874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2695 ( .a ({signal_4259, signal_2870}), .b ({signal_4386, signal_2902}), .c ({signal_4551, signal_1849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2696 ( .a ({signal_4260, signal_2871}), .b ({signal_4387, signal_2903}), .c ({signal_4552, signal_1850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2697 ( .a ({signal_4267, signal_2878}), .b ({signal_4389, signal_2904}), .c ({signal_4553, signal_2917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2698 ( .a ({signal_4266, signal_2877}), .b ({signal_4394, signal_2908}), .c ({signal_4554, signal_1857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2699 ( .a ({signal_4267, signal_2878}), .b ({signal_4395, signal_2909}), .c ({signal_4555, signal_2918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2700 ( .a ({signal_4269, signal_2880}), .b ({signal_4396, signal_2910}), .c ({signal_4556, signal_1858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2701 ( .a ({signal_4271, signal_2882}), .b ({signal_4398, signal_2911}), .c ({signal_4557, signal_2919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2702 ( .a ({signal_4277, signal_2888}), .b ({signal_4403, signal_2915}), .c ({signal_4558, signal_1865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2703 ( .a ({signal_4279, signal_2890}), .b ({signal_4404, signal_2916}), .c ({signal_4559, signal_1866}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2704 ( .a ({signal_4553, signal_2917}), .b ({signal_4702, signal_1852}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2705 ( .a ({signal_4555, signal_2918}), .b ({signal_4703, signal_1876}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2706 ( .a ({signal_4557, signal_2919}), .b ({signal_4704, signal_1860}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_159 ( .D ({signal_4830, signal_414}), .clk (signal_5060), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_162 ( .D ({signal_4911, signal_416}), .clk (signal_5060), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_165 ( .D ({signal_4706, signal_418}), .clk (signal_5060), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_168 ( .D ({signal_4832, signal_420}), .clk (signal_5060), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_171 ( .D ({signal_4834, signal_422}), .clk (signal_5060), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_174 ( .D ({signal_4836, signal_424}), .clk (signal_5060), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_177 ( .D ({signal_4838, signal_426}), .clk (signal_5060), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_180 ( .D ({signal_4708, signal_428}), .clk (signal_5060), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_183 ( .D ({signal_4840, signal_430}), .clk (signal_5060), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_186 ( .D ({signal_4913, signal_432}), .clk (signal_5060), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_189 ( .D ({signal_4710, signal_434}), .clk (signal_5060), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_192 ( .D ({signal_4842, signal_436}), .clk (signal_5060), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_195 ( .D ({signal_4844, signal_438}), .clk (signal_5060), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_198 ( .D ({signal_4846, signal_440}), .clk (signal_5060), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_201 ( .D ({signal_4848, signal_442}), .clk (signal_5060), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_204 ( .D ({signal_4712, signal_444}), .clk (signal_5060), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_207 ( .D ({signal_4850, signal_446}), .clk (signal_5060), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_210 ( .D ({signal_4915, signal_448}), .clk (signal_5060), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_213 ( .D ({signal_4714, signal_450}), .clk (signal_5060), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_216 ( .D ({signal_4852, signal_452}), .clk (signal_5060), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_219 ( .D ({signal_4854, signal_454}), .clk (signal_5060), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_222 ( .D ({signal_4856, signal_456}), .clk (signal_5060), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_225 ( .D ({signal_4858, signal_458}), .clk (signal_5060), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_228 ( .D ({signal_4716, signal_460}), .clk (signal_5060), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_231 ( .D ({signal_4860, signal_462}), .clk (signal_5060), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_234 ( .D ({signal_4917, signal_464}), .clk (signal_5060), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_237 ( .D ({signal_4718, signal_466}), .clk (signal_5060), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_240 ( .D ({signal_4862, signal_468}), .clk (signal_5060), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_243 ( .D ({signal_4864, signal_470}), .clk (signal_5060), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_246 ( .D ({signal_4866, signal_472}), .clk (signal_5060), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_249 ( .D ({signal_4868, signal_474}), .clk (signal_5060), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_252 ( .D ({signal_4720, signal_476}), .clk (signal_5060), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_255 ( .D ({signal_3433, signal_478}), .clk (signal_5060), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_258 ( .D ({signal_3435, signal_480}), .clk (signal_5060), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_261 ( .D ({signal_3437, signal_482}), .clk (signal_5060), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_264 ( .D ({signal_3439, signal_484}), .clk (signal_5060), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_267 ( .D ({signal_3441, signal_486}), .clk (signal_5060), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_270 ( .D ({signal_3443, signal_488}), .clk (signal_5060), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_273 ( .D ({signal_3445, signal_490}), .clk (signal_5060), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_276 ( .D ({signal_3447, signal_492}), .clk (signal_5060), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_279 ( .D ({signal_3449, signal_494}), .clk (signal_5060), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_282 ( .D ({signal_3451, signal_496}), .clk (signal_5060), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_285 ( .D ({signal_3453, signal_498}), .clk (signal_5060), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_288 ( .D ({signal_3455, signal_500}), .clk (signal_5060), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_291 ( .D ({signal_3457, signal_502}), .clk (signal_5060), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_294 ( .D ({signal_3459, signal_504}), .clk (signal_5060), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_297 ( .D ({signal_3461, signal_506}), .clk (signal_5060), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_300 ( .D ({signal_3463, signal_508}), .clk (signal_5060), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_303 ( .D ({signal_3465, signal_510}), .clk (signal_5060), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_306 ( .D ({signal_3467, signal_512}), .clk (signal_5060), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_309 ( .D ({signal_3469, signal_514}), .clk (signal_5060), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_312 ( .D ({signal_3471, signal_516}), .clk (signal_5060), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_315 ( .D ({signal_3473, signal_518}), .clk (signal_5060), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_318 ( .D ({signal_3475, signal_520}), .clk (signal_5060), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_321 ( .D ({signal_3477, signal_522}), .clk (signal_5060), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_324 ( .D ({signal_3479, signal_524}), .clk (signal_5060), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_327 ( .D ({signal_3481, signal_526}), .clk (signal_5060), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_330 ( .D ({signal_3483, signal_528}), .clk (signal_5060), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_333 ( .D ({signal_3485, signal_530}), .clk (signal_5060), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_336 ( .D ({signal_3487, signal_532}), .clk (signal_5060), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_339 ( .D ({signal_3489, signal_534}), .clk (signal_5060), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_342 ( .D ({signal_3491, signal_536}), .clk (signal_5060), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_345 ( .D ({signal_3493, signal_538}), .clk (signal_5060), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_348 ( .D ({signal_3495, signal_540}), .clk (signal_5060), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_351 ( .D ({signal_3497, signal_542}), .clk (signal_5060), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_354 ( .D ({signal_3499, signal_544}), .clk (signal_5060), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_357 ( .D ({signal_3501, signal_546}), .clk (signal_5060), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_360 ( .D ({signal_3503, signal_548}), .clk (signal_5060), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_363 ( .D ({signal_3505, signal_550}), .clk (signal_5060), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_366 ( .D ({signal_3507, signal_552}), .clk (signal_5060), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_369 ( .D ({signal_3509, signal_554}), .clk (signal_5060), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_372 ( .D ({signal_3511, signal_556}), .clk (signal_5060), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_375 ( .D ({signal_3513, signal_558}), .clk (signal_5060), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_378 ( .D ({signal_3515, signal_560}), .clk (signal_5060), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_381 ( .D ({signal_3517, signal_562}), .clk (signal_5060), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_384 ( .D ({signal_3519, signal_564}), .clk (signal_5060), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_387 ( .D ({signal_3521, signal_566}), .clk (signal_5060), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_390 ( .D ({signal_3523, signal_568}), .clk (signal_5060), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_393 ( .D ({signal_3525, signal_570}), .clk (signal_5060), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_396 ( .D ({signal_3527, signal_572}), .clk (signal_5060), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_399 ( .D ({signal_3529, signal_574}), .clk (signal_5060), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_402 ( .D ({signal_3531, signal_576}), .clk (signal_5060), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_405 ( .D ({signal_3533, signal_578}), .clk (signal_5060), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_408 ( .D ({signal_3535, signal_580}), .clk (signal_5060), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_411 ( .D ({signal_3537, signal_582}), .clk (signal_5060), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_414 ( .D ({signal_3539, signal_584}), .clk (signal_5060), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_417 ( .D ({signal_3541, signal_586}), .clk (signal_5060), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_420 ( .D ({signal_3543, signal_588}), .clk (signal_5060), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_423 ( .D ({signal_3545, signal_590}), .clk (signal_5060), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_426 ( .D ({signal_3547, signal_592}), .clk (signal_5060), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_429 ( .D ({signal_3549, signal_594}), .clk (signal_5060), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_432 ( .D ({signal_3551, signal_596}), .clk (signal_5060), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_435 ( .D ({signal_3553, signal_598}), .clk (signal_5060), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_438 ( .D ({signal_3555, signal_600}), .clk (signal_5060), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_441 ( .D ({signal_3557, signal_602}), .clk (signal_5060), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_444 ( .D ({signal_3559, signal_604}), .clk (signal_5060), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_447 ( .D ({signal_3561, signal_606}), .clk (signal_5060), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_450 ( .D ({signal_3563, signal_608}), .clk (signal_5060), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_453 ( .D ({signal_3565, signal_610}), .clk (signal_5060), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_456 ( .D ({signal_3567, signal_612}), .clk (signal_5060), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_459 ( .D ({signal_3569, signal_614}), .clk (signal_5060), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_462 ( .D ({signal_3571, signal_616}), .clk (signal_5060), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_465 ( .D ({signal_3573, signal_618}), .clk (signal_5060), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_468 ( .D ({signal_3575, signal_620}), .clk (signal_5060), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_471 ( .D ({signal_3577, signal_622}), .clk (signal_5060), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_474 ( .D ({signal_3579, signal_624}), .clk (signal_5060), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_477 ( .D ({signal_3581, signal_626}), .clk (signal_5060), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_480 ( .D ({signal_3583, signal_628}), .clk (signal_5060), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_483 ( .D ({signal_3585, signal_630}), .clk (signal_5060), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_486 ( .D ({signal_3587, signal_632}), .clk (signal_5060), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_489 ( .D ({signal_3589, signal_634}), .clk (signal_5060), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_492 ( .D ({signal_3591, signal_636}), .clk (signal_5060), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_495 ( .D ({signal_3593, signal_638}), .clk (signal_5060), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_498 ( .D ({signal_3595, signal_640}), .clk (signal_5060), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_501 ( .D ({signal_3597, signal_642}), .clk (signal_5060), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_504 ( .D ({signal_3599, signal_644}), .clk (signal_5060), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_507 ( .D ({signal_3601, signal_646}), .clk (signal_5060), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_510 ( .D ({signal_3603, signal_648}), .clk (signal_5060), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_513 ( .D ({signal_3605, signal_650}), .clk (signal_5060), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_516 ( .D ({signal_3607, signal_652}), .clk (signal_5060), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_519 ( .D ({signal_3609, signal_654}), .clk (signal_5060), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_522 ( .D ({signal_3611, signal_656}), .clk (signal_5060), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_525 ( .D ({signal_3613, signal_658}), .clk (signal_5060), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_528 ( .D ({signal_3615, signal_660}), .clk (signal_5060), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_531 ( .D ({signal_3617, signal_662}), .clk (signal_5060), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_534 ( .D ({signal_3619, signal_664}), .clk (signal_5060), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_537 ( .D ({signal_3621, signal_666}), .clk (signal_5060), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_540 ( .D ({signal_3623, signal_668}), .clk (signal_5060), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1368 ( .D ({signal_4746, signal_1227}), .clk (signal_5060), .Q ({signal_2921, signal_1793}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1371 ( .D ({signal_4874, signal_1229}), .clk (signal_5060), .Q ({signal_3038, signal_1792}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1374 ( .D ({signal_4748, signal_1231}), .clk (signal_5060), .Q ({signal_3071, signal_1791}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1377 ( .D ({signal_4750, signal_1233}), .clk (signal_5060), .Q ({signal_3104, signal_1790}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1380 ( .D ({signal_4752, signal_1235}), .clk (signal_5060), .Q ({signal_3137, signal_1789}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1383 ( .D ({signal_4876, signal_1237}), .clk (signal_5060), .Q ({signal_3170, signal_1788}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1386 ( .D ({signal_4878, signal_1239}), .clk (signal_5060), .Q ({signal_3203, signal_1787}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1389 ( .D ({signal_4754, signal_1241}), .clk (signal_5060), .Q ({signal_3236, signal_1786}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1392 ( .D ({signal_4756, signal_1243}), .clk (signal_5060), .Q ({signal_3269, signal_1801}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1395 ( .D ({signal_4880, signal_1245}), .clk (signal_5060), .Q ({signal_3302, signal_1800}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1398 ( .D ({signal_4758, signal_1247}), .clk (signal_5060), .Q ({signal_2954, signal_1799}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1401 ( .D ({signal_4760, signal_1249}), .clk (signal_5060), .Q ({signal_2987, signal_1798}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1404 ( .D ({signal_4762, signal_1251}), .clk (signal_5060), .Q ({signal_3014, signal_1797}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1407 ( .D ({signal_4882, signal_1253}), .clk (signal_5060), .Q ({signal_3017, signal_1796}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1410 ( .D ({signal_4884, signal_1255}), .clk (signal_5060), .Q ({signal_3020, signal_1795}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1413 ( .D ({signal_4764, signal_1257}), .clk (signal_5060), .Q ({signal_3023, signal_1794}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1416 ( .D ({signal_4766, signal_1259}), .clk (signal_5060), .Q ({signal_3026, signal_1809}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1419 ( .D ({signal_4886, signal_1261}), .clk (signal_5060), .Q ({signal_3029, signal_1808}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1422 ( .D ({signal_4768, signal_1263}), .clk (signal_5060), .Q ({signal_3032, signal_1807}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1425 ( .D ({signal_4770, signal_1265}), .clk (signal_5060), .Q ({signal_3035, signal_1806}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1428 ( .D ({signal_4772, signal_1267}), .clk (signal_5060), .Q ({signal_3041, signal_1805}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1431 ( .D ({signal_4888, signal_1269}), .clk (signal_5060), .Q ({signal_3044, signal_1804}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1434 ( .D ({signal_4890, signal_1271}), .clk (signal_5060), .Q ({signal_3047, signal_1803}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1437 ( .D ({signal_4774, signal_1273}), .clk (signal_5060), .Q ({signal_3050, signal_1802}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1440 ( .D ({signal_4892, signal_1275}), .clk (signal_5060), .Q ({signal_3053, signal_1785}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1443 ( .D ({signal_4919, signal_1277}), .clk (signal_5060), .Q ({signal_3056, signal_1784}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1446 ( .D ({signal_4894, signal_1279}), .clk (signal_5060), .Q ({signal_3059, signal_1783}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1449 ( .D ({signal_4896, signal_1281}), .clk (signal_5060), .Q ({signal_3062, signal_1782}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1452 ( .D ({signal_4898, signal_1283}), .clk (signal_5060), .Q ({signal_3065, signal_1781}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1455 ( .D ({signal_4921, signal_1285}), .clk (signal_5060), .Q ({signal_3068, signal_1780}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1458 ( .D ({signal_4923, signal_1287}), .clk (signal_5060), .Q ({signal_3074, signal_1779}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1461 ( .D ({signal_4900, signal_1289}), .clk (signal_5060), .Q ({signal_3077, signal_1778}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1464 ( .D ({signal_4590, signal_1291}), .clk (signal_5060), .Q ({signal_3080, signal_2133}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1467 ( .D ({signal_4776, signal_1293}), .clk (signal_5060), .Q ({signal_3083, signal_2132}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1470 ( .D ({signal_4592, signal_1295}), .clk (signal_5060), .Q ({signal_3086, signal_2131}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1473 ( .D ({signal_4594, signal_1297}), .clk (signal_5060), .Q ({signal_3089, signal_2130}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1476 ( .D ({signal_4596, signal_1299}), .clk (signal_5060), .Q ({signal_3092, signal_2129}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1479 ( .D ({signal_4778, signal_1301}), .clk (signal_5060), .Q ({signal_3095, signal_2128}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1482 ( .D ({signal_4780, signal_1303}), .clk (signal_5060), .Q ({signal_3098, signal_2127}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1485 ( .D ({signal_4598, signal_1305}), .clk (signal_5060), .Q ({signal_3101, signal_2126}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1488 ( .D ({signal_4600, signal_1307}), .clk (signal_5060), .Q ({signal_3107, signal_2125}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1491 ( .D ({signal_4782, signal_1309}), .clk (signal_5060), .Q ({signal_3110, signal_2124}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1494 ( .D ({signal_4602, signal_1311}), .clk (signal_5060), .Q ({signal_3113, signal_2123}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1497 ( .D ({signal_4604, signal_1313}), .clk (signal_5060), .Q ({signal_3116, signal_2122}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1500 ( .D ({signal_4606, signal_1315}), .clk (signal_5060), .Q ({signal_3119, signal_2121}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1503 ( .D ({signal_4784, signal_1317}), .clk (signal_5060), .Q ({signal_3122, signal_2120}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1506 ( .D ({signal_4786, signal_1319}), .clk (signal_5060), .Q ({signal_3125, signal_2119}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1509 ( .D ({signal_4608, signal_1321}), .clk (signal_5060), .Q ({signal_3128, signal_2118}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1512 ( .D ({signal_4610, signal_1323}), .clk (signal_5060), .Q ({signal_3131, signal_2117}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1515 ( .D ({signal_4788, signal_1325}), .clk (signal_5060), .Q ({signal_3134, signal_2116}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1518 ( .D ({signal_4612, signal_1327}), .clk (signal_5060), .Q ({signal_3140, signal_2115}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1521 ( .D ({signal_4614, signal_1329}), .clk (signal_5060), .Q ({signal_3143, signal_2114}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1524 ( .D ({signal_4616, signal_1331}), .clk (signal_5060), .Q ({signal_3146, signal_2113}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1527 ( .D ({signal_4790, signal_1333}), .clk (signal_5060), .Q ({signal_3149, signal_2112}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1530 ( .D ({signal_4792, signal_1335}), .clk (signal_5060), .Q ({signal_3152, signal_2111}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1533 ( .D ({signal_4618, signal_1337}), .clk (signal_5060), .Q ({signal_3155, signal_2110}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1536 ( .D ({signal_4794, signal_1339}), .clk (signal_5060), .Q ({signal_3158, signal_2109}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1539 ( .D ({signal_4902, signal_1341}), .clk (signal_5060), .Q ({signal_3161, signal_2108}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1542 ( .D ({signal_4796, signal_1343}), .clk (signal_5060), .Q ({signal_3164, signal_2107}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1545 ( .D ({signal_4798, signal_1345}), .clk (signal_5060), .Q ({signal_3167, signal_2106}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1548 ( .D ({signal_4800, signal_1347}), .clk (signal_5060), .Q ({signal_3173, signal_2105}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1551 ( .D ({signal_4904, signal_1349}), .clk (signal_5060), .Q ({signal_3176, signal_2104}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1554 ( .D ({signal_4906, signal_1351}), .clk (signal_5060), .Q ({signal_3179, signal_2103}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1557 ( .D ({signal_4802, signal_1353}), .clk (signal_5060), .Q ({signal_3182, signal_2102}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1560 ( .D ({signal_4416, signal_1355}), .clk (signal_5060), .Q ({signal_3185, signal_2101}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1563 ( .D ({signal_4620, signal_1357}), .clk (signal_5060), .Q ({signal_3188, signal_2100}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1566 ( .D ({signal_4418, signal_1359}), .clk (signal_5060), .Q ({signal_3191, signal_2099}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1569 ( .D ({signal_4420, signal_1361}), .clk (signal_5060), .Q ({signal_3194, signal_2098}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1572 ( .D ({signal_4422, signal_1363}), .clk (signal_5060), .Q ({signal_3197, signal_2097}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1575 ( .D ({signal_4622, signal_1365}), .clk (signal_5060), .Q ({signal_3200, signal_2096}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1578 ( .D ({signal_4624, signal_1367}), .clk (signal_5060), .Q ({signal_3206, signal_2095}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1581 ( .D ({signal_4424, signal_1369}), .clk (signal_5060), .Q ({signal_3209, signal_2094}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1584 ( .D ({signal_4426, signal_1371}), .clk (signal_5060), .Q ({signal_3212, signal_2093}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1587 ( .D ({signal_4626, signal_1373}), .clk (signal_5060), .Q ({signal_3215, signal_2092}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1590 ( .D ({signal_4428, signal_1375}), .clk (signal_5060), .Q ({signal_3218, signal_2091}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1593 ( .D ({signal_4430, signal_1377}), .clk (signal_5060), .Q ({signal_3221, signal_2090}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1596 ( .D ({signal_4432, signal_1379}), .clk (signal_5060), .Q ({signal_3224, signal_2089}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1599 ( .D ({signal_4628, signal_1381}), .clk (signal_5060), .Q ({signal_3227, signal_2088}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1602 ( .D ({signal_4630, signal_1383}), .clk (signal_5060), .Q ({signal_3230, signal_2087}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1605 ( .D ({signal_4434, signal_1385}), .clk (signal_5060), .Q ({signal_3233, signal_2086}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1608 ( .D ({signal_4436, signal_1387}), .clk (signal_5060), .Q ({signal_3239, signal_2085}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1611 ( .D ({signal_4632, signal_1389}), .clk (signal_5060), .Q ({signal_3242, signal_2084}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1614 ( .D ({signal_4438, signal_1391}), .clk (signal_5060), .Q ({signal_3245, signal_2083}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1617 ( .D ({signal_4440, signal_1393}), .clk (signal_5060), .Q ({signal_3248, signal_2082}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1620 ( .D ({signal_4442, signal_1395}), .clk (signal_5060), .Q ({signal_3251, signal_2081}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1623 ( .D ({signal_4634, signal_1397}), .clk (signal_5060), .Q ({signal_3254, signal_2080}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1626 ( .D ({signal_4636, signal_1399}), .clk (signal_5060), .Q ({signal_3257, signal_2079}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1629 ( .D ({signal_4444, signal_1401}), .clk (signal_5060), .Q ({signal_3260, signal_2078}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1632 ( .D ({signal_4638, signal_1403}), .clk (signal_5060), .Q ({signal_3263, signal_2077}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1635 ( .D ({signal_4804, signal_1405}), .clk (signal_5060), .Q ({signal_3266, signal_2076}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1638 ( .D ({signal_4640, signal_1407}), .clk (signal_5060), .Q ({signal_3272, signal_2075}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1641 ( .D ({signal_4642, signal_1409}), .clk (signal_5060), .Q ({signal_3275, signal_2074}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1644 ( .D ({signal_4644, signal_1411}), .clk (signal_5060), .Q ({signal_3278, signal_2073}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1647 ( .D ({signal_4806, signal_1413}), .clk (signal_5060), .Q ({signal_3281, signal_2072}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1650 ( .D ({signal_4808, signal_1415}), .clk (signal_5060), .Q ({signal_3284, signal_2071}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1653 ( .D ({signal_4646, signal_1417}), .clk (signal_5060), .Q ({signal_3287, signal_2070}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1656 ( .D ({signal_4284, signal_1419}), .clk (signal_5060), .Q ({signal_3290, signal_2069}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1659 ( .D ({signal_4446, signal_1421}), .clk (signal_5060), .Q ({signal_3293, signal_2068}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1662 ( .D ({signal_4286, signal_1423}), .clk (signal_5060), .Q ({signal_3296, signal_2067}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1665 ( .D ({signal_4288, signal_1425}), .clk (signal_5060), .Q ({signal_3299, signal_2066}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1668 ( .D ({signal_4290, signal_1427}), .clk (signal_5060), .Q ({signal_2924, signal_2065}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1671 ( .D ({signal_4448, signal_1429}), .clk (signal_5060), .Q ({signal_2927, signal_2064}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1674 ( .D ({signal_4450, signal_1431}), .clk (signal_5060), .Q ({signal_2930, signal_2063}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1677 ( .D ({signal_4292, signal_1433}), .clk (signal_5060), .Q ({signal_2933, signal_2062}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1680 ( .D ({signal_4294, signal_1435}), .clk (signal_5060), .Q ({signal_2936, signal_2061}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1683 ( .D ({signal_4452, signal_1437}), .clk (signal_5060), .Q ({signal_2939, signal_2060}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1686 ( .D ({signal_4296, signal_1439}), .clk (signal_5060), .Q ({signal_2942, signal_2059}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1689 ( .D ({signal_4298, signal_1441}), .clk (signal_5060), .Q ({signal_2945, signal_2058}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1692 ( .D ({signal_4300, signal_1443}), .clk (signal_5060), .Q ({signal_2948, signal_2057}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1695 ( .D ({signal_4454, signal_1445}), .clk (signal_5060), .Q ({signal_2951, signal_2056}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1698 ( .D ({signal_4456, signal_1447}), .clk (signal_5060), .Q ({signal_2957, signal_2055}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1701 ( .D ({signal_4302, signal_1449}), .clk (signal_5060), .Q ({signal_2960, signal_2054}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1704 ( .D ({signal_4304, signal_1451}), .clk (signal_5060), .Q ({signal_2963, signal_2053}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1707 ( .D ({signal_4458, signal_1453}), .clk (signal_5060), .Q ({signal_2966, signal_2052}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1710 ( .D ({signal_4306, signal_1455}), .clk (signal_5060), .Q ({signal_2969, signal_2051}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1713 ( .D ({signal_4308, signal_1457}), .clk (signal_5060), .Q ({signal_2972, signal_2050}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1716 ( .D ({signal_4310, signal_1459}), .clk (signal_5060), .Q ({signal_2975, signal_2049}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1719 ( .D ({signal_4460, signal_1461}), .clk (signal_5060), .Q ({signal_2978, signal_2048}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1722 ( .D ({signal_4462, signal_1463}), .clk (signal_5060), .Q ({signal_2981, signal_2047}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1725 ( .D ({signal_4312, signal_1465}), .clk (signal_5060), .Q ({signal_2984, signal_2046}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1728 ( .D ({signal_4464, signal_1467}), .clk (signal_5060), .Q ({signal_2990, signal_2045}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1731 ( .D ({signal_4648, signal_1469}), .clk (signal_5060), .Q ({signal_2993, signal_2044}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1734 ( .D ({signal_4466, signal_1471}), .clk (signal_5060), .Q ({signal_2996, signal_2043}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1737 ( .D ({signal_4468, signal_1473}), .clk (signal_5060), .Q ({signal_2999, signal_2042}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1740 ( .D ({signal_4470, signal_1475}), .clk (signal_5060), .Q ({signal_3002, signal_2041}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1743 ( .D ({signal_4650, signal_1477}), .clk (signal_5060), .Q ({signal_3005, signal_2040}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1746 ( .D ({signal_4652, signal_1479}), .clk (signal_5060), .Q ({signal_3008, signal_2039}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1749 ( .D ({signal_4472, signal_1481}), .clk (signal_5060), .Q ({signal_3011, signal_2038}) ) ;
    DFF_X1 cell_2035 ( .D (signal_1502), .CK (signal_5060), .Q (signal_2273), .QN () ) ;
    DFF_X1 cell_2037 ( .D (signal_1501), .CK (signal_5060), .Q (signal_2272), .QN () ) ;
    DFF_X1 cell_2039 ( .D (signal_1499), .CK (signal_5060), .Q (signal_2271), .QN () ) ;
    DFF_X1 cell_2041 ( .D (signal_1498), .CK (signal_5060), .Q (signal_2270), .QN () ) ;
    DFF_X1 cell_2056 ( .D (signal_1520), .CK (signal_5060), .Q (signal_2276), .QN () ) ;
    DFF_X1 cell_2058 ( .D (signal_1519), .CK (signal_5060), .Q (signal_2275), .QN () ) ;
    DFF_X1 cell_2060 ( .D (signal_1518), .CK (signal_5060), .Q (signal_2274), .QN () ) ;
endmodule
