/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [11:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    wire Q0 ;
    wire Q1 ;
    wire T0 ;
    wire Q2 ;
    wire T1 ;
    wire Q4 ;
    wire T2 ;
    wire L0 ;
    wire Q6 ;
    wire L1 ;
    wire Q7 ;
    wire T3 ;
    wire L2 ;
    wire L2_T1 ;
    wire L3 ;
    wire n2 ;
    wire [2:1] XX ;
    wire [3:0] YY ;
    wire new_AGEMA_signal_39 ;
    wire new_AGEMA_signal_40 ;
    wire new_AGEMA_signal_43 ;
    wire new_AGEMA_signal_44 ;
    wire new_AGEMA_signal_47 ;
    wire new_AGEMA_signal_48 ;
    wire new_AGEMA_signal_51 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_53 ;
    wire new_AGEMA_signal_54 ;
    wire new_AGEMA_signal_55 ;
    wire new_AGEMA_signal_56 ;
    wire new_AGEMA_signal_57 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_61 ;
    wire new_AGEMA_signal_62 ;
    wire new_AGEMA_signal_63 ;
    wire new_AGEMA_signal_64 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_109 ;
    wire new_AGEMA_signal_110 ;
    wire new_AGEMA_signal_111 ;
    wire new_AGEMA_signal_112 ;
    wire new_AGEMA_signal_113 ;
    wire new_AGEMA_signal_114 ;
    wire new_AGEMA_signal_115 ;
    wire new_AGEMA_signal_116 ;
    wire new_AGEMA_signal_117 ;
    wire new_AGEMA_signal_118 ;
    wire new_AGEMA_signal_119 ;
    wire new_AGEMA_signal_120 ;
    wire new_AGEMA_signal_121 ;
    wire new_AGEMA_signal_122 ;
    wire new_AGEMA_signal_123 ;
    wire new_AGEMA_signal_124 ;
    wire new_AGEMA_signal_125 ;
    wire new_AGEMA_signal_126 ;
    wire new_AGEMA_signal_127 ;
    wire new_AGEMA_signal_128 ;
    wire new_AGEMA_signal_129 ;
    wire new_AGEMA_signal_130 ;
    wire new_AGEMA_signal_131 ;
    wire new_AGEMA_signal_132 ;
    wire new_AGEMA_signal_133 ;
    wire new_AGEMA_signal_134 ;
    wire new_AGEMA_signal_135 ;
    wire new_AGEMA_signal_136 ;
    wire new_AGEMA_signal_137 ;
    wire new_AGEMA_signal_138 ;
    wire new_AGEMA_signal_139 ;
    wire new_AGEMA_signal_140 ;
    wire new_AGEMA_signal_141 ;
    wire new_AGEMA_signal_142 ;
    wire new_AGEMA_signal_143 ;
    wire new_AGEMA_signal_144 ;
    wire new_AGEMA_signal_145 ;
    wire new_AGEMA_signal_146 ;
    wire new_AGEMA_signal_147 ;
    wire new_AGEMA_signal_148 ;
    wire new_AGEMA_signal_149 ;
    wire new_AGEMA_signal_150 ;
    wire new_AGEMA_signal_151 ;
    wire new_AGEMA_signal_152 ;
    wire new_AGEMA_signal_153 ;
    wire new_AGEMA_signal_154 ;
    wire new_AGEMA_signal_155 ;
    wire new_AGEMA_signal_156 ;
    wire new_AGEMA_signal_157 ;
    wire new_AGEMA_signal_158 ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_161 ;
    wire new_AGEMA_signal_162 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_166 ;
    wire new_AGEMA_signal_167 ;
    wire new_AGEMA_signal_168 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_171 ;
    wire new_AGEMA_signal_172 ;
    wire new_AGEMA_signal_173 ;
    wire new_AGEMA_signal_174 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) U5 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR_i1_U1 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s2[3], X_s1[3], X_s0[3]}), .c ({new_AGEMA_signal_44, new_AGEMA_signal_43, XX[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR_i2_U1 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_48, new_AGEMA_signal_47, XX[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR0_U1 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_48, new_AGEMA_signal_47, XX[2]}), .c ({new_AGEMA_signal_52, new_AGEMA_signal_51, Q0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR1_U1 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_44, new_AGEMA_signal_43, XX[1]}), .c ({new_AGEMA_signal_54, new_AGEMA_signal_53, Q1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) XOR3_U1 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}), .c ({new_AGEMA_signal_56, new_AGEMA_signal_55, Q4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR5_U1 ( .a ({new_AGEMA_signal_48, new_AGEMA_signal_47, XX[2]}), .b ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}), .c ({new_AGEMA_signal_58, new_AGEMA_signal_57, Q6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) XOR6_U1 ( .a ({new_AGEMA_signal_54, new_AGEMA_signal_53, Q1}), .b ({new_AGEMA_signal_58, new_AGEMA_signal_57, Q6}), .c ({new_AGEMA_signal_66, new_AGEMA_signal_65, L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR8_U1 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}), .c ({new_AGEMA_signal_60, new_AGEMA_signal_59, L2}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_26 ( .C (clk), .D (Q0), .Q (new_AGEMA_signal_109) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C (clk), .D (new_AGEMA_signal_51), .Q (new_AGEMA_signal_111) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C (clk), .D (new_AGEMA_signal_52), .Q (new_AGEMA_signal_113) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C (clk), .D (L1), .Q (new_AGEMA_signal_115) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C (clk), .D (new_AGEMA_signal_65), .Q (new_AGEMA_signal_117) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C (clk), .D (new_AGEMA_signal_66), .Q (new_AGEMA_signal_119) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C (clk), .D (XX[2]), .Q (new_AGEMA_signal_121) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C (clk), .D (new_AGEMA_signal_47), .Q (new_AGEMA_signal_123) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C (clk), .D (new_AGEMA_signal_48), .Q (new_AGEMA_signal_125) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C (clk), .D (XX[1]), .Q (new_AGEMA_signal_127) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C (clk), .D (new_AGEMA_signal_43), .Q (new_AGEMA_signal_129) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C (clk), .D (new_AGEMA_signal_44), .Q (new_AGEMA_signal_131) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C (clk), .D (X_s0[1]), .Q (new_AGEMA_signal_133) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C (clk), .D (X_s1[1]), .Q (new_AGEMA_signal_135) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C (clk), .D (X_s2[1]), .Q (new_AGEMA_signal_137) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C (clk), .D (Q6), .Q (new_AGEMA_signal_145) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C (clk), .D (new_AGEMA_signal_57), .Q (new_AGEMA_signal_147) ) ;
    buf_clk new_AGEMA_reg_buffer_66 ( .C (clk), .D (new_AGEMA_signal_58), .Q (new_AGEMA_signal_149) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C (clk), .D (L2), .Q (new_AGEMA_signal_151) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C (clk), .D (new_AGEMA_signal_59), .Q (new_AGEMA_signal_155) ) ;
    buf_clk new_AGEMA_reg_buffer_76 ( .C (clk), .D (new_AGEMA_signal_60), .Q (new_AGEMA_signal_159) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(1)) AND1_U1 ( .a ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}), .b ({new_AGEMA_signal_54, new_AGEMA_signal_53, Q1}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_62, new_AGEMA_signal_61, T0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR2_U1 ( .a ({new_AGEMA_signal_114, new_AGEMA_signal_112, new_AGEMA_signal_110}), .b ({new_AGEMA_signal_62, new_AGEMA_signal_61, T0}), .c ({new_AGEMA_signal_68, new_AGEMA_signal_67, Q2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) AND3_U1 ( .a ({new_AGEMA_signal_40, new_AGEMA_signal_39, n2}), .b ({new_AGEMA_signal_56, new_AGEMA_signal_55, Q4}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_64, new_AGEMA_signal_63, T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR7_U1 ( .a ({new_AGEMA_signal_120, new_AGEMA_signal_118, new_AGEMA_signal_116}), .b ({new_AGEMA_signal_64, new_AGEMA_signal_63, T2}), .c ({new_AGEMA_signal_70, new_AGEMA_signal_69, Q7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR11_U1 ( .a ({new_AGEMA_signal_126, new_AGEMA_signal_124, new_AGEMA_signal_122}), .b ({new_AGEMA_signal_62, new_AGEMA_signal_61, T0}), .c ({new_AGEMA_signal_72, new_AGEMA_signal_71, L3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) XOR12_U1 ( .a ({new_AGEMA_signal_72, new_AGEMA_signal_71, L3}), .b ({new_AGEMA_signal_64, new_AGEMA_signal_63, T2}), .c ({new_AGEMA_signal_80, new_AGEMA_signal_79, YY[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) XOR13_U1 ( .a ({new_AGEMA_signal_132, new_AGEMA_signal_130, new_AGEMA_signal_128}), .b ({new_AGEMA_signal_64, new_AGEMA_signal_63, T2}), .c ({new_AGEMA_signal_74, new_AGEMA_signal_73, YY[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C (clk), .D (new_AGEMA_signal_109), .Q (new_AGEMA_signal_110) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C (clk), .D (new_AGEMA_signal_111), .Q (new_AGEMA_signal_112) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C (clk), .D (new_AGEMA_signal_113), .Q (new_AGEMA_signal_114) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C (clk), .D (new_AGEMA_signal_115), .Q (new_AGEMA_signal_116) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C (clk), .D (new_AGEMA_signal_117), .Q (new_AGEMA_signal_118) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C (clk), .D (new_AGEMA_signal_119), .Q (new_AGEMA_signal_120) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C (clk), .D (new_AGEMA_signal_121), .Q (new_AGEMA_signal_122) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C (clk), .D (new_AGEMA_signal_123), .Q (new_AGEMA_signal_124) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C (clk), .D (new_AGEMA_signal_125), .Q (new_AGEMA_signal_126) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C (clk), .D (new_AGEMA_signal_127), .Q (new_AGEMA_signal_128) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C (clk), .D (new_AGEMA_signal_129), .Q (new_AGEMA_signal_130) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C (clk), .D (new_AGEMA_signal_131), .Q (new_AGEMA_signal_132) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C (clk), .D (new_AGEMA_signal_133), .Q (new_AGEMA_signal_134) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C (clk), .D (new_AGEMA_signal_135), .Q (new_AGEMA_signal_136) ) ;
    buf_clk new_AGEMA_reg_buffer_55 ( .C (clk), .D (new_AGEMA_signal_137), .Q (new_AGEMA_signal_138) ) ;
    buf_clk new_AGEMA_reg_buffer_63 ( .C (clk), .D (new_AGEMA_signal_145), .Q (new_AGEMA_signal_146) ) ;
    buf_clk new_AGEMA_reg_buffer_65 ( .C (clk), .D (new_AGEMA_signal_147), .Q (new_AGEMA_signal_148) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C (clk), .D (new_AGEMA_signal_149), .Q (new_AGEMA_signal_150) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C (clk), .D (new_AGEMA_signal_151), .Q (new_AGEMA_signal_152) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C (clk), .D (new_AGEMA_signal_155), .Q (new_AGEMA_signal_156) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C (clk), .D (new_AGEMA_signal_159), .Q (new_AGEMA_signal_160) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_56 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_139) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C (clk), .D (new_AGEMA_signal_63), .Q (new_AGEMA_signal_141) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C (clk), .D (new_AGEMA_signal_64), .Q (new_AGEMA_signal_143) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C (clk), .D (new_AGEMA_signal_152), .Q (new_AGEMA_signal_153) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C (clk), .D (new_AGEMA_signal_156), .Q (new_AGEMA_signal_157) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C (clk), .D (new_AGEMA_signal_160), .Q (new_AGEMA_signal_161) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C (clk), .D (L3), .Q (new_AGEMA_signal_163) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C (clk), .D (new_AGEMA_signal_71), .Q (new_AGEMA_signal_165) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C (clk), .D (new_AGEMA_signal_72), .Q (new_AGEMA_signal_167) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C (clk), .D (YY[1]), .Q (new_AGEMA_signal_169) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C (clk), .D (new_AGEMA_signal_79), .Q (new_AGEMA_signal_171) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C (clk), .D (new_AGEMA_signal_80), .Q (new_AGEMA_signal_173) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C (clk), .D (YY[0]), .Q (new_AGEMA_signal_175) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C (clk), .D (new_AGEMA_signal_73), .Q (new_AGEMA_signal_177) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C (clk), .D (new_AGEMA_signal_74), .Q (new_AGEMA_signal_179) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(1)) AND2_U1 ( .a ({new_AGEMA_signal_138, new_AGEMA_signal_136, new_AGEMA_signal_134}), .b ({new_AGEMA_signal_68, new_AGEMA_signal_67, Q2}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_76, new_AGEMA_signal_75, T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR4_U1 ( .a ({new_AGEMA_signal_76, new_AGEMA_signal_75, T1}), .b ({new_AGEMA_signal_144, new_AGEMA_signal_142, new_AGEMA_signal_140}), .c ({new_AGEMA_signal_82, new_AGEMA_signal_81, L0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) AND4_U1 ( .a ({new_AGEMA_signal_150, new_AGEMA_signal_148, new_AGEMA_signal_146}), .b ({new_AGEMA_signal_70, new_AGEMA_signal_69, Q7}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_78, new_AGEMA_signal_77, T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR81_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_158, new_AGEMA_signal_154}), .b ({new_AGEMA_signal_76, new_AGEMA_signal_75, T1}), .c ({new_AGEMA_signal_84, new_AGEMA_signal_83, L2_T1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) XOR9_U1 ( .a ({new_AGEMA_signal_84, new_AGEMA_signal_83, L2_T1}), .b ({new_AGEMA_signal_168, new_AGEMA_signal_166, new_AGEMA_signal_164}), .c ({new_AGEMA_signal_86, new_AGEMA_signal_85, YY[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) XOR10_U1 ( .a ({new_AGEMA_signal_82, new_AGEMA_signal_81, L0}), .b ({new_AGEMA_signal_78, new_AGEMA_signal_77, T3}), .c ({new_AGEMA_signal_88, new_AGEMA_signal_87, YY[2]}) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C (clk), .D (new_AGEMA_signal_139), .Q (new_AGEMA_signal_140) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C (clk), .D (new_AGEMA_signal_141), .Q (new_AGEMA_signal_142) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C (clk), .D (new_AGEMA_signal_143), .Q (new_AGEMA_signal_144) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C (clk), .D (new_AGEMA_signal_153), .Q (new_AGEMA_signal_154) ) ;
    buf_clk new_AGEMA_reg_buffer_75 ( .C (clk), .D (new_AGEMA_signal_157), .Q (new_AGEMA_signal_158) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C (clk), .D (new_AGEMA_signal_161), .Q (new_AGEMA_signal_162) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C (clk), .D (new_AGEMA_signal_163), .Q (new_AGEMA_signal_164) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C (clk), .D (new_AGEMA_signal_165), .Q (new_AGEMA_signal_166) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C (clk), .D (new_AGEMA_signal_167), .Q (new_AGEMA_signal_168) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C (clk), .D (new_AGEMA_signal_169), .Q (new_AGEMA_signal_170) ) ;
    buf_clk new_AGEMA_reg_buffer_89 ( .C (clk), .D (new_AGEMA_signal_171), .Q (new_AGEMA_signal_172) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C (clk), .D (new_AGEMA_signal_173), .Q (new_AGEMA_signal_174) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C (clk), .D (new_AGEMA_signal_175), .Q (new_AGEMA_signal_176) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C (clk), .D (new_AGEMA_signal_177), .Q (new_AGEMA_signal_178) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C (clk), .D (new_AGEMA_signal_179), .Q (new_AGEMA_signal_180) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_174, new_AGEMA_signal_172, new_AGEMA_signal_170}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_180, new_AGEMA_signal_178, new_AGEMA_signal_176}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_86, new_AGEMA_signal_85, YY[3]}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_88, new_AGEMA_signal_87, YY[2]}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
