/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_BDDcudd_ClockGating_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input rst ;
    input [4109:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    output Synch ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_6373 ;

    /* cells in depth 0 */
    ClockGatingController #(17) cell_547 ( .clk (clk), .rst (rst), .GatedClk (signal_6373), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_136 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_561, signal_560, signal_559, signal_558, signal_151}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_137 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_569, signal_568, signal_567, signal_566, signal_152}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_138 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_573, signal_572, signal_571, signal_570, signal_153}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_139 ( .s ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_581, signal_580, signal_579, signal_578, signal_154}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_140 ( .s ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_585, signal_584, signal_583, signal_582, signal_155}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_141 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_589, signal_588, signal_587, signal_586, signal_156}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_142 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_593, signal_592, signal_591, signal_590, signal_157}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_143 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_597, signal_596, signal_595, signal_594, signal_158}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_144 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_601, signal_600, signal_599, signal_598, signal_159}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_145 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_605, signal_604, signal_603, signal_602, signal_160}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_146 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_609, signal_608, signal_607, signal_606, signal_161}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_147 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_613, signal_612, signal_611, signal_610, signal_162}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_148 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_617, signal_616, signal_615, signal_614, signal_163}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_149 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_621, signal_620, signal_619, signal_618, signal_164}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_150 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_625, signal_624, signal_623, signal_622, signal_165}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_151 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_629, signal_628, signal_627, signal_626, signal_166}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_152 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_633, signal_632, signal_631, signal_630, signal_167}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_153 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_637, signal_636, signal_635, signal_634, signal_168}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_154 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_641, signal_640, signal_639, signal_638, signal_169}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_155 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_645, signal_644, signal_643, signal_642, signal_170}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_156 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_649, signal_648, signal_647, signal_646, signal_171}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_157 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_653, signal_652, signal_651, signal_650, signal_172}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_158 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_657, signal_656, signal_655, signal_654, signal_173}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_159 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_661, signal_660, signal_659, signal_658, signal_174}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_160 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_665, signal_664, signal_663, signal_662, signal_175}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_161 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_669, signal_668, signal_667, signal_666, signal_176}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_162 ( .s ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_673, signal_672, signal_671, signal_670, signal_177}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_163 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_677, signal_676, signal_675, signal_674, signal_178}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_164 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_681, signal_680, signal_679, signal_678, signal_179}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_165 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_685, signal_684, signal_683, signal_682, signal_180}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_166 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_689, signal_688, signal_687, signal_686, signal_181}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_167 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_693, signal_692, signal_691, signal_690, signal_182}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_168 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_697, signal_696, signal_695, signal_694, signal_183}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_169 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_701, signal_700, signal_699, signal_698, signal_184}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_170 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({signal_705, signal_704, signal_703, signal_702, signal_185}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_171 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .c ({signal_709, signal_708, signal_707, signal_706, signal_186}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_172 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_713, signal_712, signal_711, signal_710, signal_187}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_173 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .c ({signal_717, signal_716, signal_715, signal_714, signal_188}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_174 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({signal_721, signal_720, signal_719, signal_718, signal_189}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_175 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_725, signal_724, signal_723, signal_722, signal_190}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_176 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .c ({signal_729, signal_728, signal_727, signal_726, signal_191}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_177 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .c ({signal_733, signal_732, signal_731, signal_730, signal_192}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_178 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_737, signal_736, signal_735, signal_734, signal_193}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_179 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .c ({signal_741, signal_740, signal_739, signal_738, signal_194}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_180 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .c ({signal_745, signal_744, signal_743, signal_742, signal_195}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_181 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_749, signal_748, signal_747, signal_746, signal_196}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_182 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .c ({signal_753, signal_752, signal_751, signal_750, signal_197}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_183 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .c ({signal_757, signal_756, signal_755, signal_754, signal_198}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_184 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_761, signal_760, signal_759, signal_758, signal_199}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_185 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .c ({signal_765, signal_764, signal_763, signal_762, signal_200}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_186 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .c ({signal_769, signal_768, signal_767, signal_766, signal_201}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_187 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_773, signal_772, signal_771, signal_770, signal_202}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_188 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .c ({signal_777, signal_776, signal_775, signal_774, signal_203}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_189 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .c ({signal_781, signal_780, signal_779, signal_778, signal_204}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_190 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_785, signal_784, signal_783, signal_782, signal_205}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_191 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .c ({signal_789, signal_788, signal_787, signal_786, signal_206}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_192 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .c ({signal_793, signal_792, signal_791, signal_790, signal_207}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_193 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_797, signal_796, signal_795, signal_794, signal_208}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_194 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .c ({signal_801, signal_800, signal_799, signal_798, signal_209}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_195 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .c ({signal_805, signal_804, signal_803, signal_802, signal_210}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_196 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_809, signal_808, signal_807, signal_806, signal_211}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_197 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .c ({signal_813, signal_812, signal_811, signal_810, signal_212}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_198 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .c ({signal_817, signal_816, signal_815, signal_814, signal_213}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_199 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_821, signal_820, signal_819, signal_818, signal_214}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_200 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .c ({signal_825, signal_824, signal_823, signal_822, signal_215}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_201 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .c ({signal_829, signal_828, signal_827, signal_826, signal_216}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_202 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_833, signal_832, signal_831, signal_830, signal_217}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_203 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .c ({signal_837, signal_836, signal_835, signal_834, signal_218}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_204 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .c ({signal_841, signal_840, signal_839, signal_838, signal_219}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_205 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_845, signal_844, signal_843, signal_842, signal_220}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_206 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .c ({signal_849, signal_848, signal_847, signal_846, signal_221}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_207 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .c ({signal_853, signal_852, signal_851, signal_850, signal_222}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_208 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_857, signal_856, signal_855, signal_854, signal_223}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_209 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .c ({signal_861, signal_860, signal_859, signal_858, signal_224}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_210 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .c ({signal_865, signal_864, signal_863, signal_862, signal_225}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_211 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_869, signal_868, signal_867, signal_866, signal_226}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_212 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .c ({signal_873, signal_872, signal_871, signal_870, signal_227}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_213 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .c ({signal_877, signal_876, signal_875, signal_874, signal_228}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_214 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_881, signal_880, signal_879, signal_878, signal_229}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_215 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .c ({signal_885, signal_884, signal_883, signal_882, signal_230}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_216 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .c ({signal_889, signal_888, signal_887, signal_886, signal_231}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_217 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_893, signal_892, signal_891, signal_890, signal_232}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_218 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .c ({signal_897, signal_896, signal_895, signal_894, signal_233}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_219 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .c ({signal_901, signal_900, signal_899, signal_898, signal_234}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_220 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_905, signal_904, signal_903, signal_902, signal_235}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_221 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .c ({signal_909, signal_908, signal_907, signal_906, signal_236}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_222 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .c ({signal_913, signal_912, signal_911, signal_910, signal_237}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_223 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_917, signal_916, signal_915, signal_914, signal_238}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_224 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .c ({signal_921, signal_920, signal_919, signal_918, signal_239}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_225 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890]}), .c ({signal_925, signal_924, signal_923, signal_922, signal_240}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_226 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_929, signal_928, signal_927, signal_926, signal_241}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_227 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910]}), .c ({signal_933, signal_932, signal_931, signal_930, signal_242}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_228 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .c ({signal_937, signal_936, signal_935, signal_934, signal_243}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_229 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_605, signal_604, signal_603, signal_602, signal_160}), .a ({signal_669, signal_668, signal_667, signal_666, signal_176}), .clk (clk), .r ({Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_945, signal_944, signal_943, signal_942, signal_244}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_230 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .c ({signal_949, signal_948, signal_947, signal_946, signal_245}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_231 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950]}), .c ({signal_953, signal_952, signal_951, signal_950, signal_246}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_232 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_957, signal_956, signal_955, signal_954, signal_247}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_233 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970]}), .c ({signal_961, signal_960, signal_959, signal_958, signal_248}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_234 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .c ({signal_965, signal_964, signal_963, signal_962, signal_249}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_235 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_969, signal_968, signal_967, signal_966, signal_250}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_236 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .c ({signal_973, signal_972, signal_971, signal_970, signal_251}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_237 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010]}), .c ({signal_977, signal_976, signal_975, signal_974, signal_252}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_238 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_981, signal_980, signal_979, signal_978, signal_253}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_239 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030]}), .c ({signal_985, signal_984, signal_983, signal_982, signal_254}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_240 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .c ({signal_989, signal_988, signal_987, signal_986, signal_255}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_241 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_993, signal_992, signal_991, signal_990, signal_256}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_242 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .c ({signal_997, signal_996, signal_995, signal_994, signal_257}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_243 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070]}), .c ({signal_1001, signal_1000, signal_999, signal_998, signal_258}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_244 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1005, signal_1004, signal_1003, signal_1002, signal_259}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_245 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090]}), .c ({signal_1009, signal_1008, signal_1007, signal_1006, signal_260}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_246 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .c ({signal_1013, signal_1012, signal_1011, signal_1010, signal_261}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_247 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1017, signal_1016, signal_1015, signal_1014, signal_262}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_248 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .c ({signal_1021, signal_1020, signal_1019, signal_1018, signal_263}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_249 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130]}), .c ({signal_1025, signal_1024, signal_1023, signal_1022, signal_264}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_250 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1029, signal_1028, signal_1027, signal_1026, signal_265}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_251 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150]}), .c ({signal_1033, signal_1032, signal_1031, signal_1030, signal_266}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_252 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .c ({signal_1037, signal_1036, signal_1035, signal_1034, signal_267}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_253 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1041, signal_1040, signal_1039, signal_1038, signal_268}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_254 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .c ({signal_1045, signal_1044, signal_1043, signal_1042, signal_269}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_255 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190]}), .c ({signal_1049, signal_1048, signal_1047, signal_1046, signal_270}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_256 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1053, signal_1052, signal_1051, signal_1050, signal_271}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_257 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_581, signal_580, signal_579, signal_578, signal_154}), .clk (clk), .r ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210]}), .c ({signal_1057, signal_1056, signal_1055, signal_1054, signal_272}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_258 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .c ({signal_1061, signal_1060, signal_1059, signal_1058, signal_273}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_259 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_621, signal_620, signal_619, signal_618, signal_164}), .clk (clk), .r ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_1065, signal_1064, signal_1063, signal_1062, signal_274}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_260 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .c ({signal_1069, signal_1068, signal_1067, signal_1066, signal_275}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_261 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250]}), .c ({signal_1073, signal_1072, signal_1071, signal_1070, signal_276}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_262 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_1077, signal_1076, signal_1075, signal_1074, signal_277}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_263 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270]}), .c ({signal_1081, signal_1080, signal_1079, signal_1078, signal_278}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_264 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .c ({signal_1085, signal_1084, signal_1083, signal_1082, signal_279}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_265 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_1089, signal_1088, signal_1087, signal_1086, signal_280}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_266 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .c ({signal_1093, signal_1092, signal_1091, signal_1090, signal_281}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_267 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_569, signal_568, signal_567, signal_566, signal_152}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310]}), .c ({signal_1097, signal_1096, signal_1095, signal_1094, signal_282}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_268 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_593, signal_592, signal_591, signal_590, signal_157}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_1101, signal_1100, signal_1099, signal_1098, signal_283}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_269 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330]}), .c ({signal_1105, signal_1104, signal_1103, signal_1102, signal_284}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_270 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .c ({signal_1109, signal_1108, signal_1107, signal_1106, signal_285}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_271 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_1113, signal_1112, signal_1111, signal_1110, signal_286}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_272 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .c ({signal_1117, signal_1116, signal_1115, signal_1114, signal_287}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_273 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370]}), .c ({signal_1121, signal_1120, signal_1119, signal_1118, signal_288}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_274 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_1125, signal_1124, signal_1123, signal_1122, signal_289}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_275 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390]}), .c ({signal_1129, signal_1128, signal_1127, signal_1126, signal_290}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_276 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_589, signal_588, signal_587, signal_586, signal_156}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .c ({signal_1133, signal_1132, signal_1131, signal_1130, signal_291}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_277 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_561, signal_560, signal_559, signal_558, signal_151}), .clk (clk), .r ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_1137, signal_1136, signal_1135, signal_1134, signal_292}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_278 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .c ({signal_1141, signal_1140, signal_1139, signal_1138, signal_293}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_279 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430]}), .c ({signal_1145, signal_1144, signal_1143, signal_1142, signal_294}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_280 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_1149, signal_1148, signal_1147, signal_1146, signal_295}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_281 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450]}), .c ({signal_1153, signal_1152, signal_1151, signal_1150, signal_296}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_282 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .c ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_283 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_1161, signal_1160, signal_1159, signal_1158, signal_298}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_284 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_693, signal_692, signal_691, signal_690, signal_182}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .c ({signal_1165, signal_1164, signal_1163, signal_1162, signal_299}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_285 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_673, signal_672, signal_671, signal_670, signal_177}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490]}), .c ({signal_1169, signal_1168, signal_1167, signal_1166, signal_300}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_286 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_1173, signal_1172, signal_1171, signal_1170, signal_301}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_287 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_601, signal_600, signal_599, signal_598, signal_159}), .a ({signal_609, signal_608, signal_607, signal_606, signal_161}), .clk (clk), .r ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510]}), .c ({signal_1177, signal_1176, signal_1175, signal_1174, signal_302}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_288 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .c ({signal_1181, signal_1180, signal_1179, signal_1178, signal_303}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_289 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_1185, signal_1184, signal_1183, signal_1182, signal_304}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_290 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_641, signal_640, signal_639, signal_638, signal_169}), .a ({signal_585, signal_584, signal_583, signal_582, signal_155}), .clk (clk), .r ({Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .c ({signal_1189, signal_1188, signal_1187, signal_1186, signal_305}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_291 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_681, signal_680, signal_679, signal_678, signal_179}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550]}), .c ({signal_1193, signal_1192, signal_1191, signal_1190, signal_306}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_292 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_585, signal_584, signal_583, signal_582, signal_155}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_1197, signal_1196, signal_1195, signal_1194, signal_307}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_293 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_625, signal_624, signal_623, signal_622, signal_165}), .clk (clk), .r ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570]}), .c ({signal_1201, signal_1200, signal_1199, signal_1198, signal_308}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_294 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .c ({signal_1205, signal_1204, signal_1203, signal_1202, signal_309}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_295 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_637, signal_636, signal_635, signal_634, signal_168}), .a ({signal_613, signal_612, signal_611, signal_610, signal_162}), .clk (clk), .r ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_1209, signal_1208, signal_1207, signal_1206, signal_310}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_296 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_573, signal_572, signal_571, signal_570, signal_153}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .c ({signal_1213, signal_1212, signal_1211, signal_1210, signal_311}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_297 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610]}), .c ({signal_1217, signal_1216, signal_1215, signal_1214, signal_312}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_298 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_597, signal_596, signal_595, signal_594, signal_158}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_1221, signal_1220, signal_1219, signal_1218, signal_313}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_299 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_581, signal_580, signal_579, signal_578, signal_154}), .a ({signal_589, signal_588, signal_587, signal_586, signal_156}), .clk (clk), .r ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630]}), .c ({signal_1225, signal_1224, signal_1223, signal_1222, signal_314}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_300 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .c ({signal_1229, signal_1228, signal_1227, signal_1226, signal_315}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_301 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_661, signal_660, signal_659, signal_658, signal_174}), .clk (clk), .r ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_1233, signal_1232, signal_1231, signal_1230, signal_316}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_302 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_661, signal_660, signal_659, signal_658, signal_174}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .c ({signal_1237, signal_1236, signal_1235, signal_1234, signal_317}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_303 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_625, signal_624, signal_623, signal_622, signal_165}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670]}), .c ({signal_1241, signal_1240, signal_1239, signal_1238, signal_318}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_304 ( .s ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_665, signal_664, signal_663, signal_662, signal_175}), .a ({signal_573, signal_572, signal_571, signal_570, signal_153}), .clk (clk), .r ({Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_1245, signal_1244, signal_1243, signal_1242, signal_319}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_305 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_881, signal_880, signal_879, signal_878, signal_229}), .clk (clk), .r ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690]}), .c ({signal_1249, signal_1248, signal_1247, signal_1246, signal_320}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_306 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1237, signal_1236, signal_1235, signal_1234, signal_317}), .a ({signal_905, signal_904, signal_903, signal_902, signal_235}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .c ({signal_1253, signal_1252, signal_1251, signal_1250, signal_321}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_307 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1185, signal_1184, signal_1183, signal_1182, signal_304}), .a ({signal_1133, signal_1132, signal_1131, signal_1130, signal_291}), .clk (clk), .r ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_1257, signal_1256, signal_1255, signal_1254, signal_322}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_308 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1213, signal_1212, signal_1211, signal_1210, signal_311}), .a ({signal_569, signal_568, signal_567, signal_566, signal_152}), .clk (clk), .r ({Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .c ({signal_1261, signal_1260, signal_1259, signal_1258, signal_323}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_309 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_817, signal_816, signal_815, signal_814, signal_213}), .a ({signal_981, signal_980, signal_979, signal_978, signal_253}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730]}), .c ({signal_1265, signal_1264, signal_1263, signal_1262, signal_324}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_310 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_949, signal_948, signal_947, signal_946, signal_245}), .a ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}), .clk (clk), .r ({Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_1269, signal_1268, signal_1267, signal_1266, signal_325}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_311 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_709, signal_708, signal_707, signal_706, signal_186}), .clk (clk), .r ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750]}), .c ({signal_1273, signal_1272, signal_1271, signal_1270, signal_326}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_312 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_693, signal_692, signal_691, signal_690, signal_182}), .a ({signal_1033, signal_1032, signal_1031, signal_1030, signal_266}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .c ({signal_1277, signal_1276, signal_1275, signal_1274, signal_327}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_313 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_761, signal_760, signal_759, signal_758, signal_199}), .a ({signal_869, signal_868, signal_867, signal_866, signal_226}), .clk (clk), .r ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_1281, signal_1280, signal_1279, signal_1278, signal_328}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_314 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1005, signal_1004, signal_1003, signal_1002, signal_259}), .a ({signal_1121, signal_1120, signal_1119, signal_1118, signal_288}), .clk (clk), .r ({Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .c ({signal_1285, signal_1284, signal_1283, signal_1282, signal_329}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_315 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1129, signal_1128, signal_1127, signal_1126, signal_290}), .a ({signal_1021, signal_1020, signal_1019, signal_1018, signal_263}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790]}), .c ({signal_1289, signal_1288, signal_1287, signal_1286, signal_330}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_316 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1137, signal_1136, signal_1135, signal_1134, signal_292}), .a ({signal_1237, signal_1236, signal_1235, signal_1234, signal_317}), .clk (clk), .r ({Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_1293, signal_1292, signal_1291, signal_1290, signal_331}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_317 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_825, signal_824, signal_823, signal_822, signal_215}), .a ({signal_665, signal_664, signal_663, signal_662, signal_175}), .clk (clk), .r ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810]}), .c ({signal_1297, signal_1296, signal_1295, signal_1294, signal_332}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_318 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_853, signal_852, signal_851, signal_850, signal_222}), .a ({signal_1001, signal_1000, signal_999, signal_998, signal_258}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .c ({signal_1301, signal_1300, signal_1299, signal_1298, signal_333}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_319 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_785, signal_784, signal_783, signal_782, signal_205}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_1305, signal_1304, signal_1303, signal_1302, signal_334}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_320 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_917, signal_916, signal_915, signal_914, signal_238}), .a ({signal_901, signal_900, signal_899, signal_898, signal_234}), .clk (clk), .r ({Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .c ({signal_1309, signal_1308, signal_1307, signal_1306, signal_335}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_321 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_841, signal_840, signal_839, signal_838, signal_219}), .a ({signal_817, signal_816, signal_815, signal_814, signal_213}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850]}), .c ({signal_1313, signal_1312, signal_1311, signal_1310, signal_336}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_322 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1229, signal_1228, signal_1227, signal_1226, signal_315}), .a ({signal_1093, signal_1092, signal_1091, signal_1090, signal_281}), .clk (clk), .r ({Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_1317, signal_1316, signal_1315, signal_1314, signal_337}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_323 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1141, signal_1140, signal_1139, signal_1138, signal_293}), .a ({signal_773, signal_772, signal_771, signal_770, signal_202}), .clk (clk), .r ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870]}), .c ({signal_1321, signal_1320, signal_1319, signal_1318, signal_338}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_324 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1221, signal_1220, signal_1219, signal_1218, signal_313}), .a ({signal_641, signal_640, signal_639, signal_638, signal_169}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .c ({signal_1325, signal_1324, signal_1323, signal_1322, signal_339}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_325 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_845, signal_844, signal_843, signal_842, signal_220}), .a ({signal_881, signal_880, signal_879, signal_878, signal_229}), .clk (clk), .r ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_1329, signal_1328, signal_1327, signal_1326, signal_340}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_326 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_937, signal_936, signal_935, signal_934, signal_243}), .a ({signal_913, signal_912, signal_911, signal_910, signal_237}), .clk (clk), .r ({Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .c ({signal_1333, signal_1332, signal_1331, signal_1330, signal_341}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_327 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_933, signal_932, signal_931, signal_930, signal_242}), .a ({signal_1125, signal_1124, signal_1123, signal_1122, signal_289}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910]}), .c ({signal_1337, signal_1336, signal_1335, signal_1334, signal_342}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_328 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_829, signal_828, signal_827, signal_826, signal_216}), .a ({signal_1233, signal_1232, signal_1231, signal_1230, signal_316}), .clk (clk), .r ({Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_1341, signal_1340, signal_1339, signal_1338, signal_343}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_329 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_913, signal_912, signal_911, signal_910, signal_237}), .a ({signal_1101, signal_1100, signal_1099, signal_1098, signal_283}), .clk (clk), .r ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930]}), .c ({signal_1345, signal_1344, signal_1343, signal_1342, signal_344}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_330 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1245, signal_1244, signal_1243, signal_1242, signal_319}), .a ({signal_965, signal_964, signal_963, signal_962, signal_249}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .c ({signal_1349, signal_1348, signal_1347, signal_1346, signal_345}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_331 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_989, signal_988, signal_987, signal_986, signal_255}), .a ({signal_937, signal_936, signal_935, signal_934, signal_243}), .clk (clk), .r ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_1353, signal_1352, signal_1351, signal_1350, signal_346}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_332 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_793, signal_792, signal_791, signal_790, signal_207}), .a ({signal_677, signal_676, signal_675, signal_674, signal_178}), .clk (clk), .r ({Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .c ({signal_1357, signal_1356, signal_1355, signal_1354, signal_347}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_333 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1049, signal_1048, signal_1047, signal_1046, signal_270}), .a ({signal_985, signal_984, signal_983, signal_982, signal_254}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970]}), .c ({signal_1361, signal_1360, signal_1359, signal_1358, signal_348}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_334 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1013, signal_1012, signal_1011, signal_1010, signal_261}), .a ({signal_1229, signal_1228, signal_1227, signal_1226, signal_315}), .clk (clk), .r ({Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_1365, signal_1364, signal_1363, signal_1362, signal_349}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_335 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_569, signal_568, signal_567, signal_566, signal_152}), .a ({signal_965, signal_964, signal_963, signal_962, signal_249}), .clk (clk), .r ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990]}), .c ({signal_1369, signal_1368, signal_1367, signal_1366, signal_350}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_336 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_989, signal_988, signal_987, signal_986, signal_255}), .a ({signal_1089, signal_1088, signal_1087, signal_1086, signal_280}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .c ({signal_1373, signal_1372, signal_1371, signal_1370, signal_351}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_337 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_893, signal_892, signal_891, signal_890, signal_232}), .a ({signal_729, signal_728, signal_727, signal_726, signal_191}), .clk (clk), .r ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_1377, signal_1376, signal_1375, signal_1374, signal_352}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_338 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1209, signal_1208, signal_1207, signal_1206, signal_310}), .a ({signal_1137, signal_1136, signal_1135, signal_1134, signal_292}), .clk (clk), .r ({Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .c ({signal_1381, signal_1380, signal_1379, signal_1378, signal_353}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_339 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_961, signal_960, signal_959, signal_958, signal_248}), .a ({signal_889, signal_888, signal_887, signal_886, signal_231}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030]}), .c ({signal_1385, signal_1384, signal_1383, signal_1382, signal_354}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_340 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1169, signal_1168, signal_1167, signal_1166, signal_300}), .a ({signal_1205, signal_1204, signal_1203, signal_1202, signal_309}), .clk (clk), .r ({Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_1389, signal_1388, signal_1387, signal_1386, signal_355}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_341 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_857, signal_856, signal_855, signal_854, signal_223}), .a ({signal_1109, signal_1108, signal_1107, signal_1106, signal_285}), .clk (clk), .r ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050]}), .c ({signal_1393, signal_1392, signal_1391, signal_1390, signal_356}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_342 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_917, signal_916, signal_915, signal_914, signal_238}), .a ({signal_969, signal_968, signal_967, signal_966, signal_250}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .c ({signal_1397, signal_1396, signal_1395, signal_1394, signal_357}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_343 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_909, signal_908, signal_907, signal_906, signal_236}), .a ({signal_633, signal_632, signal_631, signal_630, signal_167}), .clk (clk), .r ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_1401, signal_1400, signal_1399, signal_1398, signal_358}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_344 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1057, signal_1056, signal_1055, signal_1054, signal_272}), .a ({signal_893, signal_892, signal_891, signal_890, signal_232}), .clk (clk), .r ({Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .c ({signal_1405, signal_1404, signal_1403, signal_1402, signal_359}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_345 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_649, signal_648, signal_647, signal_646, signal_171}), .a ({signal_1185, signal_1184, signal_1183, signal_1182, signal_304}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090]}), .c ({signal_1409, signal_1408, signal_1407, signal_1406, signal_360}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_346 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1093, signal_1092, signal_1091, signal_1090, signal_281}), .a ({signal_1109, signal_1108, signal_1107, signal_1106, signal_285}), .clk (clk), .r ({Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_1413, signal_1412, signal_1411, signal_1410, signal_361}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_347 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_733, signal_732, signal_731, signal_730, signal_192}), .a ({signal_965, signal_964, signal_963, signal_962, signal_249}), .clk (clk), .r ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110]}), .c ({signal_1417, signal_1416, signal_1415, signal_1414, signal_362}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_348 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1161, signal_1160, signal_1159, signal_1158, signal_298}), .a ({signal_697, signal_696, signal_695, signal_694, signal_183}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .c ({signal_1421, signal_1420, signal_1419, signal_1418, signal_363}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_349 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_865, signal_864, signal_863, signal_862, signal_225}), .a ({signal_701, signal_700, signal_699, signal_698, signal_184}), .clk (clk), .r ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_1425, signal_1424, signal_1423, signal_1422, signal_364}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_350 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_677, signal_676, signal_675, signal_674, signal_178}), .a ({signal_1117, signal_1116, signal_1115, signal_1114, signal_287}), .clk (clk), .r ({Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .c ({signal_1429, signal_1428, signal_1427, signal_1426, signal_365}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_351 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_861, signal_860, signal_859, signal_858, signal_224}), .a ({signal_685, signal_684, signal_683, signal_682, signal_180}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150]}), .c ({signal_1433, signal_1432, signal_1431, signal_1430, signal_366}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_352 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_725, signal_724, signal_723, signal_722, signal_190}), .a ({signal_653, signal_652, signal_651, signal_650, signal_172}), .clk (clk), .r ({Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_1437, signal_1436, signal_1435, signal_1434, signal_367}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_353 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_997, signal_996, signal_995, signal_994, signal_257}), .a ({signal_753, signal_752, signal_751, signal_750, signal_197}), .clk (clk), .r ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170]}), .c ({signal_1441, signal_1440, signal_1439, signal_1438, signal_368}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_354 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_617, signal_616, signal_615, signal_614, signal_163}), .a ({signal_1025, signal_1024, signal_1023, signal_1022, signal_264}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .c ({signal_1445, signal_1444, signal_1443, signal_1442, signal_369}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_355 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1017, signal_1016, signal_1015, signal_1014, signal_262}), .a ({signal_637, signal_636, signal_635, signal_634, signal_168}), .clk (clk), .r ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_1449, signal_1448, signal_1447, signal_1446, signal_370}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_356 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_721, signal_720, signal_719, signal_718, signal_189}), .a ({signal_1201, signal_1200, signal_1199, signal_1198, signal_308}), .clk (clk), .r ({Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .c ({signal_1453, signal_1452, signal_1451, signal_1450, signal_371}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_357 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_561, signal_560, signal_559, signal_558, signal_151}), .a ({signal_969, signal_968, signal_967, signal_966, signal_250}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210]}), .c ({signal_1457, signal_1456, signal_1455, signal_1454, signal_372}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_358 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1029, signal_1028, signal_1027, signal_1026, signal_265}), .a ({signal_1021, signal_1020, signal_1019, signal_1018, signal_263}), .clk (clk), .r ({Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_1461, signal_1460, signal_1459, signal_1458, signal_373}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_359 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1081, signal_1080, signal_1079, signal_1078, signal_278}), .a ({signal_921, signal_920, signal_919, signal_918, signal_239}), .clk (clk), .r ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230]}), .c ({signal_1465, signal_1464, signal_1463, signal_1462, signal_374}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_360 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_713, signal_712, signal_711, signal_710, signal_187}), .a ({signal_821, signal_820, signal_819, signal_818, signal_214}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .c ({signal_1469, signal_1468, signal_1467, signal_1466, signal_375}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_361 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_725, signal_724, signal_723, signal_722, signal_190}), .a ({signal_749, signal_748, signal_747, signal_746, signal_196}), .clk (clk), .r ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_1473, signal_1472, signal_1471, signal_1470, signal_376}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_362 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1101, signal_1100, signal_1099, signal_1098, signal_283}), .a ({signal_645, signal_644, signal_643, signal_642, signal_170}), .clk (clk), .r ({Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .c ({signal_1477, signal_1476, signal_1475, signal_1474, signal_377}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_363 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1013, signal_1012, signal_1011, signal_1010, signal_261}), .a ({signal_1149, signal_1148, signal_1147, signal_1146, signal_295}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270]}), .c ({signal_1481, signal_1480, signal_1479, signal_1478, signal_378}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_364 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_837, signal_836, signal_835, signal_834, signal_218}), .a ({signal_717, signal_716, signal_715, signal_714, signal_188}), .clk (clk), .r ({Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_1485, signal_1484, signal_1483, signal_1482, signal_379}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_365 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1105, signal_1104, signal_1103, signal_1102, signal_284}), .a ({signal_769, signal_768, signal_767, signal_766, signal_201}), .clk (clk), .r ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290]}), .c ({signal_1489, signal_1488, signal_1487, signal_1486, signal_380}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_366 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_609, signal_608, signal_607, signal_606, signal_161}), .a ({signal_1061, signal_1060, signal_1059, signal_1058, signal_273}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .c ({signal_1493, signal_1492, signal_1491, signal_1490, signal_381}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_367 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_609, signal_608, signal_607, signal_606, signal_161}), .a ({signal_753, signal_752, signal_751, signal_750, signal_197}), .clk (clk), .r ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_1497, signal_1496, signal_1495, signal_1494, signal_382}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_368 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_765, signal_764, signal_763, signal_762, signal_200}), .a ({signal_621, signal_620, signal_619, signal_618, signal_164}), .clk (clk), .r ({Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .c ({signal_1501, signal_1500, signal_1499, signal_1498, signal_383}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_369 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1181, signal_1180, signal_1179, signal_1178, signal_303}), .a ({signal_1045, signal_1044, signal_1043, signal_1042, signal_269}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330]}), .c ({signal_1505, signal_1504, signal_1503, signal_1502, signal_384}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_370 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_961, signal_960, signal_959, signal_958, signal_248}), .a ({signal_993, signal_992, signal_991, signal_990, signal_256}), .clk (clk), .r ({Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_1509, signal_1508, signal_1507, signal_1506, signal_385}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_371 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_645, signal_644, signal_643, signal_642, signal_170}), .a ({signal_1013, signal_1012, signal_1011, signal_1010, signal_261}), .clk (clk), .r ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350]}), .c ({signal_1513, signal_1512, signal_1511, signal_1510, signal_386}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_372 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_905, signal_904, signal_903, signal_902, signal_235}), .a ({signal_1189, signal_1188, signal_1187, signal_1186, signal_305}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .c ({signal_1517, signal_1516, signal_1515, signal_1514, signal_387}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_373 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_865, signal_864, signal_863, signal_862, signal_225}), .a ({signal_685, signal_684, signal_683, signal_682, signal_180}), .clk (clk), .r ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_1521, signal_1520, signal_1519, signal_1518, signal_388}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_374 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_825, signal_824, signal_823, signal_822, signal_215}), .a ({signal_645, signal_644, signal_643, signal_642, signal_170}), .clk (clk), .r ({Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .c ({signal_1525, signal_1524, signal_1523, signal_1522, signal_389}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_375 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_957, signal_956, signal_955, signal_954, signal_247}), .a ({signal_1073, signal_1072, signal_1071, signal_1070, signal_276}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390]}), .c ({signal_1529, signal_1528, signal_1527, signal_1526, signal_390}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_376 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_833, signal_832, signal_831, signal_830, signal_217}), .a ({signal_841, signal_840, signal_839, signal_838, signal_219}), .clk (clk), .r ({Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_1533, signal_1532, signal_1531, signal_1530, signal_391}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_377 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_849, signal_848, signal_847, signal_846, signal_221}), .a ({signal_813, signal_812, signal_811, signal_810, signal_212}), .clk (clk), .r ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410]}), .c ({signal_1537, signal_1536, signal_1535, signal_1534, signal_392}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_378 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_613, signal_612, signal_611, signal_610, signal_162}), .a ({signal_977, signal_976, signal_975, signal_974, signal_252}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .c ({signal_1541, signal_1540, signal_1539, signal_1538, signal_393}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_379 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_729, signal_728, signal_727, signal_726, signal_191}), .a ({signal_777, signal_776, signal_775, signal_774, signal_203}), .clk (clk), .r ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_1545, signal_1544, signal_1543, signal_1542, signal_394}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_380 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}), .a ({signal_909, signal_908, signal_907, signal_906, signal_236}), .clk (clk), .r ({Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .c ({signal_1549, signal_1548, signal_1547, signal_1546, signal_395}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_381 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_821, signal_820, signal_819, signal_818, signal_214}), .a ({signal_569, signal_568, signal_567, signal_566, signal_152}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450]}), .c ({signal_1553, signal_1552, signal_1551, signal_1550, signal_396}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_382 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_985, signal_984, signal_983, signal_982, signal_254}), .a ({signal_721, signal_720, signal_719, signal_718, signal_189}), .clk (clk), .r ({Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_1557, signal_1556, signal_1555, signal_1554, signal_397}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_383 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_985, signal_984, signal_983, signal_982, signal_254}), .a ({signal_841, signal_840, signal_839, signal_838, signal_219}), .clk (clk), .r ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470]}), .c ({signal_1561, signal_1560, signal_1559, signal_1558, signal_398}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_384 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_805, signal_804, signal_803, signal_802, signal_210}), .a ({signal_733, signal_732, signal_731, signal_730, signal_192}), .clk (clk), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .c ({signal_1565, signal_1564, signal_1563, signal_1562, signal_399}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_385 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1081, signal_1080, signal_1079, signal_1078, signal_278}), .a ({signal_1037, signal_1036, signal_1035, signal_1034, signal_267}), .clk (clk), .r ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_1569, signal_1568, signal_1567, signal_1566, signal_400}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_386 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_813, signal_812, signal_811, signal_810, signal_212}), .a ({signal_825, signal_824, signal_823, signal_822, signal_215}), .clk (clk), .r ({Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .c ({signal_1573, signal_1572, signal_1571, signal_1570, signal_401}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_387 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1153, signal_1152, signal_1151, signal_1150, signal_296}), .a ({signal_1053, signal_1052, signal_1051, signal_1050, signal_271}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510]}), .c ({signal_1577, signal_1576, signal_1575, signal_1574, signal_402}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_388 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_657, signal_656, signal_655, signal_654, signal_173}), .a ({signal_737, signal_736, signal_735, signal_734, signal_193}), .clk (clk), .r ({Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_1581, signal_1580, signal_1579, signal_1578, signal_403}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_389 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_801, signal_800, signal_799, signal_798, signal_209}), .a ({signal_1085, signal_1084, signal_1083, signal_1082, signal_279}), .clk (clk), .r ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530]}), .c ({signal_1585, signal_1584, signal_1583, signal_1582, signal_404}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_390 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_973, signal_972, signal_971, signal_970, signal_251}), .a ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}), .clk (clk), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .c ({signal_1589, signal_1588, signal_1587, signal_1586, signal_405}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_391 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_777, signal_776, signal_775, signal_774, signal_203}), .a ({signal_597, signal_596, signal_595, signal_594, signal_158}), .clk (clk), .r ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_1593, signal_1592, signal_1591, signal_1590, signal_406}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_392 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_937, signal_936, signal_935, signal_934, signal_243}), .a ({signal_1113, signal_1112, signal_1111, signal_1110, signal_286}), .clk (clk), .r ({Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .c ({signal_1597, signal_1596, signal_1595, signal_1594, signal_407}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_393 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_901, signal_900, signal_899, signal_898, signal_234}), .a ({signal_689, signal_688, signal_687, signal_686, signal_181}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570]}), .c ({signal_1601, signal_1600, signal_1599, signal_1598, signal_408}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_394 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1145, signal_1144, signal_1143, signal_1142, signal_294}), .a ({signal_989, signal_988, signal_987, signal_986, signal_255}), .clk (clk), .r ({Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_1605, signal_1604, signal_1603, signal_1602, signal_409}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_395 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_901, signal_900, signal_899, signal_898, signal_234}), .a ({signal_1041, signal_1040, signal_1039, signal_1038, signal_268}), .clk (clk), .r ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590]}), .c ({signal_1609, signal_1608, signal_1607, signal_1606, signal_410}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_396 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_929, signal_928, signal_927, signal_926, signal_241}), .a ({signal_645, signal_644, signal_643, signal_642, signal_170}), .clk (clk), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .c ({signal_1613, signal_1612, signal_1611, signal_1610, signal_411}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_397 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_729, signal_728, signal_727, signal_726, signal_191}), .a ({signal_897, signal_896, signal_895, signal_894, signal_233}), .clk (clk), .r ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_1617, signal_1616, signal_1615, signal_1614, signal_412}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_398 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1021, signal_1020, signal_1019, signal_1018, signal_263}), .a ({signal_737, signal_736, signal_735, signal_734, signal_193}), .clk (clk), .r ({Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .c ({signal_1621, signal_1620, signal_1619, signal_1618, signal_413}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_399 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1233, signal_1232, signal_1231, signal_1230, signal_316}), .a ({signal_841, signal_840, signal_839, signal_838, signal_219}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630]}), .c ({signal_1625, signal_1624, signal_1623, signal_1622, signal_414}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_400 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_885, signal_884, signal_883, signal_882, signal_230}), .a ({signal_1217, signal_1216, signal_1215, signal_1214, signal_312}), .clk (clk), .r ({Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_1629, signal_1628, signal_1627, signal_1626, signal_415}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_401 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1077, signal_1076, signal_1075, signal_1074, signal_277}), .a ({signal_833, signal_832, signal_831, signal_830, signal_217}), .clk (clk), .r ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650]}), .c ({signal_1633, signal_1632, signal_1631, signal_1630, signal_416}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_402 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}), .a ({signal_1181, signal_1180, signal_1179, signal_1178, signal_303}), .clk (clk), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .c ({signal_1637, signal_1636, signal_1635, signal_1634, signal_417}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_403 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1173, signal_1172, signal_1171, signal_1170, signal_301}), .a ({signal_1069, signal_1068, signal_1067, signal_1066, signal_275}), .clk (clk), .r ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_1641, signal_1640, signal_1639, signal_1638, signal_418}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_404 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1025, signal_1024, signal_1023, signal_1022, signal_264}), .a ({signal_781, signal_780, signal_779, signal_778, signal_204}), .clk (clk), .r ({Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .c ({signal_1645, signal_1644, signal_1643, signal_1642, signal_419}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_405 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_745, signal_744, signal_743, signal_742, signal_195}), .a ({signal_853, signal_852, signal_851, signal_850, signal_222}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690]}), .c ({signal_1649, signal_1648, signal_1647, signal_1646, signal_420}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_406 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_877, signal_876, signal_875, signal_874, signal_228}), .a ({signal_933, signal_932, signal_931, signal_930, signal_242}), .clk (clk), .r ({Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_1653, signal_1652, signal_1651, signal_1650, signal_421}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_407 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_977, signal_976, signal_975, signal_974, signal_252}), .a ({signal_1237, signal_1236, signal_1235, signal_1234, signal_317}), .clk (clk), .r ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710]}), .c ({signal_1657, signal_1656, signal_1655, signal_1654, signal_422}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_408 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_841, signal_840, signal_839, signal_838, signal_219}), .a ({signal_713, signal_712, signal_711, signal_710, signal_187}), .clk (clk), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .c ({signal_1661, signal_1660, signal_1659, signal_1658, signal_423}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_409 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1157, signal_1156, signal_1155, signal_1154, signal_297}), .a ({signal_673, signal_672, signal_671, signal_670, signal_177}), .clk (clk), .r ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_1665, signal_1664, signal_1663, signal_1662, signal_424}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_410 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_713, signal_712, signal_711, signal_710, signal_187}), .a ({signal_669, signal_668, signal_667, signal_666, signal_176}), .clk (clk), .r ({Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .c ({signal_1669, signal_1668, signal_1667, signal_1666, signal_425}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_411 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_725, signal_724, signal_723, signal_722, signal_190}), .a ({signal_873, signal_872, signal_871, signal_870, signal_227}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750]}), .c ({signal_1673, signal_1672, signal_1671, signal_1670, signal_426}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_412 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1073, signal_1072, signal_1071, signal_1070, signal_276}), .a ({signal_593, signal_592, signal_591, signal_590, signal_157}), .clk (clk), .r ({Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_1677, signal_1676, signal_1675, signal_1674, signal_427}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_413 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_933, signal_932, signal_931, signal_930, signal_242}), .a ({signal_805, signal_804, signal_803, signal_802, signal_210}), .clk (clk), .r ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770]}), .c ({signal_1681, signal_1680, signal_1679, signal_1678, signal_428}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_414 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_757, signal_756, signal_755, signal_754, signal_198}), .a ({signal_793, signal_792, signal_791, signal_790, signal_207}), .clk (clk), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .c ({signal_1685, signal_1684, signal_1683, signal_1682, signal_429}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_415 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1025, signal_1024, signal_1023, signal_1022, signal_264}), .a ({signal_1241, signal_1240, signal_1239, signal_1238, signal_318}), .clk (clk), .r ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_1689, signal_1688, signal_1687, signal_1686, signal_430}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_416 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_669, signal_668, signal_667, signal_666, signal_176}), .a ({signal_1057, signal_1056, signal_1055, signal_1054, signal_272}), .clk (clk), .r ({Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .c ({signal_1693, signal_1692, signal_1691, signal_1690, signal_431}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_417 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1161, signal_1160, signal_1159, signal_1158, signal_298}), .a ({signal_789, signal_788, signal_787, signal_786, signal_206}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810]}), .c ({signal_1697, signal_1696, signal_1695, signal_1694, signal_432}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_418 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_925, signal_924, signal_923, signal_922, signal_240}), .a ({signal_705, signal_704, signal_703, signal_702, signal_185}), .clk (clk), .r ({Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_1701, signal_1700, signal_1699, signal_1698, signal_433}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_419 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1129, signal_1128, signal_1127, signal_1126, signal_290}), .a ({signal_925, signal_924, signal_923, signal_922, signal_240}), .clk (clk), .r ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830]}), .c ({signal_1705, signal_1704, signal_1703, signal_1702, signal_434}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_420 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1225, signal_1224, signal_1223, signal_1222, signal_314}), .a ({signal_817, signal_816, signal_815, signal_814, signal_213}), .clk (clk), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .c ({signal_1709, signal_1708, signal_1707, signal_1706, signal_435}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_421 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1009, signal_1008, signal_1007, signal_1006, signal_260}), .a ({signal_833, signal_832, signal_831, signal_830, signal_217}), .clk (clk), .r ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_1713, signal_1712, signal_1711, signal_1710, signal_436}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_422 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_741, signal_740, signal_739, signal_738, signal_194}), .a ({signal_921, signal_920, signal_919, signal_918, signal_239}), .clk (clk), .r ({Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .c ({signal_1717, signal_1716, signal_1715, signal_1714, signal_437}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_423 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_809, signal_808, signal_807, signal_806, signal_211}), .a ({signal_797, signal_796, signal_795, signal_794, signal_208}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870]}), .c ({signal_1721, signal_1720, signal_1719, signal_1718, signal_438}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_424 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_997, signal_996, signal_995, signal_994, signal_257}), .a ({signal_805, signal_804, signal_803, signal_802, signal_210}), .clk (clk), .r ({Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_1725, signal_1724, signal_1723, signal_1722, signal_439}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_425 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_629, signal_628, signal_627, signal_626, signal_166}), .a ({signal_1149, signal_1148, signal_1147, signal_1146, signal_295}), .clk (clk), .r ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890]}), .c ({signal_1729, signal_1728, signal_1727, signal_1726, signal_440}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_426 ( .s ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_1197, signal_1196, signal_1195, signal_1194, signal_307}), .a ({signal_953, signal_952, signal_951, signal_950, signal_246}), .clk (clk), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .c ({signal_1733, signal_1732, signal_1731, signal_1730, signal_441}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_427 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1353, signal_1352, signal_1351, signal_1350, signal_346}), .a ({signal_1541, signal_1540, signal_1539, signal_1538, signal_393}), .clk (clk), .r ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_1741, signal_1740, signal_1739, signal_1738, signal_442}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_428 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1345, signal_1344, signal_1343, signal_1342, signal_344}), .a ({signal_1673, signal_1672, signal_1671, signal_1670, signal_426}), .clk (clk), .r ({Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .c ({signal_1745, signal_1744, signal_1743, signal_1742, signal_443}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_429 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1525, signal_1524, signal_1523, signal_1522, signal_389}), .a ({signal_1589, signal_1588, signal_1587, signal_1586, signal_405}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930]}), .c ({signal_1749, signal_1748, signal_1747, signal_1746, signal_444}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_430 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1425, signal_1424, signal_1423, signal_1422, signal_364}), .a ({signal_1713, signal_1712, signal_1711, signal_1710, signal_436}), .clk (clk), .r ({Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_1753, signal_1752, signal_1751, signal_1750, signal_445}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_431 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1701, signal_1700, signal_1699, signal_1698, signal_433}), .a ({signal_1665, signal_1664, signal_1663, signal_1662, signal_424}), .clk (clk), .r ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950]}), .c ({signal_1757, signal_1756, signal_1755, signal_1754, signal_446}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_432 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1317, signal_1316, signal_1315, signal_1314, signal_337}), .a ({signal_1501, signal_1500, signal_1499, signal_1498, signal_383}), .clk (clk), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .c ({signal_1761, signal_1760, signal_1759, signal_1758, signal_447}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_433 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1437, signal_1436, signal_1435, signal_1434, signal_367}), .a ({signal_1657, signal_1656, signal_1655, signal_1654, signal_422}), .clk (clk), .r ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_1765, signal_1764, signal_1763, signal_1762, signal_448}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_434 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1341, signal_1340, signal_1339, signal_1338, signal_343}), .a ({signal_1577, signal_1576, signal_1575, signal_1574, signal_402}), .clk (clk), .r ({Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .c ({signal_1769, signal_1768, signal_1767, signal_1766, signal_449}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_435 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1729, signal_1728, signal_1727, signal_1726, signal_440}), .a ({signal_1265, signal_1264, signal_1263, signal_1262, signal_324}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990]}), .c ({signal_1773, signal_1772, signal_1771, signal_1770, signal_450}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_436 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1405, signal_1404, signal_1403, signal_1402, signal_359}), .a ({signal_1733, signal_1732, signal_1731, signal_1730, signal_441}), .clk (clk), .r ({Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_1777, signal_1776, signal_1775, signal_1774, signal_451}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_437 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1397, signal_1396, signal_1395, signal_1394, signal_357}), .a ({signal_1497, signal_1496, signal_1495, signal_1494, signal_382}), .clk (clk), .r ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010]}), .c ({signal_1781, signal_1780, signal_1779, signal_1778, signal_452}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_438 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1537, signal_1536, signal_1535, signal_1534, signal_392}), .a ({signal_1513, signal_1512, signal_1511, signal_1510, signal_386}), .clk (clk), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .c ({signal_1785, signal_1784, signal_1783, signal_1782, signal_453}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_439 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1293, signal_1292, signal_1291, signal_1290, signal_331}), .a ({signal_1649, signal_1648, signal_1647, signal_1646, signal_420}), .clk (clk), .r ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_1789, signal_1788, signal_1787, signal_1786, signal_454}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_440 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1629, signal_1628, signal_1627, signal_1626, signal_415}), .a ({signal_1633, signal_1632, signal_1631, signal_1630, signal_416}), .clk (clk), .r ({Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .c ({signal_1793, signal_1792, signal_1791, signal_1790, signal_455}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_441 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1553, signal_1552, signal_1551, signal_1550, signal_396}), .a ({signal_1097, signal_1096, signal_1095, signal_1094, signal_282}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050]}), .c ({signal_1797, signal_1796, signal_1795, signal_1794, signal_456}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_442 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1709, signal_1708, signal_1707, signal_1706, signal_435}), .a ({signal_1645, signal_1644, signal_1643, signal_1642, signal_419}), .clk (clk), .r ({Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_1801, signal_1800, signal_1799, signal_1798, signal_457}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_443 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1261, signal_1260, signal_1259, signal_1258, signal_323}), .a ({signal_1361, signal_1360, signal_1359, signal_1358, signal_348}), .clk (clk), .r ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070]}), .c ({signal_1805, signal_1804, signal_1803, signal_1802, signal_458}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_444 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1565, signal_1564, signal_1563, signal_1562, signal_399}), .a ({signal_1065, signal_1064, signal_1063, signal_1062, signal_274}), .clk (clk), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .c ({signal_1809, signal_1808, signal_1807, signal_1806, signal_459}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_445 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1697, signal_1696, signal_1695, signal_1694, signal_432}), .a ({signal_1193, signal_1192, signal_1191, signal_1190, signal_306}), .clk (clk), .r ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_1813, signal_1812, signal_1811, signal_1810, signal_460}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_446 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1485, signal_1484, signal_1483, signal_1482, signal_379}), .a ({signal_1273, signal_1272, signal_1271, signal_1270, signal_326}), .clk (clk), .r ({Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .c ({signal_1817, signal_1816, signal_1815, signal_1814, signal_461}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_447 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1441, signal_1440, signal_1439, signal_1438, signal_368}), .a ({signal_1373, signal_1372, signal_1371, signal_1370, signal_351}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110]}), .c ({signal_1821, signal_1820, signal_1819, signal_1818, signal_462}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_448 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1305, signal_1304, signal_1303, signal_1302, signal_334}), .a ({signal_1465, signal_1464, signal_1463, signal_1462, signal_374}), .clk (clk), .r ({Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_1825, signal_1824, signal_1823, signal_1822, signal_463}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_449 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1617, signal_1616, signal_1615, signal_1614, signal_412}), .a ({signal_1269, signal_1268, signal_1267, signal_1266, signal_325}), .clk (clk), .r ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130]}), .c ({signal_1829, signal_1828, signal_1827, signal_1826, signal_464}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_450 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1413, signal_1412, signal_1411, signal_1410, signal_361}), .a ({signal_1573, signal_1572, signal_1571, signal_1570, signal_401}), .clk (clk), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .c ({signal_1833, signal_1832, signal_1831, signal_1830, signal_465}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_451 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1277, signal_1276, signal_1275, signal_1274, signal_327}), .a ({signal_1289, signal_1288, signal_1287, signal_1286, signal_330}), .clk (clk), .r ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_1837, signal_1836, signal_1835, signal_1834, signal_466}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_452 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1249, signal_1248, signal_1247, signal_1246, signal_320}), .a ({signal_1349, signal_1348, signal_1347, signal_1346, signal_345}), .clk (clk), .r ({Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .c ({signal_1841, signal_1840, signal_1839, signal_1838, signal_467}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_453 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1601, signal_1600, signal_1599, signal_1598, signal_408}), .a ({signal_1721, signal_1720, signal_1719, signal_1718, signal_438}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170]}), .c ({signal_1845, signal_1844, signal_1843, signal_1842, signal_468}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_454 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1689, signal_1688, signal_1687, signal_1686, signal_430}), .a ({signal_1637, signal_1636, signal_1635, signal_1634, signal_417}), .clk (clk), .r ({Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_1849, signal_1848, signal_1847, signal_1846, signal_469}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_455 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1625, signal_1624, signal_1623, signal_1622, signal_414}), .a ({signal_1329, signal_1328, signal_1327, signal_1326, signal_340}), .clk (clk), .r ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190]}), .c ({signal_1853, signal_1852, signal_1851, signal_1850, signal_470}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_456 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1453, signal_1452, signal_1451, signal_1450, signal_371}), .a ({signal_1165, signal_1164, signal_1163, signal_1162, signal_299}), .clk (clk), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .c ({signal_1857, signal_1856, signal_1855, signal_1854, signal_471}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_457 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1365, signal_1364, signal_1363, signal_1362, signal_349}), .a ({signal_1369, signal_1368, signal_1367, signal_1366, signal_350}), .clk (clk), .r ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_1861, signal_1860, signal_1859, signal_1858, signal_472}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_458 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1505, signal_1504, signal_1503, signal_1502, signal_384}), .a ({signal_1517, signal_1516, signal_1515, signal_1514, signal_387}), .clk (clk), .r ({Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .c ({signal_1865, signal_1864, signal_1863, signal_1862, signal_473}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_459 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1469, signal_1468, signal_1467, signal_1466, signal_375}), .a ({signal_1333, signal_1332, signal_1331, signal_1330, signal_341}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230]}), .c ({signal_1869, signal_1868, signal_1867, signal_1866, signal_474}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_460 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1521, signal_1520, signal_1519, signal_1518, signal_388}), .a ({signal_1609, signal_1608, signal_1607, signal_1606, signal_410}), .clk (clk), .r ({Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_1873, signal_1872, signal_1871, signal_1870, signal_475}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_461 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1409, signal_1408, signal_1407, signal_1406, signal_360}), .a ({signal_1509, signal_1508, signal_1507, signal_1506, signal_385}), .clk (clk), .r ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250]}), .c ({signal_1877, signal_1876, signal_1875, signal_1874, signal_476}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_462 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1717, signal_1716, signal_1715, signal_1714, signal_437}), .a ({signal_1325, signal_1324, signal_1323, signal_1322, signal_339}), .clk (clk), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .c ({signal_1881, signal_1880, signal_1879, signal_1878, signal_477}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_463 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1581, signal_1580, signal_1579, signal_1578, signal_403}), .a ({signal_1297, signal_1296, signal_1295, signal_1294, signal_332}), .clk (clk), .r ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_1885, signal_1884, signal_1883, signal_1882, signal_478}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_464 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1309, signal_1308, signal_1307, signal_1306, signal_335}), .a ({signal_1337, signal_1336, signal_1335, signal_1334, signal_342}), .clk (clk), .r ({Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .c ({signal_1889, signal_1888, signal_1887, signal_1886, signal_479}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_465 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1313, signal_1312, signal_1311, signal_1310, signal_336}), .a ({signal_1429, signal_1428, signal_1427, signal_1426, signal_365}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290]}), .c ({signal_1893, signal_1892, signal_1891, signal_1890, signal_480}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_466 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1393, signal_1392, signal_1391, signal_1390, signal_356}), .a ({signal_1681, signal_1680, signal_1679, signal_1678, signal_428}), .clk (clk), .r ({Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_1897, signal_1896, signal_1895, signal_1894, signal_481}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_467 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1445, signal_1444, signal_1443, signal_1442, signal_369}), .a ({signal_1481, signal_1480, signal_1479, signal_1478, signal_378}), .clk (clk), .r ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310]}), .c ({signal_1901, signal_1900, signal_1899, signal_1898, signal_482}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_468 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1533, signal_1532, signal_1531, signal_1530, signal_391}), .a ({signal_1557, signal_1556, signal_1555, signal_1554, signal_397}), .clk (clk), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .c ({signal_1905, signal_1904, signal_1903, signal_1902, signal_483}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_469 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1461, signal_1460, signal_1459, signal_1458, signal_373}), .a ({signal_1281, signal_1280, signal_1279, signal_1278, signal_328}), .clk (clk), .r ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_1909, signal_1908, signal_1907, signal_1906, signal_484}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_470 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1653, signal_1652, signal_1651, signal_1650, signal_421}), .a ({signal_1473, signal_1472, signal_1471, signal_1470, signal_376}), .clk (clk), .r ({Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .c ({signal_1913, signal_1912, signal_1911, signal_1910, signal_485}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_471 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1377, signal_1376, signal_1375, signal_1374, signal_352}), .a ({signal_1433, signal_1432, signal_1431, signal_1430, signal_366}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350]}), .c ({signal_1917, signal_1916, signal_1915, signal_1914, signal_486}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_472 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1693, signal_1692, signal_1691, signal_1690, signal_431}), .a ({signal_1641, signal_1640, signal_1639, signal_1638, signal_418}), .clk (clk), .r ({Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_1921, signal_1920, signal_1919, signal_1918, signal_487}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_473 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1561, signal_1560, signal_1559, signal_1558, signal_398}), .a ({signal_1669, signal_1668, signal_1667, signal_1666, signal_425}), .clk (clk), .r ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370]}), .c ({signal_1925, signal_1924, signal_1923, signal_1922, signal_488}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_474 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1385, signal_1384, signal_1383, signal_1382, signal_354}), .a ({signal_1613, signal_1612, signal_1611, signal_1610, signal_411}), .clk (clk), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .c ({signal_1929, signal_1928, signal_1927, signal_1926, signal_489}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_475 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1381, signal_1380, signal_1379, signal_1378, signal_353}), .a ({signal_1301, signal_1300, signal_1299, signal_1298, signal_333}), .clk (clk), .r ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_1933, signal_1932, signal_1931, signal_1930, signal_490}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_476 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1417, signal_1416, signal_1415, signal_1414, signal_362}), .a ({signal_1493, signal_1492, signal_1491, signal_1490, signal_381}), .clk (clk), .r ({Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .c ({signal_1937, signal_1936, signal_1935, signal_1934, signal_491}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_477 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1489, signal_1488, signal_1487, signal_1486, signal_380}), .a ({signal_1585, signal_1584, signal_1583, signal_1582, signal_404}), .clk (clk), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410]}), .c ({signal_1941, signal_1940, signal_1939, signal_1938, signal_492}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_478 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_945, signal_944, signal_943, signal_942, signal_244}), .a ({signal_1421, signal_1420, signal_1419, signal_1418, signal_363}), .clk (clk), .r ({Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_1945, signal_1944, signal_1943, signal_1942, signal_493}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_479 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1401, signal_1400, signal_1399, signal_1398, signal_358}), .a ({signal_1549, signal_1548, signal_1547, signal_1546, signal_395}), .clk (clk), .r ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430]}), .c ({signal_1949, signal_1948, signal_1947, signal_1946, signal_494}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_480 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1725, signal_1724, signal_1723, signal_1722, signal_439}), .a ({signal_1685, signal_1684, signal_1683, signal_1682, signal_429}), .clk (clk), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .c ({signal_1953, signal_1952, signal_1951, signal_1950, signal_495}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_481 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1597, signal_1596, signal_1595, signal_1594, signal_407}), .a ({signal_1257, signal_1256, signal_1255, signal_1254, signal_322}), .clk (clk), .r ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_1957, signal_1956, signal_1955, signal_1954, signal_496}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_482 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1389, signal_1388, signal_1387, signal_1386, signal_355}), .a ({signal_1705, signal_1704, signal_1703, signal_1702, signal_434}), .clk (clk), .r ({Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .c ({signal_1961, signal_1960, signal_1959, signal_1958, signal_497}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_483 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1529, signal_1528, signal_1527, signal_1526, signal_390}), .a ({signal_1605, signal_1604, signal_1603, signal_1602, signal_409}), .clk (clk), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470]}), .c ({signal_1965, signal_1964, signal_1963, signal_1962, signal_498}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_484 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1285, signal_1284, signal_1283, signal_1282, signal_329}), .a ({signal_1477, signal_1476, signal_1475, signal_1474, signal_377}), .clk (clk), .r ({Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_1969, signal_1968, signal_1967, signal_1966, signal_499}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_485 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1253, signal_1252, signal_1251, signal_1250, signal_321}), .a ({signal_1661, signal_1660, signal_1659, signal_1658, signal_423}), .clk (clk), .r ({Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490]}), .c ({signal_1973, signal_1972, signal_1971, signal_1970, signal_500}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_486 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1621, signal_1620, signal_1619, signal_1618, signal_413}), .a ({signal_1569, signal_1568, signal_1567, signal_1566, signal_400}), .clk (clk), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500]}), .c ({signal_1977, signal_1976, signal_1975, signal_1974, signal_501}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_487 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1457, signal_1456, signal_1455, signal_1454, signal_372}), .a ({signal_1593, signal_1592, signal_1591, signal_1590, signal_406}), .clk (clk), .r ({Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_1981, signal_1980, signal_1979, signal_1978, signal_502}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_488 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1177, signal_1176, signal_1175, signal_1174, signal_302}), .a ({signal_1677, signal_1676, signal_1675, signal_1674, signal_427}), .clk (clk), .r ({Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520]}), .c ({signal_1985, signal_1984, signal_1983, signal_1982, signal_503}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_489 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1449, signal_1448, signal_1447, signal_1446, signal_370}), .a ({signal_1357, signal_1356, signal_1355, signal_1354, signal_347}), .clk (clk), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530]}), .c ({signal_1989, signal_1988, signal_1987, signal_1986, signal_504}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_490 ( .s ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_1545, signal_1544, signal_1543, signal_1542, signal_394}), .a ({signal_1321, signal_1320, signal_1319, signal_1318, signal_338}), .clk (clk), .r ({Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_1993, signal_1992, signal_1991, signal_1990, signal_505}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_491 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1873, signal_1872, signal_1871, signal_1870, signal_475}), .a ({signal_1749, signal_1748, signal_1747, signal_1746, signal_444}), .clk (clk), .r ({Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550]}), .c ({signal_2001, signal_2000, signal_1999, signal_1998, signal_506}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_492 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1773, signal_1772, signal_1771, signal_1770, signal_450}), .a ({signal_1793, signal_1792, signal_1791, signal_1790, signal_455}), .clk (clk), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560]}), .c ({signal_2005, signal_2004, signal_2003, signal_2002, signal_507}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_493 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1929, signal_1928, signal_1927, signal_1926, signal_489}), .a ({signal_1853, signal_1852, signal_1851, signal_1850, signal_470}), .clk (clk), .r ({Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_2009, signal_2008, signal_2007, signal_2006, signal_508}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_494 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1905, signal_1904, signal_1903, signal_1902, signal_483}), .a ({signal_1753, signal_1752, signal_1751, signal_1750, signal_445}), .clk (clk), .r ({Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580]}), .c ({signal_2013, signal_2012, signal_2011, signal_2010, signal_509}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_495 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1969, signal_1968, signal_1967, signal_1966, signal_499}), .a ({signal_1801, signal_1800, signal_1799, signal_1798, signal_457}), .clk (clk), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590]}), .c ({signal_2017, signal_2016, signal_2015, signal_2014, signal_510}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_496 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1893, signal_1892, signal_1891, signal_1890, signal_480}), .a ({signal_1885, signal_1884, signal_1883, signal_1882, signal_478}), .clk (clk), .r ({Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_2021, signal_2020, signal_2019, signal_2018, signal_511}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_497 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1977, signal_1976, signal_1975, signal_1974, signal_501}), .a ({signal_1877, signal_1876, signal_1875, signal_1874, signal_476}), .clk (clk), .r ({Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610]}), .c ({signal_2025, signal_2024, signal_2023, signal_2022, signal_512}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_498 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1933, signal_1932, signal_1931, signal_1930, signal_490}), .a ({signal_1845, signal_1844, signal_1843, signal_1842, signal_468}), .clk (clk), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620]}), .c ({signal_2029, signal_2028, signal_2027, signal_2026, signal_513}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_499 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1985, signal_1984, signal_1983, signal_1982, signal_503}), .a ({signal_1817, signal_1816, signal_1815, signal_1814, signal_461}), .clk (clk), .r ({Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_2033, signal_2032, signal_2031, signal_2030, signal_514}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_500 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1805, signal_1804, signal_1803, signal_1802, signal_458}), .a ({signal_1821, signal_1820, signal_1819, signal_1818, signal_462}), .clk (clk), .r ({Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640]}), .c ({signal_2037, signal_2036, signal_2035, signal_2034, signal_515}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_501 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1769, signal_1768, signal_1767, signal_1766, signal_449}), .a ({signal_1841, signal_1840, signal_1839, signal_1838, signal_467}), .clk (clk), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650]}), .c ({signal_2041, signal_2040, signal_2039, signal_2038, signal_516}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_502 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1965, signal_1964, signal_1963, signal_1962, signal_498}), .a ({signal_1937, signal_1936, signal_1935, signal_1934, signal_491}), .clk (clk), .r ({Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_2045, signal_2044, signal_2043, signal_2042, signal_517}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_503 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1781, signal_1780, signal_1779, signal_1778, signal_452}), .a ({signal_1925, signal_1924, signal_1923, signal_1922, signal_488}), .clk (clk), .r ({Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670]}), .c ({signal_2049, signal_2048, signal_2047, signal_2046, signal_518}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_504 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1941, signal_1940, signal_1939, signal_1938, signal_492}), .a ({signal_1849, signal_1848, signal_1847, signal_1846, signal_469}), .clk (clk), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680]}), .c ({signal_2053, signal_2052, signal_2051, signal_2050, signal_519}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_505 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1953, signal_1952, signal_1951, signal_1950, signal_495}), .a ({signal_1861, signal_1860, signal_1859, signal_1858, signal_472}), .clk (clk), .r ({Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_2057, signal_2056, signal_2055, signal_2054, signal_520}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_506 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1957, signal_1956, signal_1955, signal_1954, signal_496}), .a ({signal_1829, signal_1828, signal_1827, signal_1826, signal_464}), .clk (clk), .r ({Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700]}), .c ({signal_2061, signal_2060, signal_2059, signal_2058, signal_521}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_507 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1949, signal_1948, signal_1947, signal_1946, signal_494}), .a ({signal_1813, signal_1812, signal_1811, signal_1810, signal_460}), .clk (clk), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710]}), .c ({signal_2065, signal_2064, signal_2063, signal_2062, signal_522}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_508 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1865, signal_1864, signal_1863, signal_1862, signal_473}), .a ({signal_1961, signal_1960, signal_1959, signal_1958, signal_497}), .clk (clk), .r ({Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_2069, signal_2068, signal_2067, signal_2066, signal_523}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_509 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1945, signal_1944, signal_1943, signal_1942, signal_493}), .a ({signal_1809, signal_1808, signal_1807, signal_1806, signal_459}), .clk (clk), .r ({Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730]}), .c ({signal_2073, signal_2072, signal_2071, signal_2070, signal_524}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_510 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1789, signal_1788, signal_1787, signal_1786, signal_454}), .a ({signal_1981, signal_1980, signal_1979, signal_1978, signal_502}), .clk (clk), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740]}), .c ({signal_2077, signal_2076, signal_2075, signal_2074, signal_525}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_511 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1989, signal_1988, signal_1987, signal_1986, signal_504}), .a ({signal_1889, signal_1888, signal_1887, signal_1886, signal_479}), .clk (clk), .r ({Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_2081, signal_2080, signal_2079, signal_2078, signal_526}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_512 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1797, signal_1796, signal_1795, signal_1794, signal_456}), .a ({signal_1761, signal_1760, signal_1759, signal_1758, signal_447}), .clk (clk), .r ({Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760]}), .c ({signal_2085, signal_2084, signal_2083, signal_2082, signal_527}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_513 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1757, signal_1756, signal_1755, signal_1754, signal_446}), .a ({signal_1837, signal_1836, signal_1835, signal_1834, signal_466}), .clk (clk), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770]}), .c ({signal_2089, signal_2088, signal_2087, signal_2086, signal_528}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_514 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1857, signal_1856, signal_1855, signal_1854, signal_471}), .a ({signal_1913, signal_1912, signal_1911, signal_1910, signal_485}), .clk (clk), .r ({Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_2093, signal_2092, signal_2091, signal_2090, signal_529}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_515 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1901, signal_1900, signal_1899, signal_1898, signal_482}), .a ({signal_1777, signal_1776, signal_1775, signal_1774, signal_451}), .clk (clk), .r ({Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790]}), .c ({signal_2097, signal_2096, signal_2095, signal_2094, signal_530}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_516 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1765, signal_1764, signal_1763, signal_1762, signal_448}), .a ({signal_1825, signal_1824, signal_1823, signal_1822, signal_463}), .clk (clk), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800]}), .c ({signal_2101, signal_2100, signal_2099, signal_2098, signal_531}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_517 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1833, signal_1832, signal_1831, signal_1830, signal_465}), .a ({signal_1993, signal_1992, signal_1991, signal_1990, signal_505}), .clk (clk), .r ({Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_2105, signal_2104, signal_2103, signal_2102, signal_532}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_518 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1785, signal_1784, signal_1783, signal_1782, signal_453}), .a ({signal_1973, signal_1972, signal_1971, signal_1970, signal_500}), .clk (clk), .r ({Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820]}), .c ({signal_2109, signal_2108, signal_2107, signal_2106, signal_533}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_519 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1869, signal_1868, signal_1867, signal_1866, signal_474}), .a ({signal_1897, signal_1896, signal_1895, signal_1894, signal_481}), .clk (clk), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830]}), .c ({signal_2113, signal_2112, signal_2111, signal_2110, signal_534}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_520 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1881, signal_1880, signal_1879, signal_1878, signal_477}), .a ({signal_1909, signal_1908, signal_1907, signal_1906, signal_484}), .clk (clk), .r ({Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_2117, signal_2116, signal_2115, signal_2114, signal_535}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_521 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1921, signal_1920, signal_1919, signal_1918, signal_487}), .a ({signal_1741, signal_1740, signal_1739, signal_1738, signal_442}), .clk (clk), .r ({Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850]}), .c ({signal_2121, signal_2120, signal_2119, signal_2118, signal_536}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_522 ( .s ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_1917, signal_1916, signal_1915, signal_1914, signal_486}), .a ({signal_1745, signal_1744, signal_1743, signal_1742, signal_443}), .clk (clk), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860]}), .c ({signal_2125, signal_2124, signal_2123, signal_2122, signal_537}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_523 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2101, signal_2100, signal_2099, signal_2098, signal_531}), .a ({signal_2049, signal_2048, signal_2047, signal_2046, signal_518}), .clk (clk), .r ({Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_2133, signal_2132, signal_2131, signal_2130, signal_538}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_524 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2009, signal_2008, signal_2007, signal_2006, signal_508}), .a ({signal_2117, signal_2116, signal_2115, signal_2114, signal_535}), .clk (clk), .r ({Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880]}), .c ({signal_2137, signal_2136, signal_2135, signal_2134, signal_539}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_525 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2073, signal_2072, signal_2071, signal_2070, signal_524}), .a ({signal_2069, signal_2068, signal_2067, signal_2066, signal_523}), .clk (clk), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890]}), .c ({signal_2141, signal_2140, signal_2139, signal_2138, signal_540}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_526 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2053, signal_2052, signal_2051, signal_2050, signal_519}), .a ({signal_2085, signal_2084, signal_2083, signal_2082, signal_527}), .clk (clk), .r ({Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_2145, signal_2144, signal_2143, signal_2142, signal_541}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_527 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2089, signal_2088, signal_2087, signal_2086, signal_528}), .a ({signal_2001, signal_2000, signal_1999, signal_1998, signal_506}), .clk (clk), .r ({Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910]}), .c ({signal_2149, signal_2148, signal_2147, signal_2146, signal_542}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_528 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2081, signal_2080, signal_2079, signal_2078, signal_526}), .a ({signal_2125, signal_2124, signal_2123, signal_2122, signal_537}), .clk (clk), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920]}), .c ({signal_2153, signal_2152, signal_2151, signal_2150, signal_543}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_529 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2017, signal_2016, signal_2015, signal_2014, signal_510}), .a ({signal_2109, signal_2108, signal_2107, signal_2106, signal_533}), .clk (clk), .r ({Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_2157, signal_2156, signal_2155, signal_2154, signal_544}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_530 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2005, signal_2004, signal_2003, signal_2002, signal_507}), .a ({signal_2021, signal_2020, signal_2019, signal_2018, signal_511}), .clk (clk), .r ({Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940]}), .c ({signal_2161, signal_2160, signal_2159, signal_2158, signal_545}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_531 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2033, signal_2032, signal_2031, signal_2030, signal_514}), .a ({signal_2041, signal_2040, signal_2039, signal_2038, signal_516}), .clk (clk), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950]}), .c ({signal_2165, signal_2164, signal_2163, signal_2162, signal_546}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_532 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2057, signal_2056, signal_2055, signal_2054, signal_520}), .a ({signal_2077, signal_2076, signal_2075, signal_2074, signal_525}), .clk (clk), .r ({Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_2169, signal_2168, signal_2167, signal_2166, signal_547}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_533 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2025, signal_2024, signal_2023, signal_2022, signal_512}), .a ({signal_2097, signal_2096, signal_2095, signal_2094, signal_530}), .clk (clk), .r ({Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970]}), .c ({signal_2173, signal_2172, signal_2171, signal_2170, signal_548}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_534 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2037, signal_2036, signal_2035, signal_2034, signal_515}), .a ({signal_2113, signal_2112, signal_2111, signal_2110, signal_534}), .clk (clk), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980]}), .c ({signal_2177, signal_2176, signal_2175, signal_2174, signal_549}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_535 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2061, signal_2060, signal_2059, signal_2058, signal_521}), .a ({signal_2045, signal_2044, signal_2043, signal_2042, signal_517}), .clk (clk), .r ({Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_2181, signal_2180, signal_2179, signal_2178, signal_550}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_536 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2093, signal_2092, signal_2091, signal_2090, signal_529}), .a ({signal_2121, signal_2120, signal_2119, signal_2118, signal_536}), .clk (clk), .r ({Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000]}), .c ({signal_2185, signal_2184, signal_2183, signal_2182, signal_551}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_537 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2029, signal_2028, signal_2027, signal_2026, signal_513}), .a ({signal_2105, signal_2104, signal_2103, signal_2102, signal_532}), .clk (clk), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010]}), .c ({signal_2189, signal_2188, signal_2187, signal_2186, signal_552}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_538 ( .s ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_2013, signal_2012, signal_2011, signal_2010, signal_509}), .a ({signal_2065, signal_2064, signal_2063, signal_2062, signal_522}), .clk (clk), .r ({Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_2193, signal_2192, signal_2191, signal_2190, signal_553}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_539 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2137, signal_2136, signal_2135, signal_2134, signal_539}), .a ({signal_2161, signal_2160, signal_2159, signal_2158, signal_545}), .clk (clk), .r ({Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030]}), .c ({signal_2201, signal_2200, signal_2199, signal_2198, signal_145}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_540 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2173, signal_2172, signal_2171, signal_2170, signal_548}), .a ({signal_2165, signal_2164, signal_2163, signal_2162, signal_546}), .clk (clk), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040]}), .c ({signal_2205, signal_2204, signal_2203, signal_2202, signal_148}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_541 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2153, signal_2152, signal_2151, signal_2150, signal_543}), .a ({signal_2169, signal_2168, signal_2167, signal_2166, signal_547}), .clk (clk), .r ({Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_2209, signal_2208, signal_2207, signal_2206, signal_143}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_542 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2193, signal_2192, signal_2191, signal_2190, signal_553}), .a ({signal_2185, signal_2184, signal_2183, signal_2182, signal_551}), .clk (clk), .r ({Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060]}), .c ({signal_2213, signal_2212, signal_2211, signal_2210, signal_146}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_543 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2141, signal_2140, signal_2139, signal_2138, signal_540}), .a ({signal_2189, signal_2188, signal_2187, signal_2186, signal_552}), .clk (clk), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070]}), .c ({signal_2217, signal_2216, signal_2215, signal_2214, signal_149}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_544 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2181, signal_2180, signal_2179, signal_2178, signal_550}), .a ({signal_2149, signal_2148, signal_2147, signal_2146, signal_542}), .clk (clk), .r ({Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_2221, signal_2220, signal_2219, signal_2218, signal_144}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_545 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2133, signal_2132, signal_2131, signal_2130, signal_538}), .a ({signal_2177, signal_2176, signal_2175, signal_2174, signal_549}), .clk (clk), .r ({Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090]}), .c ({signal_2225, signal_2224, signal_2223, signal_2222, signal_147}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_546 ( .s ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_2157, signal_2156, signal_2155, signal_2154, signal_544}), .a ({signal_2145, signal_2144, signal_2143, signal_2142, signal_541}), .clk (clk), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100]}), .c ({signal_2229, signal_2228, signal_2227, signal_2226, signal_150}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(0)) cell_0 ( .clk (signal_6373), .D ({signal_2209, signal_2208, signal_2207, signal_2206, signal_143}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_1 ( .clk (signal_6373), .D ({signal_2221, signal_2220, signal_2219, signal_2218, signal_144}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_2 ( .clk (signal_6373), .D ({signal_2201, signal_2200, signal_2199, signal_2198, signal_145}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_3 ( .clk (signal_6373), .D ({signal_2213, signal_2212, signal_2211, signal_2210, signal_146}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_4 ( .clk (signal_6373), .D ({signal_2225, signal_2224, signal_2223, signal_2222, signal_147}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_5 ( .clk (signal_6373), .D ({signal_2205, signal_2204, signal_2203, signal_2202, signal_148}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_6 ( .clk (signal_6373), .D ({signal_2217, signal_2216, signal_2215, signal_2214, signal_149}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_7 ( .clk (signal_6373), .D ({signal_2229, signal_2228, signal_2227, signal_2226, signal_150}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
