/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [3:0] X_s3 ;
    input [23:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    output [3:0] Y_s3 ;
    wire signal_33 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_66 ;
    wire signal_67 ;
    wire signal_68 ;
    wire signal_72 ;
    wire signal_73 ;
    wire signal_74 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_83 ;
    wire signal_84 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) cell_26 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_62, signal_61, signal_60, signal_37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_27 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_68, signal_67, signal_66, signal_38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_28 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_74, signal_73, signal_72, signal_39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_29 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_80, signal_79, signal_78, signal_40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_31 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_74, signal_73, signal_72, signal_39}), .c ({signal_86, signal_85, signal_84, signal_42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_32 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_68, signal_67, signal_66, signal_38}), .c ({signal_89, signal_88, signal_87, signal_43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_33 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_74, signal_73, signal_72, signal_39}), .c ({signal_92, signal_91, signal_90, signal_44}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_34 ( .a ({signal_92, signal_91, signal_90, signal_44}), .b ({signal_95, signal_94, signal_93, signal_45}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_36 ( .a ({signal_89, signal_88, signal_87, signal_43}), .b ({signal_92, signal_91, signal_90, signal_44}), .c ({signal_101, signal_100, signal_99, signal_47}) ) ;

    /* cells in depth 1 */
    buf_clk cell_50 ( .C (clk), .D (signal_38), .Q (signal_177) ) ;
    buf_clk cell_52 ( .C (clk), .D (signal_66), .Q (signal_179) ) ;
    buf_clk cell_54 ( .C (clk), .D (signal_67), .Q (signal_181) ) ;
    buf_clk cell_56 ( .C (clk), .D (signal_68), .Q (signal_183) ) ;
    buf_clk cell_58 ( .C (clk), .D (signal_42), .Q (signal_185) ) ;
    buf_clk cell_60 ( .C (clk), .D (signal_84), .Q (signal_187) ) ;
    buf_clk cell_62 ( .C (clk), .D (signal_85), .Q (signal_189) ) ;
    buf_clk cell_64 ( .C (clk), .D (signal_86), .Q (signal_191) ) ;
    buf_clk cell_66 ( .C (clk), .D (signal_47), .Q (signal_193) ) ;
    buf_clk cell_68 ( .C (clk), .D (signal_99), .Q (signal_195) ) ;
    buf_clk cell_70 ( .C (clk), .D (signal_100), .Q (signal_197) ) ;
    buf_clk cell_72 ( .C (clk), .D (signal_101), .Q (signal_199) ) ;
    buf_clk cell_74 ( .C (clk), .D (signal_39), .Q (signal_201) ) ;
    buf_clk cell_76 ( .C (clk), .D (signal_72), .Q (signal_203) ) ;
    buf_clk cell_78 ( .C (clk), .D (signal_73), .Q (signal_205) ) ;
    buf_clk cell_80 ( .C (clk), .D (signal_74), .Q (signal_207) ) ;
    buf_clk cell_82 ( .C (clk), .D (X_s0[1]), .Q (signal_209) ) ;
    buf_clk cell_84 ( .C (clk), .D (X_s1[1]), .Q (signal_211) ) ;
    buf_clk cell_86 ( .C (clk), .D (X_s2[1]), .Q (signal_213) ) ;
    buf_clk cell_88 ( .C (clk), .D (X_s3[1]), .Q (signal_215) ) ;
    buf_clk cell_90 ( .C (clk), .D (signal_45), .Q (signal_217) ) ;
    buf_clk cell_92 ( .C (clk), .D (signal_93), .Q (signal_219) ) ;
    buf_clk cell_94 ( .C (clk), .D (signal_94), .Q (signal_221) ) ;
    buf_clk cell_96 ( .C (clk), .D (signal_95), .Q (signal_223) ) ;
    buf_clk cell_106 ( .C (clk), .D (signal_40), .Q (signal_233) ) ;
    buf_clk cell_110 ( .C (clk), .D (signal_78), .Q (signal_237) ) ;
    buf_clk cell_114 ( .C (clk), .D (signal_79), .Q (signal_241) ) ;
    buf_clk cell_118 ( .C (clk), .D (signal_80), .Q (signal_245) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_30 ( .a ({signal_62, signal_61, signal_60, signal_37}), .b ({signal_80, signal_79, signal_78, signal_40}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_83, signal_82, signal_81, signal_41}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_35 ( .a ({signal_62, signal_61, signal_60, signal_37}), .b ({signal_89, signal_88, signal_87, signal_43}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_98, signal_97, signal_96, signal_46}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_37 ( .a ({signal_184, signal_182, signal_180, signal_178}), .b ({signal_83, signal_82, signal_81, signal_41}), .c ({signal_104, signal_103, signal_102, signal_48}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_38 ( .a ({signal_104, signal_103, signal_102, signal_48}), .b ({signal_107, signal_106, signal_105, signal_36}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_39 ( .a ({signal_192, signal_190, signal_188, signal_186}), .b ({signal_98, signal_97, signal_96, signal_46}), .c ({signal_110, signal_109, signal_108, signal_49}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_40 ( .a ({signal_83, signal_82, signal_81, signal_41}), .b ({signal_200, signal_198, signal_196, signal_194}), .c ({signal_113, signal_112, signal_111, signal_50}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_41 ( .a ({signal_208, signal_206, signal_204, signal_202}), .b ({signal_98, signal_97, signal_96, signal_46}), .c ({signal_116, signal_115, signal_114, signal_51}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_44 ( .a ({signal_83, signal_82, signal_81, signal_41}), .b ({signal_116, signal_115, signal_114, signal_51}), .c ({signal_125, signal_124, signal_123, signal_54}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_45 ( .a ({signal_125, signal_124, signal_123, signal_54}), .b ({signal_128, signal_127, signal_126, signal_35}) ) ;
    buf_clk cell_51 ( .C (clk), .D (signal_177), .Q (signal_178) ) ;
    buf_clk cell_53 ( .C (clk), .D (signal_179), .Q (signal_180) ) ;
    buf_clk cell_55 ( .C (clk), .D (signal_181), .Q (signal_182) ) ;
    buf_clk cell_57 ( .C (clk), .D (signal_183), .Q (signal_184) ) ;
    buf_clk cell_59 ( .C (clk), .D (signal_185), .Q (signal_186) ) ;
    buf_clk cell_61 ( .C (clk), .D (signal_187), .Q (signal_188) ) ;
    buf_clk cell_63 ( .C (clk), .D (signal_189), .Q (signal_190) ) ;
    buf_clk cell_65 ( .C (clk), .D (signal_191), .Q (signal_192) ) ;
    buf_clk cell_67 ( .C (clk), .D (signal_193), .Q (signal_194) ) ;
    buf_clk cell_69 ( .C (clk), .D (signal_195), .Q (signal_196) ) ;
    buf_clk cell_71 ( .C (clk), .D (signal_197), .Q (signal_198) ) ;
    buf_clk cell_73 ( .C (clk), .D (signal_199), .Q (signal_200) ) ;
    buf_clk cell_75 ( .C (clk), .D (signal_201), .Q (signal_202) ) ;
    buf_clk cell_77 ( .C (clk), .D (signal_203), .Q (signal_204) ) ;
    buf_clk cell_79 ( .C (clk), .D (signal_205), .Q (signal_206) ) ;
    buf_clk cell_81 ( .C (clk), .D (signal_207), .Q (signal_208) ) ;
    buf_clk cell_83 ( .C (clk), .D (signal_209), .Q (signal_210) ) ;
    buf_clk cell_85 ( .C (clk), .D (signal_211), .Q (signal_212) ) ;
    buf_clk cell_87 ( .C (clk), .D (signal_213), .Q (signal_214) ) ;
    buf_clk cell_89 ( .C (clk), .D (signal_215), .Q (signal_216) ) ;
    buf_clk cell_91 ( .C (clk), .D (signal_217), .Q (signal_218) ) ;
    buf_clk cell_93 ( .C (clk), .D (signal_219), .Q (signal_220) ) ;
    buf_clk cell_95 ( .C (clk), .D (signal_221), .Q (signal_222) ) ;
    buf_clk cell_97 ( .C (clk), .D (signal_223), .Q (signal_224) ) ;
    buf_clk cell_107 ( .C (clk), .D (signal_233), .Q (signal_234) ) ;
    buf_clk cell_111 ( .C (clk), .D (signal_237), .Q (signal_238) ) ;
    buf_clk cell_115 ( .C (clk), .D (signal_241), .Q (signal_242) ) ;
    buf_clk cell_119 ( .C (clk), .D (signal_245), .Q (signal_246) ) ;

    /* cells in depth 3 */
    buf_clk cell_98 ( .C (clk), .D (signal_41), .Q (signal_225) ) ;
    buf_clk cell_100 ( .C (clk), .D (signal_81), .Q (signal_227) ) ;
    buf_clk cell_102 ( .C (clk), .D (signal_82), .Q (signal_229) ) ;
    buf_clk cell_104 ( .C (clk), .D (signal_83), .Q (signal_231) ) ;
    buf_clk cell_108 ( .C (clk), .D (signal_234), .Q (signal_235) ) ;
    buf_clk cell_112 ( .C (clk), .D (signal_238), .Q (signal_239) ) ;
    buf_clk cell_116 ( .C (clk), .D (signal_242), .Q (signal_243) ) ;
    buf_clk cell_120 ( .C (clk), .D (signal_246), .Q (signal_247) ) ;
    buf_clk cell_122 ( .C (clk), .D (signal_51), .Q (signal_249) ) ;
    buf_clk cell_124 ( .C (clk), .D (signal_114), .Q (signal_251) ) ;
    buf_clk cell_126 ( .C (clk), .D (signal_115), .Q (signal_253) ) ;
    buf_clk cell_128 ( .C (clk), .D (signal_116), .Q (signal_255) ) ;
    buf_clk cell_130 ( .C (clk), .D (signal_35), .Q (signal_257) ) ;
    buf_clk cell_132 ( .C (clk), .D (signal_126), .Q (signal_259) ) ;
    buf_clk cell_134 ( .C (clk), .D (signal_127), .Q (signal_261) ) ;
    buf_clk cell_136 ( .C (clk), .D (signal_128), .Q (signal_263) ) ;
    buf_clk cell_138 ( .C (clk), .D (signal_36), .Q (signal_265) ) ;
    buf_clk cell_140 ( .C (clk), .D (signal_105), .Q (signal_267) ) ;
    buf_clk cell_142 ( .C (clk), .D (signal_106), .Q (signal_269) ) ;
    buf_clk cell_144 ( .C (clk), .D (signal_107), .Q (signal_271) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_42 ( .a ({signal_216, signal_214, signal_212, signal_210}), .b ({signal_110, signal_109, signal_108, signal_49}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_119, signal_118, signal_117, signal_52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_43 ( .a ({signal_224, signal_222, signal_220, signal_218}), .b ({signal_113, signal_112, signal_111, signal_50}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_122, signal_121, signal_120, signal_53}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_46 ( .a ({signal_232, signal_230, signal_228, signal_226}), .b ({signal_119, signal_118, signal_117, signal_52}), .c ({signal_131, signal_130, signal_129, signal_55}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_47 ( .a ({signal_248, signal_244, signal_240, signal_236}), .b ({signal_119, signal_118, signal_117, signal_52}), .c ({signal_134, signal_133, signal_132, signal_56}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_48 ( .a ({signal_256, signal_254, signal_252, signal_250}), .b ({signal_134, signal_133, signal_132, signal_56}), .c ({signal_137, signal_136, signal_135, signal_33}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_49 ( .a ({signal_122, signal_121, signal_120, signal_53}), .b ({signal_131, signal_130, signal_129, signal_55}), .c ({signal_140, signal_139, signal_138, signal_34}) ) ;
    buf_clk cell_99 ( .C (clk), .D (signal_225), .Q (signal_226) ) ;
    buf_clk cell_101 ( .C (clk), .D (signal_227), .Q (signal_228) ) ;
    buf_clk cell_103 ( .C (clk), .D (signal_229), .Q (signal_230) ) ;
    buf_clk cell_105 ( .C (clk), .D (signal_231), .Q (signal_232) ) ;
    buf_clk cell_109 ( .C (clk), .D (signal_235), .Q (signal_236) ) ;
    buf_clk cell_113 ( .C (clk), .D (signal_239), .Q (signal_240) ) ;
    buf_clk cell_117 ( .C (clk), .D (signal_243), .Q (signal_244) ) ;
    buf_clk cell_121 ( .C (clk), .D (signal_247), .Q (signal_248) ) ;
    buf_clk cell_123 ( .C (clk), .D (signal_249), .Q (signal_250) ) ;
    buf_clk cell_125 ( .C (clk), .D (signal_251), .Q (signal_252) ) ;
    buf_clk cell_127 ( .C (clk), .D (signal_253), .Q (signal_254) ) ;
    buf_clk cell_129 ( .C (clk), .D (signal_255), .Q (signal_256) ) ;
    buf_clk cell_131 ( .C (clk), .D (signal_257), .Q (signal_258) ) ;
    buf_clk cell_133 ( .C (clk), .D (signal_259), .Q (signal_260) ) ;
    buf_clk cell_135 ( .C (clk), .D (signal_261), .Q (signal_262) ) ;
    buf_clk cell_137 ( .C (clk), .D (signal_263), .Q (signal_264) ) ;
    buf_clk cell_139 ( .C (clk), .D (signal_265), .Q (signal_266) ) ;
    buf_clk cell_141 ( .C (clk), .D (signal_267), .Q (signal_268) ) ;
    buf_clk cell_143 ( .C (clk), .D (signal_269), .Q (signal_270) ) ;
    buf_clk cell_145 ( .C (clk), .D (signal_271), .Q (signal_272) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_264, signal_262, signal_260, signal_258}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_272, signal_270, signal_268, signal_266}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_137, signal_136, signal_135, signal_33}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_140, signal_139, signal_138, signal_34}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
