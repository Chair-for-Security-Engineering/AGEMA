/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d2 (SI_s0, clk, SI_s1, SI_s2, Fresh, SO_s0, SO_s1, SO_s2);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [2636:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;
    wire signal_8952 ;
    wire signal_8953 ;
    wire signal_8954 ;
    wire signal_8955 ;
    wire signal_8956 ;
    wire signal_8957 ;
    wire signal_8958 ;
    wire signal_8959 ;
    wire signal_8960 ;
    wire signal_8961 ;
    wire signal_8962 ;
    wire signal_8963 ;
    wire signal_8964 ;
    wire signal_8965 ;
    wire signal_8966 ;
    wire signal_8967 ;
    wire signal_8968 ;
    wire signal_8969 ;
    wire signal_8970 ;
    wire signal_8971 ;
    wire signal_8972 ;
    wire signal_8973 ;
    wire signal_8974 ;
    wire signal_8975 ;
    wire signal_8976 ;
    wire signal_8977 ;
    wire signal_8978 ;
    wire signal_8979 ;
    wire signal_8980 ;
    wire signal_8981 ;
    wire signal_8982 ;
    wire signal_8983 ;
    wire signal_8984 ;
    wire signal_8985 ;
    wire signal_8986 ;
    wire signal_8987 ;
    wire signal_8988 ;
    wire signal_8989 ;
    wire signal_8990 ;
    wire signal_8991 ;
    wire signal_8992 ;
    wire signal_8993 ;
    wire signal_8994 ;
    wire signal_8995 ;
    wire signal_8996 ;
    wire signal_8997 ;
    wire signal_8998 ;
    wire signal_8999 ;
    wire signal_9000 ;
    wire signal_9001 ;
    wire signal_9002 ;
    wire signal_9003 ;
    wire signal_9004 ;
    wire signal_9005 ;
    wire signal_9006 ;
    wire signal_9007 ;
    wire signal_9008 ;
    wire signal_9009 ;
    wire signal_9010 ;
    wire signal_9011 ;
    wire signal_9012 ;
    wire signal_9013 ;
    wire signal_9014 ;
    wire signal_9015 ;
    wire signal_9016 ;
    wire signal_9017 ;
    wire signal_9018 ;
    wire signal_9019 ;
    wire signal_9020 ;
    wire signal_9021 ;
    wire signal_9022 ;
    wire signal_9023 ;
    wire signal_9024 ;
    wire signal_9025 ;
    wire signal_9026 ;
    wire signal_9027 ;
    wire signal_9028 ;
    wire signal_9029 ;
    wire signal_9030 ;
    wire signal_9031 ;
    wire signal_9032 ;
    wire signal_9033 ;
    wire signal_9034 ;
    wire signal_9035 ;
    wire signal_9036 ;
    wire signal_9037 ;
    wire signal_9038 ;
    wire signal_9039 ;
    wire signal_9040 ;
    wire signal_9041 ;
    wire signal_9042 ;
    wire signal_9043 ;
    wire signal_9044 ;
    wire signal_9045 ;
    wire signal_9046 ;
    wire signal_9047 ;
    wire signal_9048 ;
    wire signal_9049 ;
    wire signal_9050 ;
    wire signal_9051 ;
    wire signal_9052 ;
    wire signal_9053 ;
    wire signal_9054 ;
    wire signal_9055 ;
    wire signal_9056 ;
    wire signal_9057 ;
    wire signal_9058 ;
    wire signal_9059 ;
    wire signal_9060 ;
    wire signal_9061 ;
    wire signal_9062 ;
    wire signal_9063 ;
    wire signal_9064 ;
    wire signal_9065 ;
    wire signal_9066 ;
    wire signal_9067 ;
    wire signal_9068 ;
    wire signal_9069 ;
    wire signal_9070 ;
    wire signal_9071 ;
    wire signal_9072 ;
    wire signal_9073 ;
    wire signal_9074 ;
    wire signal_9075 ;
    wire signal_9076 ;
    wire signal_9077 ;
    wire signal_9078 ;
    wire signal_9079 ;
    wire signal_9080 ;
    wire signal_9081 ;
    wire signal_9082 ;
    wire signal_9083 ;
    wire signal_9084 ;
    wire signal_9085 ;
    wire signal_9086 ;
    wire signal_9087 ;
    wire signal_9088 ;
    wire signal_9089 ;
    wire signal_9090 ;
    wire signal_9091 ;
    wire signal_9092 ;
    wire signal_9093 ;
    wire signal_9094 ;
    wire signal_9095 ;
    wire signal_9096 ;
    wire signal_9097 ;
    wire signal_9098 ;
    wire signal_9099 ;
    wire signal_9100 ;
    wire signal_9101 ;
    wire signal_9102 ;
    wire signal_9103 ;
    wire signal_9104 ;
    wire signal_9105 ;
    wire signal_9106 ;
    wire signal_9107 ;
    wire signal_9108 ;
    wire signal_9109 ;
    wire signal_9110 ;
    wire signal_9111 ;
    wire signal_9112 ;
    wire signal_9113 ;
    wire signal_9114 ;
    wire signal_9115 ;
    wire signal_9116 ;
    wire signal_9117 ;
    wire signal_9118 ;
    wire signal_9119 ;
    wire signal_9120 ;
    wire signal_9121 ;
    wire signal_9122 ;
    wire signal_9123 ;
    wire signal_9124 ;
    wire signal_9125 ;
    wire signal_9126 ;
    wire signal_9127 ;
    wire signal_9128 ;
    wire signal_9129 ;
    wire signal_9130 ;
    wire signal_9131 ;
    wire signal_9132 ;
    wire signal_9133 ;
    wire signal_9134 ;
    wire signal_9135 ;
    wire signal_9136 ;
    wire signal_9137 ;
    wire signal_9138 ;
    wire signal_9139 ;
    wire signal_9140 ;
    wire signal_9141 ;
    wire signal_9142 ;
    wire signal_9143 ;
    wire signal_9144 ;
    wire signal_9145 ;
    wire signal_9146 ;
    wire signal_9147 ;
    wire signal_9148 ;
    wire signal_9149 ;
    wire signal_9150 ;
    wire signal_9151 ;
    wire signal_9152 ;
    wire signal_9153 ;
    wire signal_9154 ;
    wire signal_9155 ;
    wire signal_9156 ;
    wire signal_9157 ;
    wire signal_9158 ;
    wire signal_9159 ;
    wire signal_9160 ;
    wire signal_9161 ;
    wire signal_9162 ;
    wire signal_9163 ;
    wire signal_9164 ;
    wire signal_9165 ;
    wire signal_9166 ;
    wire signal_9167 ;
    wire signal_9168 ;
    wire signal_9169 ;
    wire signal_9170 ;
    wire signal_9171 ;
    wire signal_9172 ;
    wire signal_9173 ;
    wire signal_9174 ;
    wire signal_9175 ;
    wire signal_9176 ;
    wire signal_9177 ;
    wire signal_9178 ;
    wire signal_9179 ;
    wire signal_9180 ;
    wire signal_9181 ;
    wire signal_9182 ;
    wire signal_9183 ;
    wire signal_9184 ;
    wire signal_9185 ;
    wire signal_9186 ;
    wire signal_9187 ;
    wire signal_9188 ;
    wire signal_9189 ;
    wire signal_9190 ;
    wire signal_9191 ;
    wire signal_9192 ;
    wire signal_9193 ;
    wire signal_9194 ;
    wire signal_9195 ;
    wire signal_9196 ;
    wire signal_9197 ;
    wire signal_9198 ;
    wire signal_9199 ;
    wire signal_9200 ;
    wire signal_9201 ;
    wire signal_9202 ;
    wire signal_9203 ;
    wire signal_9204 ;
    wire signal_9205 ;
    wire signal_9206 ;
    wire signal_9207 ;
    wire signal_9208 ;
    wire signal_9209 ;
    wire signal_9210 ;
    wire signal_9211 ;
    wire signal_9212 ;
    wire signal_9213 ;
    wire signal_9214 ;
    wire signal_9215 ;
    wire signal_9216 ;
    wire signal_9217 ;
    wire signal_9218 ;
    wire signal_9219 ;
    wire signal_9220 ;
    wire signal_9221 ;
    wire signal_9222 ;
    wire signal_9223 ;
    wire signal_9224 ;
    wire signal_9225 ;
    wire signal_9226 ;
    wire signal_9227 ;
    wire signal_9228 ;
    wire signal_9229 ;
    wire signal_9230 ;
    wire signal_9231 ;
    wire signal_9232 ;
    wire signal_9233 ;
    wire signal_9234 ;
    wire signal_9235 ;
    wire signal_9236 ;
    wire signal_9237 ;
    wire signal_9238 ;
    wire signal_9239 ;
    wire signal_9240 ;
    wire signal_9241 ;
    wire signal_9242 ;
    wire signal_9243 ;
    wire signal_9244 ;
    wire signal_9245 ;
    wire signal_9246 ;
    wire signal_9247 ;
    wire signal_9248 ;
    wire signal_9249 ;
    wire signal_9250 ;
    wire signal_9251 ;
    wire signal_9252 ;
    wire signal_9253 ;
    wire signal_9254 ;
    wire signal_9255 ;
    wire signal_9256 ;
    wire signal_9257 ;
    wire signal_9258 ;
    wire signal_9259 ;
    wire signal_9260 ;
    wire signal_9261 ;
    wire signal_9262 ;
    wire signal_9263 ;
    wire signal_9264 ;
    wire signal_9265 ;
    wire signal_9266 ;
    wire signal_9267 ;
    wire signal_9268 ;
    wire signal_9269 ;
    wire signal_9270 ;
    wire signal_9271 ;
    wire signal_9272 ;
    wire signal_9273 ;
    wire signal_9274 ;
    wire signal_9275 ;
    wire signal_9276 ;
    wire signal_9277 ;
    wire signal_9278 ;
    wire signal_9279 ;
    wire signal_9280 ;
    wire signal_9281 ;
    wire signal_9282 ;
    wire signal_9283 ;
    wire signal_9284 ;
    wire signal_9285 ;
    wire signal_9286 ;
    wire signal_9287 ;
    wire signal_9288 ;
    wire signal_9289 ;
    wire signal_9290 ;
    wire signal_9291 ;
    wire signal_9292 ;
    wire signal_9293 ;
    wire signal_9294 ;
    wire signal_9295 ;
    wire signal_9296 ;
    wire signal_9297 ;
    wire signal_9298 ;
    wire signal_9299 ;
    wire signal_9300 ;
    wire signal_9301 ;
    wire signal_9302 ;
    wire signal_9303 ;
    wire signal_9304 ;
    wire signal_9305 ;
    wire signal_9306 ;
    wire signal_9307 ;
    wire signal_9308 ;
    wire signal_9309 ;
    wire signal_9310 ;
    wire signal_9311 ;
    wire signal_9312 ;
    wire signal_9313 ;
    wire signal_9314 ;
    wire signal_9315 ;
    wire signal_9316 ;
    wire signal_9317 ;
    wire signal_9318 ;
    wire signal_9319 ;
    wire signal_9320 ;
    wire signal_9321 ;
    wire signal_9322 ;
    wire signal_9323 ;
    wire signal_9324 ;
    wire signal_9325 ;
    wire signal_9326 ;
    wire signal_9327 ;
    wire signal_9328 ;
    wire signal_9329 ;
    wire signal_9330 ;
    wire signal_9331 ;
    wire signal_9332 ;
    wire signal_9333 ;
    wire signal_9334 ;
    wire signal_9335 ;
    wire signal_9336 ;
    wire signal_9337 ;
    wire signal_9338 ;
    wire signal_9339 ;
    wire signal_9340 ;
    wire signal_9341 ;
    wire signal_9342 ;
    wire signal_9343 ;
    wire signal_9344 ;
    wire signal_9345 ;
    wire signal_9346 ;
    wire signal_9347 ;
    wire signal_9348 ;
    wire signal_9349 ;
    wire signal_9350 ;
    wire signal_9351 ;
    wire signal_9352 ;
    wire signal_9353 ;
    wire signal_9354 ;
    wire signal_9355 ;
    wire signal_9356 ;
    wire signal_9357 ;
    wire signal_9358 ;
    wire signal_9359 ;
    wire signal_9360 ;
    wire signal_9361 ;
    wire signal_9362 ;
    wire signal_9363 ;
    wire signal_9364 ;
    wire signal_9365 ;
    wire signal_9366 ;
    wire signal_9367 ;
    wire signal_9368 ;
    wire signal_9369 ;
    wire signal_9370 ;
    wire signal_9371 ;
    wire signal_9372 ;
    wire signal_9373 ;
    wire signal_9374 ;
    wire signal_9375 ;
    wire signal_9376 ;
    wire signal_9377 ;
    wire signal_9378 ;
    wire signal_9379 ;
    wire signal_9380 ;
    wire signal_9381 ;
    wire signal_9382 ;
    wire signal_9383 ;
    wire signal_9384 ;
    wire signal_9385 ;
    wire signal_9386 ;
    wire signal_9387 ;
    wire signal_9388 ;
    wire signal_9389 ;
    wire signal_9390 ;
    wire signal_9391 ;
    wire signal_9392 ;
    wire signal_9393 ;
    wire signal_9394 ;
    wire signal_9395 ;
    wire signal_9396 ;
    wire signal_9397 ;
    wire signal_9398 ;
    wire signal_9399 ;
    wire signal_9400 ;
    wire signal_9401 ;
    wire signal_9402 ;
    wire signal_9403 ;
    wire signal_9404 ;
    wire signal_9405 ;
    wire signal_9406 ;
    wire signal_9407 ;
    wire signal_9408 ;
    wire signal_9409 ;
    wire signal_9410 ;
    wire signal_9411 ;
    wire signal_9412 ;
    wire signal_9413 ;
    wire signal_9414 ;
    wire signal_9415 ;
    wire signal_9416 ;
    wire signal_9417 ;
    wire signal_9418 ;
    wire signal_9419 ;
    wire signal_9420 ;
    wire signal_9421 ;
    wire signal_9422 ;
    wire signal_9423 ;
    wire signal_9424 ;
    wire signal_9425 ;
    wire signal_9426 ;
    wire signal_9427 ;
    wire signal_9428 ;
    wire signal_9429 ;
    wire signal_9430 ;
    wire signal_9431 ;
    wire signal_9432 ;
    wire signal_9433 ;
    wire signal_9434 ;
    wire signal_9435 ;
    wire signal_9436 ;
    wire signal_9437 ;
    wire signal_9438 ;
    wire signal_9439 ;
    wire signal_9440 ;
    wire signal_9441 ;
    wire signal_9442 ;
    wire signal_9443 ;
    wire signal_9444 ;
    wire signal_9445 ;
    wire signal_9446 ;
    wire signal_9447 ;
    wire signal_9448 ;
    wire signal_9449 ;
    wire signal_9450 ;
    wire signal_9451 ;
    wire signal_9452 ;
    wire signal_9453 ;
    wire signal_9454 ;
    wire signal_9455 ;
    wire signal_9456 ;
    wire signal_9457 ;
    wire signal_9458 ;
    wire signal_9459 ;
    wire signal_9460 ;
    wire signal_9461 ;
    wire signal_9462 ;
    wire signal_9463 ;
    wire signal_9464 ;
    wire signal_9465 ;
    wire signal_9466 ;
    wire signal_9467 ;
    wire signal_9468 ;
    wire signal_9469 ;
    wire signal_9470 ;
    wire signal_9471 ;
    wire signal_9472 ;
    wire signal_9473 ;
    wire signal_9474 ;
    wire signal_9475 ;
    wire signal_9476 ;
    wire signal_9477 ;
    wire signal_9478 ;
    wire signal_9479 ;
    wire signal_9480 ;
    wire signal_9481 ;
    wire signal_9482 ;
    wire signal_9483 ;
    wire signal_9484 ;
    wire signal_9485 ;
    wire signal_9486 ;
    wire signal_9487 ;
    wire signal_9488 ;
    wire signal_9489 ;
    wire signal_9490 ;
    wire signal_9491 ;
    wire signal_9492 ;
    wire signal_9493 ;
    wire signal_9494 ;
    wire signal_9495 ;
    wire signal_9496 ;
    wire signal_9497 ;
    wire signal_9498 ;
    wire signal_9499 ;
    wire signal_9500 ;
    wire signal_9501 ;
    wire signal_9502 ;
    wire signal_9503 ;
    wire signal_9504 ;
    wire signal_9505 ;
    wire signal_9506 ;
    wire signal_9507 ;
    wire signal_9508 ;
    wire signal_9509 ;
    wire signal_9510 ;
    wire signal_9511 ;
    wire signal_9512 ;
    wire signal_9513 ;
    wire signal_9514 ;
    wire signal_9515 ;
    wire signal_9516 ;
    wire signal_9517 ;
    wire signal_9518 ;
    wire signal_9519 ;
    wire signal_9520 ;
    wire signal_9521 ;
    wire signal_9522 ;
    wire signal_9523 ;
    wire signal_9524 ;
    wire signal_9525 ;
    wire signal_9526 ;
    wire signal_9527 ;
    wire signal_9528 ;
    wire signal_9529 ;
    wire signal_9530 ;
    wire signal_9531 ;
    wire signal_9532 ;
    wire signal_9533 ;
    wire signal_9534 ;
    wire signal_9535 ;
    wire signal_9536 ;
    wire signal_9537 ;
    wire signal_9538 ;
    wire signal_9539 ;
    wire signal_9540 ;
    wire signal_9541 ;
    wire signal_9542 ;
    wire signal_9543 ;
    wire signal_9544 ;
    wire signal_9545 ;
    wire signal_9546 ;
    wire signal_9547 ;
    wire signal_9548 ;
    wire signal_9549 ;
    wire signal_9550 ;
    wire signal_9551 ;
    wire signal_9552 ;
    wire signal_9553 ;
    wire signal_9554 ;
    wire signal_9555 ;
    wire signal_9556 ;
    wire signal_9557 ;
    wire signal_9558 ;
    wire signal_9559 ;
    wire signal_9560 ;
    wire signal_9561 ;
    wire signal_9562 ;
    wire signal_9563 ;
    wire signal_9564 ;
    wire signal_9565 ;
    wire signal_9566 ;
    wire signal_9567 ;
    wire signal_9568 ;
    wire signal_9569 ;
    wire signal_9570 ;
    wire signal_9571 ;
    wire signal_9572 ;
    wire signal_9573 ;
    wire signal_9574 ;
    wire signal_9575 ;
    wire signal_9576 ;
    wire signal_9577 ;
    wire signal_9578 ;
    wire signal_9579 ;
    wire signal_9580 ;
    wire signal_9581 ;
    wire signal_9582 ;
    wire signal_9583 ;
    wire signal_9584 ;
    wire signal_9585 ;
    wire signal_9586 ;
    wire signal_9587 ;
    wire signal_9588 ;
    wire signal_9589 ;
    wire signal_9590 ;
    wire signal_9591 ;
    wire signal_9592 ;
    wire signal_9593 ;
    wire signal_9594 ;
    wire signal_9595 ;
    wire signal_9596 ;
    wire signal_9597 ;
    wire signal_9598 ;
    wire signal_9599 ;
    wire signal_9600 ;
    wire signal_9601 ;
    wire signal_9602 ;
    wire signal_9603 ;
    wire signal_9604 ;
    wire signal_9605 ;
    wire signal_9606 ;
    wire signal_9607 ;
    wire signal_9608 ;
    wire signal_9609 ;
    wire signal_9610 ;
    wire signal_9611 ;
    wire signal_9612 ;
    wire signal_9613 ;
    wire signal_9614 ;
    wire signal_9615 ;
    wire signal_9616 ;
    wire signal_9617 ;
    wire signal_9618 ;
    wire signal_9619 ;
    wire signal_9620 ;
    wire signal_9621 ;
    wire signal_9622 ;
    wire signal_9623 ;
    wire signal_9624 ;
    wire signal_9625 ;
    wire signal_9626 ;
    wire signal_9627 ;
    wire signal_9628 ;
    wire signal_9629 ;
    wire signal_9630 ;
    wire signal_9631 ;
    wire signal_9632 ;
    wire signal_9633 ;
    wire signal_9634 ;
    wire signal_9635 ;
    wire signal_9636 ;
    wire signal_9637 ;
    wire signal_9638 ;
    wire signal_9639 ;
    wire signal_9640 ;
    wire signal_9641 ;
    wire signal_9642 ;
    wire signal_9643 ;
    wire signal_9644 ;
    wire signal_9645 ;
    wire signal_9646 ;
    wire signal_9647 ;
    wire signal_9648 ;
    wire signal_9649 ;
    wire signal_9650 ;
    wire signal_9651 ;
    wire signal_9652 ;
    wire signal_9653 ;
    wire signal_9654 ;
    wire signal_9655 ;
    wire signal_9656 ;
    wire signal_9657 ;
    wire signal_9658 ;
    wire signal_9659 ;
    wire signal_9660 ;
    wire signal_9661 ;
    wire signal_9662 ;
    wire signal_9663 ;
    wire signal_9664 ;
    wire signal_9665 ;
    wire signal_9666 ;
    wire signal_9667 ;
    wire signal_9668 ;
    wire signal_9669 ;
    wire signal_9670 ;
    wire signal_9671 ;
    wire signal_9672 ;
    wire signal_9673 ;
    wire signal_9674 ;
    wire signal_9675 ;
    wire signal_9676 ;
    wire signal_9677 ;
    wire signal_9678 ;
    wire signal_9679 ;
    wire signal_9680 ;
    wire signal_9681 ;
    wire signal_9682 ;
    wire signal_9683 ;
    wire signal_9684 ;
    wire signal_9685 ;
    wire signal_9686 ;
    wire signal_9687 ;
    wire signal_9688 ;
    wire signal_9689 ;
    wire signal_9690 ;
    wire signal_9691 ;
    wire signal_9692 ;
    wire signal_9693 ;
    wire signal_9694 ;
    wire signal_9695 ;
    wire signal_9696 ;
    wire signal_9697 ;
    wire signal_9698 ;
    wire signal_9699 ;
    wire signal_9700 ;
    wire signal_9701 ;
    wire signal_9702 ;
    wire signal_9703 ;
    wire signal_9704 ;
    wire signal_9705 ;
    wire signal_9706 ;
    wire signal_9707 ;
    wire signal_9708 ;
    wire signal_9709 ;
    wire signal_9710 ;
    wire signal_9711 ;
    wire signal_9712 ;
    wire signal_9713 ;
    wire signal_9714 ;
    wire signal_9715 ;
    wire signal_9716 ;
    wire signal_9717 ;
    wire signal_9718 ;
    wire signal_9719 ;
    wire signal_9720 ;
    wire signal_9721 ;
    wire signal_9722 ;
    wire signal_9723 ;
    wire signal_9724 ;
    wire signal_9725 ;
    wire signal_9726 ;
    wire signal_9727 ;
    wire signal_9728 ;
    wire signal_9729 ;
    wire signal_9730 ;
    wire signal_9731 ;
    wire signal_9732 ;
    wire signal_9733 ;
    wire signal_9734 ;
    wire signal_9735 ;
    wire signal_9736 ;
    wire signal_9737 ;
    wire signal_9738 ;
    wire signal_9739 ;
    wire signal_9740 ;
    wire signal_9741 ;
    wire signal_9742 ;
    wire signal_9743 ;
    wire signal_9744 ;
    wire signal_9745 ;
    wire signal_9746 ;
    wire signal_9747 ;
    wire signal_9748 ;
    wire signal_9749 ;
    wire signal_9750 ;
    wire signal_9751 ;
    wire signal_9752 ;
    wire signal_9753 ;
    wire signal_9754 ;
    wire signal_9755 ;
    wire signal_9756 ;
    wire signal_9757 ;
    wire signal_9758 ;
    wire signal_9759 ;
    wire signal_9760 ;
    wire signal_9761 ;
    wire signal_9762 ;
    wire signal_9763 ;
    wire signal_9764 ;
    wire signal_9765 ;
    wire signal_9766 ;
    wire signal_9767 ;
    wire signal_9768 ;
    wire signal_9769 ;
    wire signal_9770 ;
    wire signal_9771 ;
    wire signal_9772 ;
    wire signal_9773 ;
    wire signal_9774 ;
    wire signal_9775 ;
    wire signal_9776 ;
    wire signal_9777 ;
    wire signal_9778 ;
    wire signal_9779 ;
    wire signal_9780 ;
    wire signal_9781 ;
    wire signal_9782 ;
    wire signal_9783 ;
    wire signal_9784 ;
    wire signal_9785 ;
    wire signal_9786 ;
    wire signal_9787 ;
    wire signal_9788 ;
    wire signal_9789 ;
    wire signal_9790 ;
    wire signal_9791 ;
    wire signal_9792 ;
    wire signal_9793 ;
    wire signal_9794 ;
    wire signal_9795 ;
    wire signal_9796 ;
    wire signal_9797 ;
    wire signal_9798 ;
    wire signal_9799 ;
    wire signal_9800 ;
    wire signal_9801 ;
    wire signal_9802 ;
    wire signal_9803 ;
    wire signal_9804 ;
    wire signal_9805 ;
    wire signal_9806 ;
    wire signal_9807 ;
    wire signal_9808 ;
    wire signal_9809 ;
    wire signal_9810 ;
    wire signal_9811 ;
    wire signal_9812 ;
    wire signal_9813 ;
    wire signal_9814 ;
    wire signal_9815 ;
    wire signal_9816 ;
    wire signal_9817 ;
    wire signal_9818 ;
    wire signal_9819 ;
    wire signal_9820 ;
    wire signal_9821 ;
    wire signal_9822 ;
    wire signal_9823 ;
    wire signal_9824 ;
    wire signal_9825 ;
    wire signal_9826 ;
    wire signal_9827 ;
    wire signal_9828 ;
    wire signal_9829 ;
    wire signal_9830 ;
    wire signal_9831 ;
    wire signal_9832 ;
    wire signal_9833 ;
    wire signal_9834 ;
    wire signal_9835 ;
    wire signal_9836 ;
    wire signal_9837 ;
    wire signal_9838 ;
    wire signal_9839 ;
    wire signal_9840 ;
    wire signal_9841 ;
    wire signal_9842 ;
    wire signal_9843 ;
    wire signal_9844 ;
    wire signal_9845 ;
    wire signal_9846 ;
    wire signal_9847 ;
    wire signal_9848 ;
    wire signal_9849 ;
    wire signal_9850 ;
    wire signal_9851 ;
    wire signal_9852 ;
    wire signal_9853 ;
    wire signal_9854 ;
    wire signal_9855 ;
    wire signal_9856 ;
    wire signal_9857 ;
    wire signal_9858 ;
    wire signal_9859 ;
    wire signal_9860 ;
    wire signal_9861 ;
    wire signal_9862 ;
    wire signal_9863 ;
    wire signal_9864 ;
    wire signal_9865 ;
    wire signal_9866 ;
    wire signal_9867 ;
    wire signal_9868 ;
    wire signal_9869 ;
    wire signal_9870 ;
    wire signal_9871 ;
    wire signal_9872 ;
    wire signal_9873 ;
    wire signal_9874 ;
    wire signal_9875 ;
    wire signal_9876 ;
    wire signal_9877 ;
    wire signal_9878 ;
    wire signal_9879 ;
    wire signal_9880 ;
    wire signal_9881 ;
    wire signal_9882 ;
    wire signal_9883 ;
    wire signal_9884 ;
    wire signal_9885 ;
    wire signal_9886 ;
    wire signal_9887 ;
    wire signal_9888 ;
    wire signal_9889 ;
    wire signal_9890 ;
    wire signal_9891 ;
    wire signal_9892 ;
    wire signal_9893 ;
    wire signal_9894 ;
    wire signal_9895 ;
    wire signal_9896 ;
    wire signal_9897 ;
    wire signal_9898 ;
    wire signal_9899 ;
    wire signal_9900 ;
    wire signal_9901 ;
    wire signal_9902 ;
    wire signal_9903 ;
    wire signal_9904 ;
    wire signal_9905 ;
    wire signal_9906 ;
    wire signal_9907 ;
    wire signal_9908 ;
    wire signal_9909 ;
    wire signal_9910 ;
    wire signal_9911 ;
    wire signal_9912 ;
    wire signal_9913 ;
    wire signal_9914 ;
    wire signal_9915 ;
    wire signal_9916 ;
    wire signal_9917 ;
    wire signal_9918 ;
    wire signal_9919 ;
    wire signal_9920 ;
    wire signal_9921 ;
    wire signal_9922 ;
    wire signal_9923 ;
    wire signal_9924 ;
    wire signal_9925 ;
    wire signal_9926 ;
    wire signal_9927 ;
    wire signal_9928 ;
    wire signal_9929 ;
    wire signal_9930 ;
    wire signal_9931 ;
    wire signal_9932 ;
    wire signal_9933 ;
    wire signal_9934 ;
    wire signal_9935 ;
    wire signal_9936 ;
    wire signal_9937 ;
    wire signal_9938 ;
    wire signal_9939 ;
    wire signal_9940 ;
    wire signal_9941 ;
    wire signal_9942 ;
    wire signal_9943 ;
    wire signal_9944 ;
    wire signal_9945 ;
    wire signal_9946 ;
    wire signal_9947 ;
    wire signal_9948 ;
    wire signal_9949 ;
    wire signal_9950 ;
    wire signal_9951 ;
    wire signal_9952 ;
    wire signal_9953 ;
    wire signal_9954 ;
    wire signal_9955 ;
    wire signal_9956 ;
    wire signal_9957 ;
    wire signal_9958 ;
    wire signal_9959 ;
    wire signal_9960 ;
    wire signal_9961 ;
    wire signal_9962 ;
    wire signal_9963 ;
    wire signal_9964 ;
    wire signal_9965 ;
    wire signal_9966 ;
    wire signal_9967 ;
    wire signal_9968 ;
    wire signal_9969 ;
    wire signal_9970 ;
    wire signal_9971 ;
    wire signal_9972 ;
    wire signal_9973 ;
    wire signal_9974 ;
    wire signal_9975 ;
    wire signal_9976 ;
    wire signal_9977 ;
    wire signal_9978 ;
    wire signal_9979 ;
    wire signal_9980 ;
    wire signal_9981 ;
    wire signal_9982 ;
    wire signal_9983 ;
    wire signal_9984 ;
    wire signal_9985 ;
    wire signal_9986 ;
    wire signal_9987 ;
    wire signal_9988 ;
    wire signal_9989 ;
    wire signal_9990 ;
    wire signal_9991 ;
    wire signal_9992 ;
    wire signal_9993 ;
    wire signal_9994 ;
    wire signal_9995 ;
    wire signal_9996 ;
    wire signal_9997 ;
    wire signal_9998 ;
    wire signal_9999 ;
    wire signal_10000 ;
    wire signal_10001 ;
    wire signal_10002 ;
    wire signal_10003 ;
    wire signal_10004 ;
    wire signal_10005 ;
    wire signal_10006 ;
    wire signal_10007 ;
    wire signal_10008 ;
    wire signal_10009 ;
    wire signal_10010 ;
    wire signal_10011 ;
    wire signal_10012 ;
    wire signal_10013 ;
    wire signal_10014 ;
    wire signal_10015 ;
    wire signal_10016 ;
    wire signal_10017 ;
    wire signal_10018 ;
    wire signal_10019 ;
    wire signal_10020 ;
    wire signal_10021 ;
    wire signal_10022 ;
    wire signal_10023 ;
    wire signal_10024 ;
    wire signal_10025 ;
    wire signal_10026 ;
    wire signal_10027 ;
    wire signal_10028 ;
    wire signal_10029 ;
    wire signal_10030 ;
    wire signal_10031 ;
    wire signal_10032 ;
    wire signal_10033 ;
    wire signal_10034 ;
    wire signal_10035 ;
    wire signal_10036 ;
    wire signal_10037 ;
    wire signal_10038 ;
    wire signal_10039 ;
    wire signal_10040 ;
    wire signal_10041 ;
    wire signal_10042 ;
    wire signal_10043 ;
    wire signal_10044 ;
    wire signal_10045 ;
    wire signal_10046 ;
    wire signal_10047 ;
    wire signal_10048 ;
    wire signal_10049 ;
    wire signal_10050 ;
    wire signal_10051 ;
    wire signal_10052 ;
    wire signal_10053 ;
    wire signal_10054 ;
    wire signal_10055 ;
    wire signal_10056 ;
    wire signal_10057 ;
    wire signal_10058 ;
    wire signal_10059 ;
    wire signal_10060 ;
    wire signal_10061 ;
    wire signal_10062 ;
    wire signal_10063 ;
    wire signal_10064 ;
    wire signal_10065 ;
    wire signal_10066 ;
    wire signal_10067 ;
    wire signal_10068 ;
    wire signal_10069 ;
    wire signal_10070 ;
    wire signal_10071 ;
    wire signal_10072 ;
    wire signal_10073 ;
    wire signal_10074 ;
    wire signal_10075 ;
    wire signal_10076 ;
    wire signal_10077 ;
    wire signal_10078 ;
    wire signal_10079 ;
    wire signal_10080 ;
    wire signal_10081 ;
    wire signal_10082 ;
    wire signal_10083 ;
    wire signal_10084 ;
    wire signal_10085 ;
    wire signal_10086 ;
    wire signal_10087 ;
    wire signal_10088 ;
    wire signal_10089 ;
    wire signal_10090 ;
    wire signal_10091 ;
    wire signal_10092 ;
    wire signal_10093 ;
    wire signal_10094 ;
    wire signal_10095 ;
    wire signal_10096 ;
    wire signal_10097 ;
    wire signal_10098 ;
    wire signal_10099 ;
    wire signal_10100 ;
    wire signal_10101 ;
    wire signal_10102 ;
    wire signal_10103 ;
    wire signal_10104 ;
    wire signal_10105 ;
    wire signal_10106 ;
    wire signal_10107 ;
    wire signal_10108 ;
    wire signal_10109 ;
    wire signal_10110 ;
    wire signal_10111 ;
    wire signal_10112 ;
    wire signal_10113 ;
    wire signal_10114 ;
    wire signal_10115 ;
    wire signal_10116 ;
    wire signal_10117 ;
    wire signal_10118 ;
    wire signal_10119 ;
    wire signal_10120 ;
    wire signal_10121 ;
    wire signal_10122 ;
    wire signal_10123 ;
    wire signal_10124 ;
    wire signal_10125 ;
    wire signal_10126 ;
    wire signal_10127 ;
    wire signal_10128 ;
    wire signal_10129 ;
    wire signal_10130 ;
    wire signal_10131 ;
    wire signal_10132 ;
    wire signal_10133 ;
    wire signal_10134 ;
    wire signal_10135 ;
    wire signal_10136 ;
    wire signal_10137 ;
    wire signal_10138 ;
    wire signal_10139 ;
    wire signal_10140 ;
    wire signal_10141 ;
    wire signal_10142 ;
    wire signal_10143 ;
    wire signal_10144 ;
    wire signal_10145 ;
    wire signal_10146 ;
    wire signal_10147 ;
    wire signal_10148 ;
    wire signal_10149 ;
    wire signal_10150 ;
    wire signal_10151 ;
    wire signal_10152 ;
    wire signal_10153 ;
    wire signal_10154 ;
    wire signal_10155 ;
    wire signal_10156 ;
    wire signal_10157 ;
    wire signal_10158 ;
    wire signal_10159 ;
    wire signal_10160 ;
    wire signal_10161 ;
    wire signal_10162 ;
    wire signal_10163 ;
    wire signal_10164 ;
    wire signal_10165 ;
    wire signal_10166 ;
    wire signal_10167 ;
    wire signal_10168 ;
    wire signal_10169 ;
    wire signal_10170 ;
    wire signal_10171 ;
    wire signal_10172 ;
    wire signal_10173 ;
    wire signal_10174 ;
    wire signal_10175 ;
    wire signal_10176 ;
    wire signal_10177 ;
    wire signal_10178 ;
    wire signal_10179 ;
    wire signal_10180 ;
    wire signal_10181 ;
    wire signal_10182 ;
    wire signal_10183 ;
    wire signal_10184 ;
    wire signal_10185 ;
    wire signal_10186 ;
    wire signal_10187 ;
    wire signal_10188 ;
    wire signal_10189 ;
    wire signal_10190 ;
    wire signal_10191 ;
    wire signal_10192 ;
    wire signal_10193 ;
    wire signal_10194 ;
    wire signal_10195 ;
    wire signal_10196 ;
    wire signal_10197 ;
    wire signal_10198 ;
    wire signal_10199 ;
    wire signal_10200 ;
    wire signal_10201 ;
    wire signal_10202 ;
    wire signal_10203 ;
    wire signal_10204 ;
    wire signal_10205 ;
    wire signal_10206 ;
    wire signal_10207 ;
    wire signal_10208 ;
    wire signal_10209 ;
    wire signal_10210 ;
    wire signal_10211 ;
    wire signal_10212 ;
    wire signal_10213 ;
    wire signal_10214 ;
    wire signal_10215 ;
    wire signal_10216 ;
    wire signal_10217 ;
    wire signal_10218 ;
    wire signal_10219 ;
    wire signal_10220 ;
    wire signal_10221 ;
    wire signal_10222 ;
    wire signal_10223 ;
    wire signal_10224 ;
    wire signal_10225 ;
    wire signal_10226 ;
    wire signal_10227 ;
    wire signal_10228 ;
    wire signal_10229 ;
    wire signal_10230 ;
    wire signal_10231 ;
    wire signal_10232 ;
    wire signal_10233 ;
    wire signal_10234 ;
    wire signal_10235 ;
    wire signal_10236 ;
    wire signal_10237 ;
    wire signal_10238 ;
    wire signal_10239 ;
    wire signal_10240 ;
    wire signal_10241 ;
    wire signal_10242 ;
    wire signal_10243 ;
    wire signal_10244 ;
    wire signal_10245 ;
    wire signal_10246 ;
    wire signal_10247 ;
    wire signal_10248 ;
    wire signal_10249 ;
    wire signal_10250 ;
    wire signal_10251 ;
    wire signal_10252 ;
    wire signal_10253 ;
    wire signal_10254 ;
    wire signal_10255 ;
    wire signal_10256 ;
    wire signal_10257 ;
    wire signal_10258 ;
    wire signal_10259 ;
    wire signal_10260 ;
    wire signal_10261 ;
    wire signal_10262 ;
    wire signal_10263 ;
    wire signal_10264 ;
    wire signal_10265 ;
    wire signal_10266 ;
    wire signal_10267 ;
    wire signal_10268 ;
    wire signal_10269 ;
    wire signal_10270 ;
    wire signal_10271 ;
    wire signal_10272 ;
    wire signal_10273 ;
    wire signal_10274 ;
    wire signal_10275 ;
    wire signal_10276 ;
    wire signal_10277 ;
    wire signal_10278 ;
    wire signal_10279 ;
    wire signal_10280 ;
    wire signal_10281 ;
    wire signal_10282 ;
    wire signal_10283 ;
    wire signal_10284 ;
    wire signal_10285 ;
    wire signal_10286 ;
    wire signal_10287 ;
    wire signal_10288 ;
    wire signal_10289 ;
    wire signal_10290 ;
    wire signal_10291 ;
    wire signal_10292 ;
    wire signal_10293 ;
    wire signal_10294 ;
    wire signal_10295 ;
    wire signal_10296 ;
    wire signal_10297 ;
    wire signal_10298 ;
    wire signal_10299 ;
    wire signal_10300 ;
    wire signal_10301 ;
    wire signal_10302 ;
    wire signal_10303 ;
    wire signal_10304 ;
    wire signal_10305 ;
    wire signal_10306 ;
    wire signal_10307 ;
    wire signal_10308 ;
    wire signal_10309 ;
    wire signal_10310 ;
    wire signal_10311 ;
    wire signal_10312 ;
    wire signal_10313 ;
    wire signal_10314 ;
    wire signal_10315 ;
    wire signal_10316 ;
    wire signal_10317 ;
    wire signal_10318 ;
    wire signal_10319 ;
    wire signal_10320 ;
    wire signal_10321 ;
    wire signal_10322 ;
    wire signal_10323 ;
    wire signal_10324 ;
    wire signal_10325 ;
    wire signal_10326 ;
    wire signal_10327 ;
    wire signal_10328 ;
    wire signal_10329 ;
    wire signal_10330 ;
    wire signal_10331 ;
    wire signal_10332 ;
    wire signal_10333 ;
    wire signal_10334 ;
    wire signal_10335 ;
    wire signal_10336 ;
    wire signal_10337 ;
    wire signal_10338 ;
    wire signal_10339 ;
    wire signal_10340 ;
    wire signal_10341 ;
    wire signal_10342 ;
    wire signal_10343 ;
    wire signal_10344 ;
    wire signal_10345 ;
    wire signal_10346 ;
    wire signal_10347 ;
    wire signal_10348 ;
    wire signal_10349 ;
    wire signal_10350 ;
    wire signal_10351 ;
    wire signal_10352 ;
    wire signal_10353 ;
    wire signal_10354 ;
    wire signal_10355 ;
    wire signal_10356 ;
    wire signal_10357 ;
    wire signal_10358 ;
    wire signal_10359 ;
    wire signal_10360 ;
    wire signal_10361 ;
    wire signal_10362 ;
    wire signal_10363 ;
    wire signal_10364 ;
    wire signal_10365 ;
    wire signal_10366 ;
    wire signal_10367 ;
    wire signal_10368 ;
    wire signal_10369 ;
    wire signal_10370 ;
    wire signal_10371 ;
    wire signal_10372 ;
    wire signal_10373 ;
    wire signal_10374 ;
    wire signal_10375 ;
    wire signal_10376 ;
    wire signal_10377 ;
    wire signal_10378 ;
    wire signal_10379 ;
    wire signal_10380 ;
    wire signal_10381 ;
    wire signal_10382 ;
    wire signal_10383 ;
    wire signal_10384 ;
    wire signal_10385 ;
    wire signal_10386 ;
    wire signal_10387 ;
    wire signal_10388 ;
    wire signal_10389 ;
    wire signal_10390 ;
    wire signal_10391 ;
    wire signal_10392 ;
    wire signal_10393 ;
    wire signal_10394 ;
    wire signal_10395 ;
    wire signal_10396 ;
    wire signal_10397 ;
    wire signal_10398 ;
    wire signal_10399 ;
    wire signal_10400 ;
    wire signal_10401 ;
    wire signal_10402 ;
    wire signal_10403 ;
    wire signal_10404 ;
    wire signal_10405 ;
    wire signal_10406 ;
    wire signal_10407 ;
    wire signal_10408 ;
    wire signal_10409 ;
    wire signal_10410 ;
    wire signal_10411 ;
    wire signal_10412 ;
    wire signal_10413 ;
    wire signal_10414 ;
    wire signal_10415 ;
    wire signal_10416 ;
    wire signal_10417 ;
    wire signal_10418 ;
    wire signal_10419 ;
    wire signal_10420 ;
    wire signal_10421 ;
    wire signal_10422 ;
    wire signal_10423 ;
    wire signal_10424 ;
    wire signal_10425 ;
    wire signal_10426 ;
    wire signal_10427 ;
    wire signal_10428 ;
    wire signal_10429 ;
    wire signal_10430 ;
    wire signal_10431 ;
    wire signal_10432 ;
    wire signal_10433 ;
    wire signal_10434 ;
    wire signal_10435 ;
    wire signal_10436 ;
    wire signal_10437 ;
    wire signal_10438 ;
    wire signal_10439 ;
    wire signal_10440 ;
    wire signal_10441 ;
    wire signal_10442 ;
    wire signal_10443 ;
    wire signal_10444 ;
    wire signal_10445 ;
    wire signal_10446 ;
    wire signal_10447 ;
    wire signal_10448 ;
    wire signal_10449 ;
    wire signal_10450 ;
    wire signal_10451 ;
    wire signal_10452 ;
    wire signal_10453 ;
    wire signal_10454 ;
    wire signal_10455 ;
    wire signal_10456 ;
    wire signal_10457 ;
    wire signal_10458 ;
    wire signal_10459 ;
    wire signal_10460 ;
    wire signal_10461 ;
    wire signal_10462 ;
    wire signal_10463 ;
    wire signal_10464 ;
    wire signal_10465 ;
    wire signal_10466 ;
    wire signal_10467 ;
    wire signal_10468 ;
    wire signal_10469 ;
    wire signal_10470 ;
    wire signal_10471 ;
    wire signal_10472 ;
    wire signal_10473 ;
    wire signal_10474 ;
    wire signal_10475 ;
    wire signal_10476 ;
    wire signal_10477 ;
    wire signal_10478 ;
    wire signal_10479 ;
    wire signal_10480 ;
    wire signal_10481 ;
    wire signal_10482 ;
    wire signal_10483 ;
    wire signal_10484 ;
    wire signal_10485 ;
    wire signal_10486 ;
    wire signal_10487 ;
    wire signal_10488 ;
    wire signal_10489 ;
    wire signal_10490 ;
    wire signal_10491 ;
    wire signal_10492 ;
    wire signal_10493 ;
    wire signal_10494 ;
    wire signal_10495 ;
    wire signal_10496 ;
    wire signal_10497 ;
    wire signal_10498 ;
    wire signal_10499 ;
    wire signal_10500 ;
    wire signal_10501 ;
    wire signal_10502 ;
    wire signal_10503 ;
    wire signal_10504 ;
    wire signal_10505 ;
    wire signal_10506 ;
    wire signal_10507 ;
    wire signal_10508 ;
    wire signal_10509 ;
    wire signal_10510 ;
    wire signal_10511 ;
    wire signal_10512 ;
    wire signal_10513 ;
    wire signal_10514 ;
    wire signal_10515 ;
    wire signal_10516 ;
    wire signal_10517 ;
    wire signal_10518 ;
    wire signal_10519 ;
    wire signal_10520 ;
    wire signal_10521 ;
    wire signal_10522 ;
    wire signal_10523 ;
    wire signal_10524 ;
    wire signal_10525 ;
    wire signal_10526 ;
    wire signal_10527 ;
    wire signal_10528 ;
    wire signal_10529 ;
    wire signal_10530 ;
    wire signal_10531 ;
    wire signal_10532 ;
    wire signal_10533 ;
    wire signal_10534 ;
    wire signal_10535 ;
    wire signal_10536 ;
    wire signal_10537 ;
    wire signal_10538 ;
    wire signal_10539 ;
    wire signal_10540 ;
    wire signal_10541 ;
    wire signal_10542 ;
    wire signal_10543 ;
    wire signal_10544 ;
    wire signal_10545 ;
    wire signal_10546 ;
    wire signal_10547 ;
    wire signal_10548 ;
    wire signal_10549 ;
    wire signal_10550 ;
    wire signal_10551 ;
    wire signal_10552 ;
    wire signal_10553 ;
    wire signal_10554 ;
    wire signal_10555 ;
    wire signal_10556 ;
    wire signal_10557 ;
    wire signal_10558 ;
    wire signal_10559 ;
    wire signal_10560 ;
    wire signal_10561 ;
    wire signal_10562 ;
    wire signal_10563 ;
    wire signal_10564 ;
    wire signal_10565 ;
    wire signal_10566 ;
    wire signal_10567 ;
    wire signal_10568 ;
    wire signal_10569 ;
    wire signal_10570 ;
    wire signal_10571 ;
    wire signal_10572 ;
    wire signal_10573 ;
    wire signal_10574 ;
    wire signal_10575 ;
    wire signal_10576 ;
    wire signal_10577 ;
    wire signal_10578 ;
    wire signal_10579 ;
    wire signal_10580 ;
    wire signal_10581 ;
    wire signal_10582 ;
    wire signal_10583 ;
    wire signal_10584 ;
    wire signal_10585 ;
    wire signal_10586 ;
    wire signal_10587 ;
    wire signal_10588 ;
    wire signal_10589 ;
    wire signal_10590 ;
    wire signal_10591 ;
    wire signal_10592 ;
    wire signal_10593 ;
    wire signal_10594 ;
    wire signal_10595 ;
    wire signal_10596 ;
    wire signal_10597 ;
    wire signal_10598 ;
    wire signal_10599 ;
    wire signal_10600 ;
    wire signal_10601 ;
    wire signal_10602 ;
    wire signal_10603 ;
    wire signal_10604 ;
    wire signal_10605 ;
    wire signal_10606 ;
    wire signal_10607 ;
    wire signal_10608 ;
    wire signal_10609 ;
    wire signal_10610 ;
    wire signal_10611 ;
    wire signal_10612 ;
    wire signal_10613 ;
    wire signal_10614 ;
    wire signal_10615 ;
    wire signal_10616 ;
    wire signal_10617 ;
    wire signal_10618 ;
    wire signal_10619 ;
    wire signal_10620 ;
    wire signal_10621 ;
    wire signal_10622 ;
    wire signal_10623 ;
    wire signal_10624 ;
    wire signal_10625 ;
    wire signal_10626 ;
    wire signal_10627 ;
    wire signal_10628 ;
    wire signal_10629 ;
    wire signal_10630 ;
    wire signal_10631 ;
    wire signal_10632 ;
    wire signal_10633 ;
    wire signal_10634 ;
    wire signal_10635 ;
    wire signal_10636 ;
    wire signal_10637 ;
    wire signal_10638 ;
    wire signal_10639 ;
    wire signal_10640 ;
    wire signal_10641 ;
    wire signal_10642 ;
    wire signal_10643 ;
    wire signal_10644 ;
    wire signal_10645 ;
    wire signal_10646 ;
    wire signal_10647 ;
    wire signal_10648 ;
    wire signal_10649 ;
    wire signal_10650 ;
    wire signal_10651 ;
    wire signal_10652 ;
    wire signal_10653 ;
    wire signal_10654 ;
    wire signal_10655 ;
    wire signal_10656 ;
    wire signal_10657 ;
    wire signal_10658 ;
    wire signal_10659 ;
    wire signal_10660 ;
    wire signal_10661 ;
    wire signal_10662 ;
    wire signal_10663 ;
    wire signal_10664 ;
    wire signal_10665 ;
    wire signal_10666 ;
    wire signal_10667 ;
    wire signal_10668 ;
    wire signal_10669 ;
    wire signal_10670 ;
    wire signal_10671 ;
    wire signal_10672 ;
    wire signal_10673 ;
    wire signal_10674 ;
    wire signal_10675 ;
    wire signal_10676 ;
    wire signal_10677 ;
    wire signal_10678 ;
    wire signal_10679 ;
    wire signal_10680 ;
    wire signal_10681 ;
    wire signal_10682 ;
    wire signal_10683 ;
    wire signal_10684 ;
    wire signal_10685 ;
    wire signal_10686 ;
    wire signal_10687 ;
    wire signal_10688 ;
    wire signal_10689 ;
    wire signal_10690 ;
    wire signal_10691 ;
    wire signal_10692 ;
    wire signal_10693 ;
    wire signal_10694 ;
    wire signal_10695 ;
    wire signal_10696 ;
    wire signal_10697 ;
    wire signal_10698 ;
    wire signal_10699 ;
    wire signal_10700 ;
    wire signal_10701 ;
    wire signal_10702 ;
    wire signal_10703 ;
    wire signal_10704 ;
    wire signal_10705 ;
    wire signal_10706 ;
    wire signal_10707 ;
    wire signal_10708 ;
    wire signal_10709 ;
    wire signal_10710 ;
    wire signal_10711 ;
    wire signal_10712 ;
    wire signal_10713 ;
    wire signal_10714 ;
    wire signal_10715 ;
    wire signal_10716 ;
    wire signal_10717 ;
    wire signal_10718 ;
    wire signal_10719 ;
    wire signal_10720 ;
    wire signal_10721 ;
    wire signal_10722 ;
    wire signal_10723 ;
    wire signal_10724 ;
    wire signal_10725 ;
    wire signal_10726 ;
    wire signal_10727 ;
    wire signal_10728 ;
    wire signal_10729 ;
    wire signal_10730 ;
    wire signal_10731 ;
    wire signal_10732 ;
    wire signal_10733 ;
    wire signal_10734 ;
    wire signal_10735 ;
    wire signal_10736 ;
    wire signal_10737 ;
    wire signal_10738 ;
    wire signal_10739 ;
    wire signal_10740 ;
    wire signal_10741 ;
    wire signal_10742 ;
    wire signal_10743 ;
    wire signal_10744 ;
    wire signal_10745 ;
    wire signal_10746 ;
    wire signal_10747 ;
    wire signal_10748 ;
    wire signal_10749 ;
    wire signal_10750 ;
    wire signal_10751 ;
    wire signal_10752 ;
    wire signal_10753 ;
    wire signal_10754 ;
    wire signal_10755 ;
    wire signal_10756 ;
    wire signal_10757 ;
    wire signal_10758 ;
    wire signal_10759 ;
    wire signal_10760 ;
    wire signal_10761 ;
    wire signal_10762 ;
    wire signal_10763 ;
    wire signal_10764 ;
    wire signal_10765 ;
    wire signal_10766 ;
    wire signal_10767 ;
    wire signal_10768 ;
    wire signal_10769 ;
    wire signal_10770 ;
    wire signal_10771 ;
    wire signal_10772 ;
    wire signal_10773 ;
    wire signal_10774 ;
    wire signal_10775 ;
    wire signal_10776 ;
    wire signal_10777 ;
    wire signal_10778 ;
    wire signal_10779 ;
    wire signal_10780 ;
    wire signal_10781 ;
    wire signal_10782 ;
    wire signal_10783 ;
    wire signal_10784 ;
    wire signal_10785 ;
    wire signal_10786 ;
    wire signal_10787 ;
    wire signal_10788 ;
    wire signal_10789 ;
    wire signal_10790 ;
    wire signal_10791 ;
    wire signal_10792 ;
    wire signal_10793 ;
    wire signal_10794 ;
    wire signal_10795 ;
    wire signal_10796 ;
    wire signal_10797 ;
    wire signal_10798 ;
    wire signal_10799 ;
    wire signal_10800 ;
    wire signal_10801 ;
    wire signal_10802 ;
    wire signal_10803 ;
    wire signal_10804 ;
    wire signal_10805 ;
    wire signal_10806 ;
    wire signal_10807 ;
    wire signal_10808 ;
    wire signal_10809 ;
    wire signal_10810 ;
    wire signal_10811 ;
    wire signal_10812 ;
    wire signal_10813 ;
    wire signal_10814 ;
    wire signal_10815 ;
    wire signal_10816 ;
    wire signal_10817 ;
    wire signal_10818 ;
    wire signal_10819 ;
    wire signal_10820 ;
    wire signal_10821 ;
    wire signal_10822 ;
    wire signal_10823 ;
    wire signal_10824 ;
    wire signal_10825 ;
    wire signal_10826 ;
    wire signal_10827 ;
    wire signal_10828 ;
    wire signal_10829 ;
    wire signal_10830 ;
    wire signal_10831 ;
    wire signal_10832 ;
    wire signal_10833 ;
    wire signal_10834 ;
    wire signal_10835 ;
    wire signal_10836 ;
    wire signal_10837 ;
    wire signal_10838 ;
    wire signal_10839 ;
    wire signal_10840 ;
    wire signal_10841 ;
    wire signal_10842 ;
    wire signal_10843 ;
    wire signal_10844 ;
    wire signal_10845 ;
    wire signal_10846 ;
    wire signal_10847 ;
    wire signal_10848 ;
    wire signal_10849 ;
    wire signal_10850 ;
    wire signal_10851 ;
    wire signal_10852 ;
    wire signal_10853 ;
    wire signal_10854 ;
    wire signal_10855 ;
    wire signal_10856 ;
    wire signal_10857 ;
    wire signal_10858 ;
    wire signal_10859 ;
    wire signal_10860 ;
    wire signal_10861 ;
    wire signal_10862 ;
    wire signal_10863 ;
    wire signal_10864 ;
    wire signal_10865 ;
    wire signal_10866 ;
    wire signal_10867 ;
    wire signal_10868 ;
    wire signal_10869 ;
    wire signal_10870 ;
    wire signal_10871 ;
    wire signal_10872 ;
    wire signal_10873 ;
    wire signal_10874 ;
    wire signal_10875 ;
    wire signal_10876 ;
    wire signal_10877 ;
    wire signal_10878 ;
    wire signal_10879 ;
    wire signal_10880 ;
    wire signal_10881 ;
    wire signal_10882 ;
    wire signal_10883 ;
    wire signal_10884 ;
    wire signal_10885 ;
    wire signal_10886 ;
    wire signal_10887 ;
    wire signal_10888 ;
    wire signal_10889 ;
    wire signal_10890 ;
    wire signal_10891 ;
    wire signal_10892 ;
    wire signal_10893 ;
    wire signal_10894 ;
    wire signal_10895 ;
    wire signal_10896 ;
    wire signal_10897 ;
    wire signal_10898 ;
    wire signal_10899 ;
    wire signal_10900 ;
    wire signal_10901 ;
    wire signal_10902 ;
    wire signal_10903 ;
    wire signal_10904 ;
    wire signal_10905 ;
    wire signal_10906 ;
    wire signal_10907 ;
    wire signal_10908 ;
    wire signal_10909 ;
    wire signal_10910 ;
    wire signal_10911 ;
    wire signal_10912 ;
    wire signal_10913 ;
    wire signal_10914 ;
    wire signal_10915 ;
    wire signal_10916 ;
    wire signal_10917 ;
    wire signal_10918 ;
    wire signal_10919 ;
    wire signal_10920 ;
    wire signal_10921 ;
    wire signal_10922 ;
    wire signal_10923 ;
    wire signal_10924 ;
    wire signal_10925 ;
    wire signal_10926 ;
    wire signal_10927 ;
    wire signal_10928 ;
    wire signal_10929 ;
    wire signal_10930 ;
    wire signal_10931 ;
    wire signal_10932 ;
    wire signal_10933 ;
    wire signal_10934 ;
    wire signal_10935 ;
    wire signal_10936 ;
    wire signal_10937 ;
    wire signal_10938 ;
    wire signal_10939 ;
    wire signal_10940 ;
    wire signal_10941 ;
    wire signal_10942 ;
    wire signal_10943 ;
    wire signal_10944 ;
    wire signal_10945 ;
    wire signal_10946 ;
    wire signal_10947 ;
    wire signal_10948 ;
    wire signal_10949 ;
    wire signal_10950 ;
    wire signal_10951 ;
    wire signal_10952 ;
    wire signal_10953 ;
    wire signal_10954 ;
    wire signal_10955 ;
    wire signal_10956 ;
    wire signal_10957 ;
    wire signal_10958 ;
    wire signal_10959 ;
    wire signal_10960 ;
    wire signal_10961 ;
    wire signal_10962 ;
    wire signal_10963 ;
    wire signal_10964 ;
    wire signal_10965 ;
    wire signal_10966 ;
    wire signal_10967 ;
    wire signal_10968 ;
    wire signal_10969 ;
    wire signal_10970 ;
    wire signal_10971 ;
    wire signal_10972 ;
    wire signal_10973 ;
    wire signal_10974 ;
    wire signal_10975 ;
    wire signal_10976 ;
    wire signal_10977 ;
    wire signal_10978 ;
    wire signal_10979 ;
    wire signal_10980 ;
    wire signal_10981 ;
    wire signal_10982 ;
    wire signal_10983 ;
    wire signal_10984 ;
    wire signal_10985 ;
    wire signal_10986 ;
    wire signal_10987 ;
    wire signal_10988 ;
    wire signal_10989 ;
    wire signal_10990 ;
    wire signal_10991 ;
    wire signal_10992 ;
    wire signal_10993 ;
    wire signal_10994 ;
    wire signal_10995 ;
    wire signal_10996 ;
    wire signal_10997 ;
    wire signal_10998 ;
    wire signal_10999 ;
    wire signal_11000 ;
    wire signal_11001 ;
    wire signal_11002 ;
    wire signal_11003 ;
    wire signal_11004 ;
    wire signal_11005 ;
    wire signal_11006 ;
    wire signal_11007 ;
    wire signal_11008 ;
    wire signal_11009 ;
    wire signal_11010 ;
    wire signal_11011 ;
    wire signal_11012 ;
    wire signal_11013 ;
    wire signal_11014 ;
    wire signal_11015 ;
    wire signal_11016 ;
    wire signal_11017 ;
    wire signal_11018 ;
    wire signal_11019 ;
    wire signal_11020 ;
    wire signal_11021 ;
    wire signal_11022 ;
    wire signal_11023 ;
    wire signal_11024 ;
    wire signal_11025 ;
    wire signal_11026 ;
    wire signal_11027 ;
    wire signal_11028 ;
    wire signal_11029 ;
    wire signal_11030 ;
    wire signal_11031 ;
    wire signal_11032 ;
    wire signal_11033 ;
    wire signal_11034 ;
    wire signal_11035 ;
    wire signal_11036 ;
    wire signal_11037 ;
    wire signal_11038 ;
    wire signal_11039 ;
    wire signal_11040 ;
    wire signal_11041 ;
    wire signal_11042 ;
    wire signal_11043 ;
    wire signal_11044 ;
    wire signal_11045 ;
    wire signal_11046 ;
    wire signal_11047 ;
    wire signal_11048 ;
    wire signal_11049 ;
    wire signal_11050 ;
    wire signal_11051 ;
    wire signal_11052 ;
    wire signal_11053 ;
    wire signal_11054 ;
    wire signal_11055 ;
    wire signal_11056 ;
    wire signal_11057 ;
    wire signal_11058 ;
    wire signal_11059 ;
    wire signal_11060 ;
    wire signal_11061 ;
    wire signal_11062 ;
    wire signal_11063 ;
    wire signal_11064 ;
    wire signal_11065 ;
    wire signal_11066 ;
    wire signal_11067 ;
    wire signal_11068 ;
    wire signal_11069 ;
    wire signal_11070 ;
    wire signal_11071 ;
    wire signal_11072 ;
    wire signal_11073 ;
    wire signal_11074 ;
    wire signal_11075 ;
    wire signal_11076 ;
    wire signal_11077 ;
    wire signal_11078 ;
    wire signal_11079 ;
    wire signal_11080 ;
    wire signal_11081 ;
    wire signal_11082 ;
    wire signal_11083 ;
    wire signal_11084 ;
    wire signal_11085 ;
    wire signal_11086 ;
    wire signal_11087 ;
    wire signal_11088 ;
    wire signal_11089 ;
    wire signal_11090 ;
    wire signal_11091 ;
    wire signal_11092 ;
    wire signal_11093 ;
    wire signal_11094 ;
    wire signal_11095 ;
    wire signal_11096 ;
    wire signal_11097 ;
    wire signal_11098 ;
    wire signal_11099 ;
    wire signal_11100 ;
    wire signal_11101 ;
    wire signal_11102 ;
    wire signal_11103 ;
    wire signal_11104 ;
    wire signal_11105 ;
    wire signal_11106 ;
    wire signal_11107 ;
    wire signal_11108 ;
    wire signal_11109 ;
    wire signal_11110 ;
    wire signal_11111 ;
    wire signal_11112 ;
    wire signal_11113 ;
    wire signal_11114 ;
    wire signal_11115 ;
    wire signal_11116 ;
    wire signal_11117 ;
    wire signal_11118 ;
    wire signal_11119 ;
    wire signal_11120 ;
    wire signal_11121 ;
    wire signal_11122 ;
    wire signal_11123 ;
    wire signal_11124 ;
    wire signal_11125 ;
    wire signal_11126 ;
    wire signal_11127 ;
    wire signal_11128 ;
    wire signal_11129 ;
    wire signal_11130 ;
    wire signal_11131 ;
    wire signal_11132 ;
    wire signal_11133 ;
    wire signal_11134 ;
    wire signal_11135 ;
    wire signal_11136 ;
    wire signal_11137 ;
    wire signal_11138 ;
    wire signal_11139 ;
    wire signal_11140 ;
    wire signal_11141 ;
    wire signal_11142 ;
    wire signal_11143 ;
    wire signal_11144 ;
    wire signal_11145 ;
    wire signal_11146 ;
    wire signal_11147 ;
    wire signal_11148 ;
    wire signal_11149 ;
    wire signal_11150 ;
    wire signal_11151 ;
    wire signal_11152 ;
    wire signal_11153 ;
    wire signal_11154 ;
    wire signal_11155 ;
    wire signal_11156 ;
    wire signal_11157 ;
    wire signal_11158 ;
    wire signal_11159 ;
    wire signal_11160 ;
    wire signal_11161 ;
    wire signal_11162 ;
    wire signal_11163 ;
    wire signal_11164 ;
    wire signal_11165 ;
    wire signal_11166 ;
    wire signal_11167 ;
    wire signal_11168 ;
    wire signal_11169 ;
    wire signal_11170 ;
    wire signal_11171 ;
    wire signal_11172 ;
    wire signal_11173 ;
    wire signal_11174 ;
    wire signal_11175 ;
    wire signal_11176 ;
    wire signal_11177 ;
    wire signal_11178 ;
    wire signal_11179 ;
    wire signal_11180 ;
    wire signal_11181 ;
    wire signal_11182 ;
    wire signal_11183 ;
    wire signal_11184 ;
    wire signal_11185 ;
    wire signal_11186 ;
    wire signal_11187 ;
    wire signal_11188 ;
    wire signal_11189 ;
    wire signal_11190 ;
    wire signal_11191 ;
    wire signal_11192 ;
    wire signal_11193 ;
    wire signal_11194 ;
    wire signal_11195 ;
    wire signal_11196 ;
    wire signal_11197 ;
    wire signal_11198 ;
    wire signal_11199 ;
    wire signal_11200 ;
    wire signal_11201 ;
    wire signal_11202 ;
    wire signal_11203 ;
    wire signal_11204 ;
    wire signal_11205 ;
    wire signal_11206 ;
    wire signal_11207 ;
    wire signal_11208 ;
    wire signal_11209 ;
    wire signal_11210 ;
    wire signal_11211 ;
    wire signal_11212 ;
    wire signal_11213 ;
    wire signal_11214 ;
    wire signal_11215 ;
    wire signal_11216 ;
    wire signal_11217 ;
    wire signal_11218 ;
    wire signal_11219 ;
    wire signal_11220 ;
    wire signal_11221 ;
    wire signal_11222 ;
    wire signal_11223 ;
    wire signal_11224 ;
    wire signal_11225 ;
    wire signal_11226 ;
    wire signal_11227 ;
    wire signal_11228 ;
    wire signal_11229 ;
    wire signal_11230 ;
    wire signal_11231 ;
    wire signal_11232 ;
    wire signal_11233 ;
    wire signal_11234 ;
    wire signal_11235 ;
    wire signal_11236 ;
    wire signal_11237 ;
    wire signal_11238 ;
    wire signal_11239 ;
    wire signal_11240 ;
    wire signal_11241 ;
    wire signal_11242 ;
    wire signal_11243 ;
    wire signal_11244 ;
    wire signal_11245 ;
    wire signal_11246 ;
    wire signal_11247 ;
    wire signal_11248 ;
    wire signal_11249 ;
    wire signal_11250 ;
    wire signal_11251 ;
    wire signal_11252 ;
    wire signal_11253 ;
    wire signal_11254 ;
    wire signal_11255 ;
    wire signal_11256 ;
    wire signal_11257 ;
    wire signal_11258 ;
    wire signal_11259 ;
    wire signal_11260 ;
    wire signal_11261 ;
    wire signal_11262 ;
    wire signal_11263 ;
    wire signal_11264 ;
    wire signal_11265 ;
    wire signal_11266 ;
    wire signal_11267 ;
    wire signal_11268 ;
    wire signal_11269 ;
    wire signal_11270 ;
    wire signal_11271 ;
    wire signal_11272 ;
    wire signal_11273 ;
    wire signal_11274 ;
    wire signal_11275 ;
    wire signal_11276 ;
    wire signal_11277 ;
    wire signal_11278 ;
    wire signal_11279 ;
    wire signal_11280 ;
    wire signal_11281 ;
    wire signal_11282 ;
    wire signal_11283 ;
    wire signal_11284 ;
    wire signal_11285 ;
    wire signal_11286 ;
    wire signal_11287 ;
    wire signal_11288 ;
    wire signal_11289 ;
    wire signal_11290 ;
    wire signal_11291 ;
    wire signal_11292 ;
    wire signal_11293 ;
    wire signal_11294 ;
    wire signal_11295 ;
    wire signal_11296 ;
    wire signal_11297 ;
    wire signal_11298 ;
    wire signal_11299 ;
    wire signal_11300 ;
    wire signal_11301 ;
    wire signal_11302 ;
    wire signal_11303 ;
    wire signal_11304 ;
    wire signal_11305 ;
    wire signal_11306 ;
    wire signal_11307 ;
    wire signal_11308 ;
    wire signal_11309 ;
    wire signal_11310 ;
    wire signal_11311 ;
    wire signal_11312 ;
    wire signal_11313 ;
    wire signal_11314 ;
    wire signal_11315 ;
    wire signal_11316 ;
    wire signal_11317 ;
    wire signal_11318 ;
    wire signal_11319 ;
    wire signal_11320 ;
    wire signal_11321 ;
    wire signal_11322 ;
    wire signal_11323 ;
    wire signal_11324 ;
    wire signal_11325 ;
    wire signal_11326 ;
    wire signal_11327 ;
    wire signal_11328 ;
    wire signal_11329 ;
    wire signal_11330 ;
    wire signal_11331 ;
    wire signal_11332 ;
    wire signal_11333 ;
    wire signal_11334 ;
    wire signal_11335 ;
    wire signal_11336 ;
    wire signal_11337 ;
    wire signal_11338 ;
    wire signal_11339 ;
    wire signal_11340 ;
    wire signal_11341 ;
    wire signal_11342 ;
    wire signal_11343 ;
    wire signal_11344 ;
    wire signal_11345 ;
    wire signal_11346 ;
    wire signal_11347 ;
    wire signal_11348 ;
    wire signal_11349 ;
    wire signal_11350 ;
    wire signal_11351 ;
    wire signal_11352 ;
    wire signal_11353 ;
    wire signal_11354 ;
    wire signal_11355 ;
    wire signal_11356 ;
    wire signal_11357 ;
    wire signal_11358 ;
    wire signal_11359 ;
    wire signal_11360 ;
    wire signal_11361 ;
    wire signal_11362 ;
    wire signal_11363 ;
    wire signal_11364 ;
    wire signal_11365 ;
    wire signal_11366 ;
    wire signal_11367 ;
    wire signal_11368 ;
    wire signal_11369 ;
    wire signal_11370 ;
    wire signal_11371 ;
    wire signal_11372 ;
    wire signal_11373 ;
    wire signal_11374 ;
    wire signal_11375 ;
    wire signal_11376 ;
    wire signal_11377 ;
    wire signal_11378 ;
    wire signal_11379 ;
    wire signal_11380 ;
    wire signal_11381 ;
    wire signal_11382 ;
    wire signal_11383 ;
    wire signal_11384 ;
    wire signal_11385 ;
    wire signal_11386 ;
    wire signal_11387 ;
    wire signal_11388 ;
    wire signal_11389 ;
    wire signal_11390 ;
    wire signal_11391 ;
    wire signal_11392 ;
    wire signal_11393 ;
    wire signal_11394 ;
    wire signal_11395 ;
    wire signal_11396 ;
    wire signal_11397 ;
    wire signal_11398 ;
    wire signal_11399 ;
    wire signal_11400 ;
    wire signal_11401 ;
    wire signal_11402 ;
    wire signal_11403 ;
    wire signal_11404 ;
    wire signal_11405 ;
    wire signal_11406 ;
    wire signal_11407 ;
    wire signal_11408 ;
    wire signal_11409 ;
    wire signal_11410 ;
    wire signal_11411 ;
    wire signal_11412 ;
    wire signal_11413 ;
    wire signal_11414 ;
    wire signal_11415 ;
    wire signal_11416 ;
    wire signal_11417 ;
    wire signal_11418 ;
    wire signal_11419 ;
    wire signal_11420 ;
    wire signal_11421 ;
    wire signal_11422 ;
    wire signal_11423 ;
    wire signal_11424 ;
    wire signal_11425 ;
    wire signal_11426 ;
    wire signal_11427 ;
    wire signal_11428 ;
    wire signal_11429 ;
    wire signal_11430 ;
    wire signal_11431 ;
    wire signal_11432 ;
    wire signal_11433 ;
    wire signal_11434 ;
    wire signal_11435 ;
    wire signal_11436 ;
    wire signal_11437 ;
    wire signal_11438 ;
    wire signal_11439 ;
    wire signal_11440 ;
    wire signal_11441 ;
    wire signal_11442 ;
    wire signal_11443 ;
    wire signal_11444 ;
    wire signal_11445 ;
    wire signal_11446 ;
    wire signal_11447 ;
    wire signal_11448 ;
    wire signal_11449 ;
    wire signal_11450 ;
    wire signal_11451 ;
    wire signal_11452 ;
    wire signal_11453 ;
    wire signal_11454 ;
    wire signal_11455 ;
    wire signal_11456 ;
    wire signal_11457 ;
    wire signal_11458 ;
    wire signal_11459 ;
    wire signal_11460 ;
    wire signal_11461 ;
    wire signal_11462 ;
    wire signal_11463 ;
    wire signal_11464 ;
    wire signal_11465 ;
    wire signal_11466 ;
    wire signal_11467 ;
    wire signal_11468 ;
    wire signal_11469 ;
    wire signal_11470 ;
    wire signal_11471 ;
    wire signal_11472 ;
    wire signal_11473 ;
    wire signal_11474 ;
    wire signal_11475 ;
    wire signal_11476 ;
    wire signal_11477 ;
    wire signal_11478 ;
    wire signal_11479 ;
    wire signal_11480 ;
    wire signal_11481 ;
    wire signal_11482 ;
    wire signal_11483 ;
    wire signal_11484 ;
    wire signal_11485 ;
    wire signal_11486 ;
    wire signal_11487 ;
    wire signal_11488 ;
    wire signal_11489 ;
    wire signal_11490 ;
    wire signal_11491 ;
    wire signal_11492 ;
    wire signal_11493 ;
    wire signal_11494 ;
    wire signal_11495 ;
    wire signal_11496 ;
    wire signal_11497 ;
    wire signal_11498 ;
    wire signal_11499 ;
    wire signal_11500 ;
    wire signal_11501 ;
    wire signal_11502 ;
    wire signal_11503 ;
    wire signal_11504 ;
    wire signal_11505 ;
    wire signal_11506 ;
    wire signal_11507 ;
    wire signal_11508 ;
    wire signal_11509 ;
    wire signal_11510 ;
    wire signal_11511 ;
    wire signal_11512 ;
    wire signal_11513 ;
    wire signal_11514 ;
    wire signal_11515 ;
    wire signal_11516 ;
    wire signal_11517 ;
    wire signal_11518 ;
    wire signal_11519 ;
    wire signal_11520 ;
    wire signal_11521 ;
    wire signal_11522 ;
    wire signal_11523 ;
    wire signal_11524 ;
    wire signal_11525 ;
    wire signal_11526 ;
    wire signal_11527 ;
    wire signal_11528 ;
    wire signal_11529 ;
    wire signal_11530 ;
    wire signal_11531 ;
    wire signal_11532 ;
    wire signal_11533 ;
    wire signal_11534 ;
    wire signal_11535 ;
    wire signal_11536 ;
    wire signal_11537 ;
    wire signal_11538 ;
    wire signal_11539 ;
    wire signal_11540 ;
    wire signal_11541 ;
    wire signal_11542 ;
    wire signal_11543 ;
    wire signal_11544 ;
    wire signal_11545 ;
    wire signal_11546 ;
    wire signal_11547 ;
    wire signal_11548 ;
    wire signal_11549 ;
    wire signal_11550 ;
    wire signal_11551 ;
    wire signal_11552 ;
    wire signal_11553 ;
    wire signal_11554 ;
    wire signal_11555 ;
    wire signal_11556 ;
    wire signal_11557 ;
    wire signal_11558 ;
    wire signal_11559 ;
    wire signal_11560 ;
    wire signal_11561 ;
    wire signal_11562 ;
    wire signal_11563 ;
    wire signal_11564 ;
    wire signal_11565 ;
    wire signal_11566 ;
    wire signal_11567 ;
    wire signal_11568 ;
    wire signal_11569 ;
    wire signal_11570 ;
    wire signal_11571 ;
    wire signal_11572 ;
    wire signal_11573 ;
    wire signal_11574 ;
    wire signal_11575 ;
    wire signal_11576 ;
    wire signal_11577 ;
    wire signal_11578 ;
    wire signal_11579 ;
    wire signal_11580 ;
    wire signal_11581 ;
    wire signal_11582 ;
    wire signal_11583 ;
    wire signal_11584 ;
    wire signal_11585 ;
    wire signal_11586 ;
    wire signal_11587 ;
    wire signal_11588 ;
    wire signal_11589 ;
    wire signal_11590 ;
    wire signal_11591 ;
    wire signal_11592 ;
    wire signal_11593 ;
    wire signal_11594 ;
    wire signal_11595 ;
    wire signal_11596 ;
    wire signal_11597 ;
    wire signal_11598 ;
    wire signal_11599 ;
    wire signal_11600 ;
    wire signal_11601 ;
    wire signal_11602 ;
    wire signal_11603 ;
    wire signal_11604 ;
    wire signal_11605 ;
    wire signal_11606 ;
    wire signal_11607 ;
    wire signal_11608 ;
    wire signal_11609 ;
    wire signal_11610 ;
    wire signal_11611 ;
    wire signal_11612 ;
    wire signal_11613 ;
    wire signal_11614 ;
    wire signal_11615 ;
    wire signal_11616 ;
    wire signal_11617 ;
    wire signal_11618 ;
    wire signal_11619 ;
    wire signal_11620 ;
    wire signal_11621 ;
    wire signal_11622 ;
    wire signal_11623 ;
    wire signal_11624 ;
    wire signal_11625 ;
    wire signal_11626 ;
    wire signal_11627 ;
    wire signal_11628 ;
    wire signal_11629 ;
    wire signal_11630 ;
    wire signal_11631 ;
    wire signal_11632 ;
    wire signal_11633 ;
    wire signal_11634 ;
    wire signal_11635 ;
    wire signal_11636 ;
    wire signal_11637 ;
    wire signal_11638 ;
    wire signal_11639 ;
    wire signal_11640 ;
    wire signal_11641 ;
    wire signal_11642 ;
    wire signal_11643 ;
    wire signal_11644 ;
    wire signal_11645 ;
    wire signal_11646 ;
    wire signal_11647 ;
    wire signal_11648 ;
    wire signal_11649 ;
    wire signal_11650 ;
    wire signal_11651 ;
    wire signal_11652 ;
    wire signal_11653 ;
    wire signal_11654 ;
    wire signal_11655 ;
    wire signal_11656 ;
    wire signal_11657 ;
    wire signal_11658 ;
    wire signal_11659 ;
    wire signal_11660 ;
    wire signal_11661 ;
    wire signal_11662 ;
    wire signal_11663 ;
    wire signal_11664 ;
    wire signal_11665 ;
    wire signal_11666 ;
    wire signal_11667 ;
    wire signal_11668 ;
    wire signal_11669 ;
    wire signal_11670 ;
    wire signal_11671 ;
    wire signal_11672 ;
    wire signal_11673 ;
    wire signal_11674 ;
    wire signal_11675 ;
    wire signal_11676 ;
    wire signal_11677 ;
    wire signal_11678 ;
    wire signal_11679 ;
    wire signal_11680 ;
    wire signal_11681 ;
    wire signal_11682 ;
    wire signal_11683 ;
    wire signal_11684 ;
    wire signal_11685 ;
    wire signal_11686 ;
    wire signal_11687 ;
    wire signal_11688 ;
    wire signal_11689 ;
    wire signal_11690 ;
    wire signal_11691 ;
    wire signal_11692 ;
    wire signal_11693 ;
    wire signal_11694 ;
    wire signal_11695 ;
    wire signal_11696 ;
    wire signal_11697 ;
    wire signal_11698 ;
    wire signal_11699 ;
    wire signal_11700 ;
    wire signal_11701 ;
    wire signal_11702 ;
    wire signal_11703 ;
    wire signal_11704 ;
    wire signal_11705 ;
    wire signal_11706 ;
    wire signal_11707 ;
    wire signal_11708 ;
    wire signal_11709 ;
    wire signal_11710 ;
    wire signal_11711 ;
    wire signal_11712 ;
    wire signal_11713 ;
    wire signal_11714 ;
    wire signal_11715 ;
    wire signal_11716 ;
    wire signal_11717 ;
    wire signal_11718 ;
    wire signal_11719 ;
    wire signal_11720 ;
    wire signal_11721 ;
    wire signal_11722 ;
    wire signal_11723 ;
    wire signal_11724 ;
    wire signal_11725 ;
    wire signal_11726 ;
    wire signal_11727 ;
    wire signal_11728 ;
    wire signal_11729 ;
    wire signal_11730 ;
    wire signal_11731 ;
    wire signal_11732 ;
    wire signal_11733 ;
    wire signal_11734 ;
    wire signal_11735 ;
    wire signal_11736 ;
    wire signal_11737 ;
    wire signal_11738 ;
    wire signal_11739 ;
    wire signal_11740 ;
    wire signal_11741 ;
    wire signal_11742 ;
    wire signal_11743 ;
    wire signal_11744 ;
    wire signal_11745 ;
    wire signal_11746 ;
    wire signal_11747 ;
    wire signal_11748 ;
    wire signal_11749 ;
    wire signal_11750 ;
    wire signal_11751 ;
    wire signal_11752 ;
    wire signal_11753 ;
    wire signal_11754 ;
    wire signal_11755 ;
    wire signal_11756 ;
    wire signal_11757 ;
    wire signal_11758 ;
    wire signal_11759 ;
    wire signal_11760 ;
    wire signal_11761 ;
    wire signal_11762 ;
    wire signal_11763 ;
    wire signal_11764 ;
    wire signal_11765 ;
    wire signal_11766 ;
    wire signal_11767 ;
    wire signal_11768 ;
    wire signal_11769 ;
    wire signal_11770 ;
    wire signal_11771 ;
    wire signal_11772 ;
    wire signal_11773 ;
    wire signal_11774 ;
    wire signal_11775 ;
    wire signal_11776 ;
    wire signal_11777 ;
    wire signal_11778 ;
    wire signal_11779 ;
    wire signal_11780 ;
    wire signal_11781 ;
    wire signal_11782 ;
    wire signal_11783 ;
    wire signal_11784 ;
    wire signal_11785 ;
    wire signal_11786 ;
    wire signal_11787 ;
    wire signal_11788 ;
    wire signal_11789 ;
    wire signal_11790 ;
    wire signal_11791 ;
    wire signal_11792 ;
    wire signal_11793 ;
    wire signal_11794 ;
    wire signal_11795 ;
    wire signal_11796 ;
    wire signal_11797 ;
    wire signal_11798 ;
    wire signal_11799 ;
    wire signal_11800 ;
    wire signal_11801 ;
    wire signal_11802 ;
    wire signal_11803 ;
    wire signal_11804 ;
    wire signal_11805 ;
    wire signal_11806 ;
    wire signal_11807 ;
    wire signal_11808 ;
    wire signal_11809 ;
    wire signal_11810 ;
    wire signal_11811 ;
    wire signal_11812 ;
    wire signal_11813 ;
    wire signal_11814 ;
    wire signal_11815 ;
    wire signal_11816 ;
    wire signal_11817 ;
    wire signal_11818 ;
    wire signal_11819 ;
    wire signal_11820 ;
    wire signal_11821 ;
    wire signal_11822 ;
    wire signal_11823 ;
    wire signal_11824 ;
    wire signal_11825 ;
    wire signal_11826 ;
    wire signal_11827 ;
    wire signal_11828 ;
    wire signal_11829 ;
    wire signal_11830 ;
    wire signal_11831 ;
    wire signal_11832 ;
    wire signal_11833 ;
    wire signal_11834 ;
    wire signal_11835 ;
    wire signal_11836 ;
    wire signal_11837 ;
    wire signal_11838 ;
    wire signal_11839 ;
    wire signal_11840 ;
    wire signal_11841 ;
    wire signal_11842 ;
    wire signal_11843 ;
    wire signal_11844 ;
    wire signal_11845 ;
    wire signal_11846 ;
    wire signal_11847 ;
    wire signal_11848 ;
    wire signal_11849 ;
    wire signal_11850 ;
    wire signal_11851 ;
    wire signal_11852 ;
    wire signal_11853 ;
    wire signal_11854 ;
    wire signal_11855 ;
    wire signal_11856 ;
    wire signal_11857 ;
    wire signal_11858 ;
    wire signal_11859 ;
    wire signal_11860 ;
    wire signal_11861 ;
    wire signal_11862 ;
    wire signal_11863 ;
    wire signal_11864 ;
    wire signal_11865 ;
    wire signal_11866 ;
    wire signal_11867 ;
    wire signal_11868 ;
    wire signal_11869 ;
    wire signal_11870 ;
    wire signal_11871 ;
    wire signal_11872 ;
    wire signal_11873 ;
    wire signal_11874 ;
    wire signal_11875 ;
    wire signal_11876 ;
    wire signal_11877 ;
    wire signal_11878 ;
    wire signal_11879 ;
    wire signal_11880 ;
    wire signal_11881 ;
    wire signal_11882 ;
    wire signal_11883 ;
    wire signal_11884 ;
    wire signal_11885 ;
    wire signal_11886 ;
    wire signal_11887 ;
    wire signal_11888 ;
    wire signal_11889 ;
    wire signal_11890 ;
    wire signal_11891 ;
    wire signal_11892 ;
    wire signal_11893 ;
    wire signal_11894 ;
    wire signal_11895 ;
    wire signal_11896 ;
    wire signal_11897 ;
    wire signal_11898 ;
    wire signal_11899 ;
    wire signal_11900 ;
    wire signal_11901 ;
    wire signal_11902 ;
    wire signal_11903 ;
    wire signal_11904 ;
    wire signal_11905 ;
    wire signal_11906 ;
    wire signal_11907 ;
    wire signal_11908 ;
    wire signal_11909 ;
    wire signal_11910 ;
    wire signal_11911 ;
    wire signal_11912 ;
    wire signal_11913 ;
    wire signal_11914 ;
    wire signal_11915 ;
    wire signal_11916 ;
    wire signal_11917 ;
    wire signal_11918 ;
    wire signal_11919 ;
    wire signal_11920 ;
    wire signal_11921 ;
    wire signal_11922 ;
    wire signal_11923 ;
    wire signal_11924 ;
    wire signal_11925 ;
    wire signal_11926 ;
    wire signal_11927 ;
    wire signal_11928 ;
    wire signal_11929 ;
    wire signal_11930 ;
    wire signal_11931 ;
    wire signal_11932 ;
    wire signal_11933 ;
    wire signal_11934 ;
    wire signal_11935 ;
    wire signal_11936 ;
    wire signal_11937 ;
    wire signal_11938 ;
    wire signal_11939 ;
    wire signal_11940 ;
    wire signal_11941 ;
    wire signal_11942 ;
    wire signal_11943 ;
    wire signal_11944 ;
    wire signal_11945 ;
    wire signal_11946 ;
    wire signal_11947 ;
    wire signal_11948 ;
    wire signal_11949 ;
    wire signal_11950 ;
    wire signal_11951 ;
    wire signal_11952 ;
    wire signal_11953 ;
    wire signal_11954 ;
    wire signal_11955 ;
    wire signal_11956 ;
    wire signal_11957 ;
    wire signal_11958 ;
    wire signal_11959 ;
    wire signal_11960 ;
    wire signal_11961 ;
    wire signal_11962 ;
    wire signal_11963 ;
    wire signal_11964 ;
    wire signal_11965 ;
    wire signal_11966 ;
    wire signal_11967 ;
    wire signal_11968 ;
    wire signal_11969 ;
    wire signal_11970 ;
    wire signal_11971 ;
    wire signal_11972 ;
    wire signal_11973 ;
    wire signal_11974 ;
    wire signal_11975 ;
    wire signal_11976 ;
    wire signal_11977 ;
    wire signal_11978 ;
    wire signal_11979 ;
    wire signal_11980 ;
    wire signal_11981 ;
    wire signal_11982 ;
    wire signal_11983 ;
    wire signal_11984 ;
    wire signal_11985 ;
    wire signal_11986 ;
    wire signal_11987 ;
    wire signal_11988 ;
    wire signal_11989 ;
    wire signal_11990 ;
    wire signal_11991 ;
    wire signal_11992 ;
    wire signal_11993 ;
    wire signal_11994 ;
    wire signal_11995 ;
    wire signal_11996 ;
    wire signal_11997 ;
    wire signal_11998 ;
    wire signal_11999 ;
    wire signal_12000 ;
    wire signal_12001 ;
    wire signal_12002 ;
    wire signal_12003 ;
    wire signal_12004 ;
    wire signal_12005 ;
    wire signal_12006 ;
    wire signal_12007 ;
    wire signal_12008 ;
    wire signal_12009 ;
    wire signal_12010 ;
    wire signal_12011 ;
    wire signal_12012 ;
    wire signal_12013 ;
    wire signal_12014 ;
    wire signal_12015 ;
    wire signal_12016 ;
    wire signal_12017 ;
    wire signal_12018 ;
    wire signal_12019 ;
    wire signal_12020 ;
    wire signal_12021 ;
    wire signal_12022 ;
    wire signal_12023 ;
    wire signal_12024 ;
    wire signal_12025 ;
    wire signal_12026 ;
    wire signal_12027 ;
    wire signal_12028 ;
    wire signal_12029 ;
    wire signal_12030 ;
    wire signal_12031 ;
    wire signal_12032 ;
    wire signal_12033 ;
    wire signal_12034 ;
    wire signal_12035 ;
    wire signal_12036 ;
    wire signal_12037 ;
    wire signal_12038 ;
    wire signal_12039 ;
    wire signal_12040 ;
    wire signal_12041 ;
    wire signal_12042 ;
    wire signal_12043 ;
    wire signal_12044 ;
    wire signal_12045 ;
    wire signal_12046 ;
    wire signal_12047 ;
    wire signal_12048 ;
    wire signal_12049 ;
    wire signal_12050 ;
    wire signal_12051 ;
    wire signal_12052 ;
    wire signal_12053 ;
    wire signal_12054 ;
    wire signal_12055 ;
    wire signal_12056 ;
    wire signal_12057 ;
    wire signal_12058 ;
    wire signal_12059 ;
    wire signal_12060 ;
    wire signal_12061 ;
    wire signal_12062 ;
    wire signal_12063 ;
    wire signal_12064 ;
    wire signal_12065 ;
    wire signal_12066 ;
    wire signal_12067 ;
    wire signal_12068 ;
    wire signal_12069 ;
    wire signal_12070 ;
    wire signal_12071 ;
    wire signal_12072 ;
    wire signal_12073 ;
    wire signal_12074 ;
    wire signal_12075 ;
    wire signal_12076 ;
    wire signal_12077 ;
    wire signal_12078 ;
    wire signal_12079 ;
    wire signal_12080 ;
    wire signal_12081 ;
    wire signal_12082 ;
    wire signal_12083 ;
    wire signal_12084 ;
    wire signal_12085 ;
    wire signal_12086 ;
    wire signal_12087 ;
    wire signal_12088 ;
    wire signal_12089 ;
    wire signal_12090 ;
    wire signal_12091 ;
    wire signal_12092 ;
    wire signal_12093 ;
    wire signal_12094 ;
    wire signal_12095 ;
    wire signal_12096 ;
    wire signal_12097 ;
    wire signal_12098 ;
    wire signal_12099 ;
    wire signal_12100 ;
    wire signal_12101 ;
    wire signal_12102 ;
    wire signal_12103 ;
    wire signal_12104 ;
    wire signal_12105 ;
    wire signal_12106 ;
    wire signal_12107 ;
    wire signal_12108 ;
    wire signal_12109 ;
    wire signal_12110 ;
    wire signal_12111 ;
    wire signal_12112 ;
    wire signal_12113 ;
    wire signal_12114 ;
    wire signal_12115 ;
    wire signal_12116 ;
    wire signal_12117 ;
    wire signal_12118 ;
    wire signal_12119 ;
    wire signal_12120 ;
    wire signal_12121 ;
    wire signal_12122 ;
    wire signal_12123 ;
    wire signal_12124 ;
    wire signal_12125 ;
    wire signal_12126 ;
    wire signal_12127 ;
    wire signal_12128 ;
    wire signal_12129 ;
    wire signal_12130 ;
    wire signal_12131 ;
    wire signal_12132 ;
    wire signal_12133 ;
    wire signal_12134 ;
    wire signal_12135 ;
    wire signal_12136 ;
    wire signal_12137 ;
    wire signal_12138 ;
    wire signal_12139 ;
    wire signal_12140 ;
    wire signal_12141 ;
    wire signal_12142 ;
    wire signal_12143 ;
    wire signal_12144 ;
    wire signal_12145 ;
    wire signal_12146 ;
    wire signal_12147 ;
    wire signal_12148 ;
    wire signal_12149 ;
    wire signal_12150 ;
    wire signal_12151 ;
    wire signal_12152 ;
    wire signal_12153 ;
    wire signal_12154 ;
    wire signal_12155 ;
    wire signal_12156 ;
    wire signal_12157 ;
    wire signal_12158 ;
    wire signal_12159 ;
    wire signal_12160 ;
    wire signal_12161 ;
    wire signal_12162 ;
    wire signal_12163 ;
    wire signal_12164 ;
    wire signal_12165 ;
    wire signal_12166 ;
    wire signal_12167 ;
    wire signal_12168 ;
    wire signal_12169 ;
    wire signal_12170 ;
    wire signal_12171 ;
    wire signal_12172 ;
    wire signal_12173 ;
    wire signal_12174 ;
    wire signal_12175 ;
    wire signal_12176 ;
    wire signal_12177 ;
    wire signal_12178 ;
    wire signal_12179 ;
    wire signal_12180 ;
    wire signal_12181 ;
    wire signal_12182 ;
    wire signal_12183 ;
    wire signal_12184 ;
    wire signal_12185 ;
    wire signal_12186 ;
    wire signal_12187 ;
    wire signal_12188 ;
    wire signal_12189 ;
    wire signal_12190 ;
    wire signal_12191 ;
    wire signal_12192 ;
    wire signal_12193 ;
    wire signal_12194 ;
    wire signal_12195 ;
    wire signal_12196 ;
    wire signal_12197 ;
    wire signal_12198 ;
    wire signal_12199 ;
    wire signal_12200 ;
    wire signal_12201 ;
    wire signal_12202 ;
    wire signal_12203 ;
    wire signal_12204 ;
    wire signal_12205 ;
    wire signal_12206 ;
    wire signal_12207 ;
    wire signal_12208 ;
    wire signal_12209 ;
    wire signal_12210 ;
    wire signal_12211 ;
    wire signal_12212 ;
    wire signal_12213 ;
    wire signal_12214 ;
    wire signal_12215 ;
    wire signal_12216 ;
    wire signal_12217 ;
    wire signal_12218 ;
    wire signal_12219 ;
    wire signal_12220 ;
    wire signal_12221 ;
    wire signal_12222 ;
    wire signal_12223 ;
    wire signal_12224 ;
    wire signal_12225 ;
    wire signal_12226 ;
    wire signal_12227 ;
    wire signal_12228 ;
    wire signal_12229 ;
    wire signal_12230 ;
    wire signal_12231 ;
    wire signal_12232 ;
    wire signal_12233 ;
    wire signal_12234 ;
    wire signal_12235 ;
    wire signal_12236 ;
    wire signal_12237 ;
    wire signal_12238 ;
    wire signal_12239 ;
    wire signal_12240 ;
    wire signal_12241 ;
    wire signal_12242 ;
    wire signal_12243 ;
    wire signal_12244 ;
    wire signal_12245 ;
    wire signal_12246 ;
    wire signal_12247 ;
    wire signal_12248 ;
    wire signal_12249 ;
    wire signal_12250 ;
    wire signal_12251 ;
    wire signal_12252 ;
    wire signal_12253 ;
    wire signal_12254 ;
    wire signal_12255 ;
    wire signal_12256 ;
    wire signal_12257 ;
    wire signal_12258 ;
    wire signal_12259 ;
    wire signal_12260 ;
    wire signal_12261 ;
    wire signal_12262 ;
    wire signal_12263 ;
    wire signal_12264 ;
    wire signal_12265 ;
    wire signal_12266 ;
    wire signal_12267 ;
    wire signal_12268 ;
    wire signal_12269 ;
    wire signal_12270 ;
    wire signal_12271 ;
    wire signal_12272 ;
    wire signal_12273 ;
    wire signal_12274 ;
    wire signal_12275 ;
    wire signal_12276 ;
    wire signal_12277 ;
    wire signal_12278 ;
    wire signal_12279 ;
    wire signal_12280 ;
    wire signal_12281 ;
    wire signal_12282 ;
    wire signal_12283 ;
    wire signal_12284 ;
    wire signal_12285 ;
    wire signal_12286 ;
    wire signal_12287 ;
    wire signal_12288 ;
    wire signal_12289 ;
    wire signal_12290 ;
    wire signal_12291 ;
    wire signal_12292 ;
    wire signal_12293 ;
    wire signal_12294 ;
    wire signal_12295 ;
    wire signal_12296 ;
    wire signal_12297 ;
    wire signal_12298 ;
    wire signal_12299 ;
    wire signal_12300 ;
    wire signal_12301 ;
    wire signal_12302 ;
    wire signal_12303 ;
    wire signal_12304 ;
    wire signal_12305 ;
    wire signal_12306 ;
    wire signal_12307 ;
    wire signal_12308 ;
    wire signal_12309 ;
    wire signal_12310 ;
    wire signal_12311 ;
    wire signal_12312 ;
    wire signal_12313 ;
    wire signal_12314 ;
    wire signal_12315 ;
    wire signal_12316 ;
    wire signal_12317 ;
    wire signal_12318 ;
    wire signal_12319 ;
    wire signal_12320 ;
    wire signal_12321 ;
    wire signal_12322 ;
    wire signal_12323 ;
    wire signal_12324 ;
    wire signal_12325 ;
    wire signal_12326 ;
    wire signal_12327 ;
    wire signal_12328 ;
    wire signal_12329 ;
    wire signal_12330 ;
    wire signal_12331 ;
    wire signal_12332 ;
    wire signal_12333 ;
    wire signal_12334 ;
    wire signal_12335 ;
    wire signal_12336 ;
    wire signal_12337 ;
    wire signal_12338 ;
    wire signal_12339 ;
    wire signal_12340 ;
    wire signal_12341 ;
    wire signal_12342 ;
    wire signal_12343 ;
    wire signal_12344 ;
    wire signal_12345 ;
    wire signal_12346 ;
    wire signal_12347 ;
    wire signal_12348 ;
    wire signal_12349 ;
    wire signal_12350 ;
    wire signal_12351 ;
    wire signal_12352 ;
    wire signal_12353 ;
    wire signal_12354 ;
    wire signal_12355 ;
    wire signal_12356 ;
    wire signal_12357 ;
    wire signal_12358 ;
    wire signal_12359 ;
    wire signal_12360 ;
    wire signal_12361 ;
    wire signal_12362 ;
    wire signal_12363 ;
    wire signal_12364 ;
    wire signal_12365 ;
    wire signal_12366 ;
    wire signal_12367 ;
    wire signal_12368 ;
    wire signal_12369 ;
    wire signal_12370 ;
    wire signal_12371 ;
    wire signal_12372 ;
    wire signal_12373 ;
    wire signal_12374 ;
    wire signal_12375 ;
    wire signal_12376 ;
    wire signal_12377 ;
    wire signal_12378 ;
    wire signal_12379 ;
    wire signal_12380 ;
    wire signal_12381 ;
    wire signal_12382 ;
    wire signal_12383 ;
    wire signal_12384 ;
    wire signal_12385 ;
    wire signal_12386 ;
    wire signal_12387 ;
    wire signal_12388 ;
    wire signal_12389 ;
    wire signal_12390 ;
    wire signal_12391 ;
    wire signal_12392 ;
    wire signal_12393 ;
    wire signal_12394 ;
    wire signal_12395 ;
    wire signal_12396 ;
    wire signal_12397 ;
    wire signal_12398 ;
    wire signal_12399 ;
    wire signal_12400 ;
    wire signal_12401 ;
    wire signal_12402 ;
    wire signal_12403 ;
    wire signal_12404 ;
    wire signal_12405 ;
    wire signal_12406 ;
    wire signal_12407 ;
    wire signal_12408 ;
    wire signal_12409 ;
    wire signal_12410 ;
    wire signal_12411 ;
    wire signal_12412 ;
    wire signal_12413 ;
    wire signal_12414 ;
    wire signal_12415 ;
    wire signal_12416 ;
    wire signal_12417 ;
    wire signal_12418 ;
    wire signal_12419 ;
    wire signal_12420 ;
    wire signal_12421 ;
    wire signal_12422 ;
    wire signal_12423 ;
    wire signal_12424 ;
    wire signal_12425 ;
    wire signal_12426 ;
    wire signal_12427 ;
    wire signal_12428 ;
    wire signal_12429 ;
    wire signal_12430 ;
    wire signal_12431 ;
    wire signal_12432 ;
    wire signal_12433 ;
    wire signal_12434 ;
    wire signal_12435 ;
    wire signal_12436 ;
    wire signal_12437 ;
    wire signal_12438 ;
    wire signal_12439 ;
    wire signal_12440 ;
    wire signal_12441 ;
    wire signal_12442 ;
    wire signal_12443 ;
    wire signal_12444 ;
    wire signal_12445 ;
    wire signal_12446 ;
    wire signal_12447 ;
    wire signal_12448 ;
    wire signal_12449 ;
    wire signal_12450 ;
    wire signal_12451 ;
    wire signal_12452 ;
    wire signal_12453 ;
    wire signal_12454 ;
    wire signal_12455 ;
    wire signal_12456 ;
    wire signal_12457 ;
    wire signal_12458 ;
    wire signal_12459 ;
    wire signal_12460 ;
    wire signal_12461 ;
    wire signal_12462 ;
    wire signal_12463 ;
    wire signal_12464 ;
    wire signal_12465 ;
    wire signal_12466 ;
    wire signal_12467 ;
    wire signal_12468 ;
    wire signal_12469 ;
    wire signal_12470 ;
    wire signal_12471 ;
    wire signal_12472 ;
    wire signal_12473 ;
    wire signal_12474 ;
    wire signal_12475 ;
    wire signal_12476 ;
    wire signal_12477 ;
    wire signal_12478 ;
    wire signal_12479 ;
    wire signal_12480 ;
    wire signal_12481 ;
    wire signal_12482 ;
    wire signal_12483 ;
    wire signal_12484 ;
    wire signal_12485 ;
    wire signal_12486 ;
    wire signal_12487 ;
    wire signal_12488 ;
    wire signal_12489 ;
    wire signal_12490 ;
    wire signal_12491 ;
    wire signal_12492 ;
    wire signal_12493 ;
    wire signal_12494 ;
    wire signal_12495 ;
    wire signal_12496 ;
    wire signal_12497 ;
    wire signal_12498 ;
    wire signal_12499 ;
    wire signal_12500 ;
    wire signal_12501 ;
    wire signal_12502 ;
    wire signal_12503 ;
    wire signal_12504 ;
    wire signal_12505 ;
    wire signal_12506 ;
    wire signal_12507 ;
    wire signal_12508 ;
    wire signal_12509 ;
    wire signal_12510 ;
    wire signal_12511 ;
    wire signal_12512 ;
    wire signal_12513 ;
    wire signal_12514 ;
    wire signal_12515 ;
    wire signal_12516 ;
    wire signal_12517 ;
    wire signal_12518 ;
    wire signal_12519 ;
    wire signal_12520 ;
    wire signal_12521 ;
    wire signal_12522 ;
    wire signal_12523 ;
    wire signal_12524 ;
    wire signal_12525 ;
    wire signal_12526 ;
    wire signal_12527 ;
    wire signal_12528 ;
    wire signal_12529 ;
    wire signal_12530 ;
    wire signal_12531 ;
    wire signal_12532 ;
    wire signal_12533 ;
    wire signal_12534 ;
    wire signal_12535 ;
    wire signal_12536 ;
    wire signal_12537 ;
    wire signal_12538 ;
    wire signal_12539 ;
    wire signal_12540 ;
    wire signal_12541 ;
    wire signal_12542 ;
    wire signal_12543 ;
    wire signal_12544 ;
    wire signal_12545 ;
    wire signal_12546 ;
    wire signal_12547 ;
    wire signal_12548 ;
    wire signal_12549 ;
    wire signal_12550 ;
    wire signal_12551 ;
    wire signal_12552 ;
    wire signal_12553 ;
    wire signal_12554 ;
    wire signal_12555 ;
    wire signal_12556 ;
    wire signal_12557 ;
    wire signal_12558 ;
    wire signal_12559 ;
    wire signal_12560 ;
    wire signal_12561 ;
    wire signal_12562 ;
    wire signal_12563 ;
    wire signal_12564 ;
    wire signal_12565 ;
    wire signal_12566 ;
    wire signal_12567 ;
    wire signal_12568 ;
    wire signal_12569 ;
    wire signal_12570 ;
    wire signal_12571 ;
    wire signal_12572 ;
    wire signal_12573 ;
    wire signal_12574 ;
    wire signal_12575 ;
    wire signal_12576 ;
    wire signal_12577 ;
    wire signal_12578 ;
    wire signal_12579 ;
    wire signal_12580 ;
    wire signal_12581 ;
    wire signal_12582 ;
    wire signal_12583 ;
    wire signal_12584 ;
    wire signal_12585 ;
    wire signal_12586 ;
    wire signal_12587 ;
    wire signal_12588 ;
    wire signal_12589 ;
    wire signal_12590 ;
    wire signal_12591 ;
    wire signal_12592 ;
    wire signal_12593 ;
    wire signal_12594 ;
    wire signal_12595 ;
    wire signal_12596 ;
    wire signal_12597 ;
    wire signal_12598 ;
    wire signal_12599 ;
    wire signal_12600 ;
    wire signal_12601 ;
    wire signal_12602 ;
    wire signal_12603 ;
    wire signal_12604 ;
    wire signal_12605 ;
    wire signal_12606 ;
    wire signal_12607 ;
    wire signal_12608 ;
    wire signal_12609 ;
    wire signal_12610 ;
    wire signal_12611 ;
    wire signal_12612 ;
    wire signal_12613 ;
    wire signal_12614 ;
    wire signal_12615 ;
    wire signal_12616 ;
    wire signal_12617 ;
    wire signal_12618 ;
    wire signal_12619 ;
    wire signal_12620 ;
    wire signal_12621 ;
    wire signal_12622 ;
    wire signal_12623 ;
    wire signal_12624 ;
    wire signal_12625 ;
    wire signal_12626 ;
    wire signal_12627 ;
    wire signal_12628 ;
    wire signal_12629 ;
    wire signal_12630 ;
    wire signal_12631 ;
    wire signal_12632 ;
    wire signal_12633 ;
    wire signal_12634 ;
    wire signal_12635 ;
    wire signal_12636 ;
    wire signal_12637 ;
    wire signal_12638 ;
    wire signal_12639 ;
    wire signal_12640 ;
    wire signal_12641 ;
    wire signal_12642 ;
    wire signal_12643 ;
    wire signal_12644 ;
    wire signal_12645 ;
    wire signal_12646 ;
    wire signal_12647 ;
    wire signal_12648 ;
    wire signal_12649 ;
    wire signal_12650 ;
    wire signal_12651 ;
    wire signal_12652 ;
    wire signal_12653 ;
    wire signal_12654 ;
    wire signal_12655 ;
    wire signal_12656 ;
    wire signal_12657 ;
    wire signal_12658 ;
    wire signal_12659 ;
    wire signal_12660 ;
    wire signal_12661 ;
    wire signal_12662 ;
    wire signal_12663 ;
    wire signal_12664 ;
    wire signal_12665 ;
    wire signal_12666 ;
    wire signal_12667 ;
    wire signal_12668 ;
    wire signal_12669 ;
    wire signal_12670 ;
    wire signal_12671 ;
    wire signal_12672 ;
    wire signal_12673 ;
    wire signal_12674 ;
    wire signal_12675 ;
    wire signal_12676 ;
    wire signal_12677 ;
    wire signal_12678 ;
    wire signal_12679 ;
    wire signal_12680 ;
    wire signal_12681 ;
    wire signal_12682 ;
    wire signal_12683 ;
    wire signal_12684 ;
    wire signal_12685 ;
    wire signal_12686 ;
    wire signal_12687 ;
    wire signal_12688 ;
    wire signal_12689 ;
    wire signal_12690 ;
    wire signal_12691 ;
    wire signal_12692 ;
    wire signal_12693 ;
    wire signal_12694 ;
    wire signal_12695 ;
    wire signal_12696 ;
    wire signal_12697 ;
    wire signal_12698 ;
    wire signal_12699 ;
    wire signal_12700 ;
    wire signal_12701 ;
    wire signal_12702 ;
    wire signal_12703 ;
    wire signal_12704 ;
    wire signal_12705 ;
    wire signal_12706 ;
    wire signal_12707 ;
    wire signal_12708 ;
    wire signal_12709 ;
    wire signal_12710 ;
    wire signal_12711 ;
    wire signal_12712 ;
    wire signal_12713 ;
    wire signal_12714 ;
    wire signal_12715 ;
    wire signal_12716 ;
    wire signal_12717 ;
    wire signal_12718 ;
    wire signal_12719 ;
    wire signal_12720 ;
    wire signal_12721 ;
    wire signal_12722 ;
    wire signal_12723 ;
    wire signal_12724 ;
    wire signal_12725 ;
    wire signal_12726 ;
    wire signal_12727 ;
    wire signal_12728 ;
    wire signal_12729 ;
    wire signal_12730 ;
    wire signal_12731 ;
    wire signal_12732 ;
    wire signal_12733 ;
    wire signal_12734 ;
    wire signal_12735 ;
    wire signal_12736 ;
    wire signal_12737 ;
    wire signal_12738 ;
    wire signal_12739 ;
    wire signal_12740 ;
    wire signal_12741 ;
    wire signal_12742 ;
    wire signal_12743 ;
    wire signal_12744 ;
    wire signal_12745 ;
    wire signal_12746 ;
    wire signal_12747 ;
    wire signal_12748 ;
    wire signal_12749 ;
    wire signal_12750 ;
    wire signal_12751 ;
    wire signal_12752 ;
    wire signal_12753 ;
    wire signal_12754 ;
    wire signal_12755 ;
    wire signal_12756 ;
    wire signal_12757 ;
    wire signal_12758 ;
    wire signal_12759 ;
    wire signal_12760 ;
    wire signal_12761 ;
    wire signal_12762 ;
    wire signal_12763 ;
    wire signal_12764 ;
    wire signal_12765 ;
    wire signal_12766 ;
    wire signal_12767 ;
    wire signal_12768 ;
    wire signal_12769 ;
    wire signal_12770 ;
    wire signal_12771 ;
    wire signal_12772 ;
    wire signal_12773 ;
    wire signal_12774 ;
    wire signal_12775 ;
    wire signal_12776 ;
    wire signal_12777 ;
    wire signal_12778 ;
    wire signal_12779 ;
    wire signal_12780 ;
    wire signal_12781 ;
    wire signal_12782 ;
    wire signal_12783 ;
    wire signal_12784 ;
    wire signal_12785 ;
    wire signal_12786 ;
    wire signal_12787 ;
    wire signal_12788 ;
    wire signal_12789 ;
    wire signal_12790 ;
    wire signal_12791 ;
    wire signal_12792 ;
    wire signal_12793 ;
    wire signal_12794 ;
    wire signal_12795 ;
    wire signal_12796 ;
    wire signal_12797 ;
    wire signal_12798 ;
    wire signal_12799 ;
    wire signal_12800 ;
    wire signal_12801 ;
    wire signal_12802 ;
    wire signal_12803 ;
    wire signal_12804 ;
    wire signal_12805 ;
    wire signal_12806 ;
    wire signal_12807 ;
    wire signal_12808 ;
    wire signal_12809 ;
    wire signal_12810 ;
    wire signal_12811 ;
    wire signal_12812 ;
    wire signal_12813 ;
    wire signal_12814 ;
    wire signal_12815 ;
    wire signal_12816 ;
    wire signal_12817 ;
    wire signal_12818 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) cell_927 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2395, signal_2394, signal_942}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_928 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2399, signal_2398, signal_943}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_929 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2403, signal_2402, signal_944}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_930 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2407, signal_2406, signal_945}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_931 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2411, signal_2410, signal_946}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_932 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2415, signal_2414, signal_947}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_933 ( .a ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2419, signal_2418, signal_948}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_934 ( .a ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2423, signal_2422, signal_949}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_949 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .c ({signal_2453, signal_2452, signal_964}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_950 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .c ({signal_2455, signal_2454, signal_965}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_962 ( .a ({signal_2453, signal_2452, signal_964}), .b ({signal_2479, signal_2478, signal_977}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_963 ( .a ({signal_2455, signal_2454, signal_965}), .b ({signal_2481, signal_2480, signal_978}) ) ;

    /* cells in depth 1 */
    buf_clk cell_2385 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( signal_7977 ) ) ;
    buf_clk cell_2387 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( signal_7979 ) ) ;
    buf_clk cell_2389 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( signal_7981 ) ) ;
    buf_clk cell_2391 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_7983 ) ) ;
    buf_clk cell_2393 ( .C ( clk ), .D ( signal_2422 ), .Q ( signal_7985 ) ) ;
    buf_clk cell_2395 ( .C ( clk ), .D ( signal_2423 ), .Q ( signal_7987 ) ) ;
    buf_clk cell_2397 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_7989 ) ) ;
    buf_clk cell_2399 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_7991 ) ) ;
    buf_clk cell_2401 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_7993 ) ) ;
    buf_clk cell_2403 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_7995 ) ) ;
    buf_clk cell_2405 ( .C ( clk ), .D ( signal_2402 ), .Q ( signal_7997 ) ) ;
    buf_clk cell_2407 ( .C ( clk ), .D ( signal_2403 ), .Q ( signal_7999 ) ) ;
    buf_clk cell_2409 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_8001 ) ) ;
    buf_clk cell_2411 ( .C ( clk ), .D ( signal_2394 ), .Q ( signal_8003 ) ) ;
    buf_clk cell_2413 ( .C ( clk ), .D ( signal_2395 ), .Q ( signal_8005 ) ) ;
    buf_clk cell_2415 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_8007 ) ) ;
    buf_clk cell_2417 ( .C ( clk ), .D ( signal_2410 ), .Q ( signal_8009 ) ) ;
    buf_clk cell_2419 ( .C ( clk ), .D ( signal_2411 ), .Q ( signal_8011 ) ) ;
    buf_clk cell_2421 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_8013 ) ) ;
    buf_clk cell_2423 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_8015 ) ) ;
    buf_clk cell_2425 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_8017 ) ) ;
    buf_clk cell_2427 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( signal_8019 ) ) ;
    buf_clk cell_2429 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( signal_8021 ) ) ;
    buf_clk cell_2431 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( signal_8023 ) ) ;
    buf_clk cell_2433 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_8025 ) ) ;
    buf_clk cell_2435 ( .C ( clk ), .D ( signal_2406 ), .Q ( signal_8027 ) ) ;
    buf_clk cell_2437 ( .C ( clk ), .D ( signal_2407 ), .Q ( signal_8029 ) ) ;
    buf_clk cell_2439 ( .C ( clk ), .D ( signal_948 ), .Q ( signal_8031 ) ) ;
    buf_clk cell_2441 ( .C ( clk ), .D ( signal_2418 ), .Q ( signal_8033 ) ) ;
    buf_clk cell_2443 ( .C ( clk ), .D ( signal_2419 ), .Q ( signal_8035 ) ) ;
    buf_clk cell_2445 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( signal_8037 ) ) ;
    buf_clk cell_2447 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( signal_8039 ) ) ;
    buf_clk cell_2449 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( signal_8041 ) ) ;
    buf_clk cell_2451 ( .C ( clk ), .D ( signal_978 ), .Q ( signal_8043 ) ) ;
    buf_clk cell_2453 ( .C ( clk ), .D ( signal_2480 ), .Q ( signal_8045 ) ) ;
    buf_clk cell_2455 ( .C ( clk ), .D ( signal_2481 ), .Q ( signal_8047 ) ) ;
    buf_clk cell_2457 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_8049 ) ) ;
    buf_clk cell_2459 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_8051 ) ) ;
    buf_clk cell_2461 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_8053 ) ) ;
    buf_clk cell_2463 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_8055 ) ) ;
    buf_clk cell_2467 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_8059 ) ) ;
    buf_clk cell_2471 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_8063 ) ) ;
    buf_clk cell_2679 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_8271 ) ) ;
    buf_clk cell_2683 ( .C ( clk ), .D ( signal_2398 ), .Q ( signal_8275 ) ) ;
    buf_clk cell_2687 ( .C ( clk ), .D ( signal_2399 ), .Q ( signal_8279 ) ) ;
    buf_clk cell_2889 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( signal_8481 ) ) ;
    buf_clk cell_2895 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( signal_8487 ) ) ;
    buf_clk cell_2901 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( signal_8493 ) ) ;
    buf_clk cell_3177 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_8769 ) ) ;
    buf_clk cell_3183 ( .C ( clk ), .D ( signal_2414 ), .Q ( signal_8775 ) ) ;
    buf_clk cell_3189 ( .C ( clk ), .D ( signal_2415 ), .Q ( signal_8781 ) ) ;
    buf_clk cell_3399 ( .C ( clk ), .D ( signal_977 ), .Q ( signal_8991 ) ) ;
    buf_clk cell_3407 ( .C ( clk ), .D ( signal_2478 ), .Q ( signal_8999 ) ) ;
    buf_clk cell_3415 ( .C ( clk ), .D ( signal_2479 ), .Q ( signal_9007 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_935 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_2425, signal_2424, signal_950}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_936 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_2427, signal_2426, signal_951}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_937 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_2429, signal_2428, signal_952}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_938 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_2431, signal_2430, signal_953}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_939 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_2433, signal_2432, signal_954}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_940 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_2435, signal_2434, signal_955}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_941 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_2437, signal_2436, signal_956}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_942 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_2439, signal_2438, signal_957}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_943 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_2441, signal_2440, signal_958}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_944 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_2443, signal_2442, signal_959}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_945 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_2445, signal_2444, signal_960}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_946 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_2447, signal_2446, signal_961}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_947 ( .a ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_2449, signal_2448, signal_962}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_948 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_2451, signal_2450, signal_963}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_951 ( .a ({signal_2425, signal_2424, signal_950}), .b ({signal_2457, signal_2456, signal_966}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_952 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2459, signal_2458, signal_967}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_953 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2461, signal_2460, signal_968}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_954 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2463, signal_2462, signal_969}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_955 ( .a ({signal_2433, signal_2432, signal_954}), .b ({signal_2465, signal_2464, signal_970}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_956 ( .a ({signal_2437, signal_2436, signal_956}), .b ({signal_2467, signal_2466, signal_971}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_957 ( .a ({signal_2439, signal_2438, signal_957}), .b ({signal_2469, signal_2468, signal_972}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_958 ( .a ({signal_2443, signal_2442, signal_959}), .b ({signal_2471, signal_2470, signal_973}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_959 ( .a ({signal_2445, signal_2444, signal_960}), .b ({signal_2473, signal_2472, signal_974}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_960 ( .a ({signal_2447, signal_2446, signal_961}), .b ({signal_2475, signal_2474, signal_975}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_961 ( .a ({signal_2449, signal_2448, signal_962}), .b ({signal_2477, signal_2476, signal_976}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_964 ( .a ({signal_2399, signal_2398, signal_943}), .b ({signal_2403, signal_2402, signal_944}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_2483, signal_2482, signal_979}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_965 ( .a ({signal_2419, signal_2418, signal_948}), .b ({signal_2423, signal_2422, signal_949}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_2485, signal_2484, signal_980}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_966 ( .a ({signal_2407, signal_2406, signal_945}), .b ({signal_2411, signal_2410, signal_946}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_2487, signal_2486, signal_981}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_967 ( .a ({signal_2403, signal_2402, signal_944}), .b ({signal_2411, signal_2410, signal_946}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_2489, signal_2488, signal_982}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_968 ( .a ({signal_2403, signal_2402, signal_944}), .b ({signal_2407, signal_2406, signal_945}), .clk ( clk ), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_2491, signal_2490, signal_983}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_969 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2399, signal_2398, signal_943}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_2493, signal_2492, signal_984}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_970 ( .a ({signal_2395, signal_2394, signal_942}), .b ({SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_2495, signal_2494, signal_985}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_971 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2411, signal_2410, signal_946}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_2497, signal_2496, signal_986}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_972 ( .a ({signal_2415, signal_2414, signal_947}), .b ({signal_2423, signal_2422, signal_949}), .clk ( clk ), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_2499, signal_2498, signal_987}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_973 ( .a ({signal_2415, signal_2414, signal_947}), .b ({signal_2419, signal_2418, signal_948}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_2501, signal_2500, signal_988}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_974 ( .a ({signal_2415, signal_2414, signal_947}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_2503, signal_2502, signal_989}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_975 ( .a ({signal_2399, signal_2398, signal_943}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_2505, signal_2504, signal_990}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_976 ( .a ({signal_2407, signal_2406, signal_945}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_2507, signal_2506, signal_991}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_977 ( .a ({signal_2419, signal_2418, signal_948}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_2509, signal_2508, signal_992}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_978 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2403, signal_2402, signal_944}), .clk ( clk ), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_2511, signal_2510, signal_993}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_979 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2411, signal_2410, signal_946}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_2513, signal_2512, signal_994}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_980 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2403, signal_2402, signal_944}), .clk ( clk ), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_2515, signal_2514, signal_995}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_981 ( .a ({signal_2403, signal_2402, signal_944}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_2517, signal_2516, signal_996}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_982 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2415, signal_2414, signal_947}), .clk ( clk ), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_2519, signal_2518, signal_997}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_983 ( .a ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2423, signal_2422, signal_949}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_2521, signal_2520, signal_998}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_984 ( .a ({signal_2395, signal_2394, signal_942}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_2523, signal_2522, signal_999}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_985 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2419, signal_2418, signal_948}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({signal_2525, signal_2524, signal_1000}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_986 ( .a ({signal_2395, signal_2394, signal_942}), .b ({signal_2399, signal_2398, signal_943}), .clk ( clk ), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_2527, signal_2526, signal_1001}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_987 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2407, signal_2406, signal_945}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({signal_2529, signal_2528, signal_1002}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_989 ( .a ({signal_2411, signal_2410, signal_946}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_2533, signal_2532, signal_1004}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_990 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2407, signal_2406, signal_945}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({signal_2535, signal_2534, signal_1005}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_991 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2415, signal_2414, signal_947}), .clk ( clk ), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_2537, signal_2536, signal_1006}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_992 ( .a ({signal_2403, signal_2402, signal_944}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({signal_2539, signal_2538, signal_1007}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_993 ( .a ({signal_2415, signal_2414, signal_947}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_2541, signal_2540, signal_1008}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_994 ( .a ({signal_2411, signal_2410, signal_946}), .b ({signal_2415, signal_2414, signal_947}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({signal_2543, signal_2542, signal_1009}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_995 ( .a ({signal_2395, signal_2394, signal_942}), .b ({signal_2403, signal_2402, signal_944}), .clk ( clk ), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_2545, signal_2544, signal_1010}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_996 ( .a ({signal_2403, signal_2402, signal_944}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({signal_2547, signal_2546, signal_1011}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_997 ( .a ({signal_2407, signal_2406, signal_945}), .b ({signal_2415, signal_2414, signal_947}), .clk ( clk ), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_2549, signal_2548, signal_1012}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_998 ( .a ({signal_2407, signal_2406, signal_945}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({signal_2551, signal_2550, signal_1013}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1000 ( .a ({signal_2407, signal_2406, signal_945}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_2555, signal_2554, signal_1015}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1001 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2419, signal_2418, signal_948}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({signal_2557, signal_2556, signal_1016}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1002 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2411, signal_2410, signal_946}), .clk ( clk ), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_2559, signal_2558, signal_1017}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1003 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2423, signal_2422, signal_949}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({signal_2561, signal_2560, signal_1018}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1016 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_2587, signal_2586, signal_1031}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1017 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2589, signal_2588, signal_1032}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1018 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2591, signal_2590, signal_1033}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1019 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2593, signal_2592, signal_1034}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1020 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2595, signal_2594, signal_1035}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1021 ( .a ({signal_2499, signal_2498, signal_987}), .b ({signal_2597, signal_2596, signal_1036}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1022 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2599, signal_2598, signal_1037}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1023 ( .a ({signal_2503, signal_2502, signal_989}), .b ({signal_2601, signal_2600, signal_1038}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1024 ( .a ({signal_2505, signal_2504, signal_990}), .b ({signal_2603, signal_2602, signal_1039}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1025 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2605, signal_2604, signal_1040}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1026 ( .a ({signal_2509, signal_2508, signal_992}), .b ({signal_2607, signal_2606, signal_1041}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1027 ( .a ({signal_2511, signal_2510, signal_993}), .b ({signal_2609, signal_2608, signal_1042}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1028 ( .a ({signal_2515, signal_2514, signal_995}), .b ({signal_2611, signal_2610, signal_1043}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1029 ( .a ({signal_2517, signal_2516, signal_996}), .b ({signal_2613, signal_2612, signal_1044}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1030 ( .a ({signal_2519, signal_2518, signal_997}), .b ({signal_2615, signal_2614, signal_1045}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1031 ( .a ({signal_2521, signal_2520, signal_998}), .b ({signal_2617, signal_2616, signal_1046}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1032 ( .a ({signal_2525, signal_2524, signal_1000}), .b ({signal_2619, signal_2618, signal_1047}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1034 ( .a ({signal_2533, signal_2532, signal_1004}), .b ({signal_2623, signal_2622, signal_1049}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1035 ( .a ({signal_2535, signal_2534, signal_1005}), .b ({signal_2625, signal_2624, signal_1050}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1036 ( .a ({signal_2537, signal_2536, signal_1006}), .b ({signal_2627, signal_2626, signal_1051}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1037 ( .a ({signal_2541, signal_2540, signal_1008}), .b ({signal_2629, signal_2628, signal_1052}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1038 ( .a ({signal_2543, signal_2542, signal_1009}), .b ({signal_2631, signal_2630, signal_1053}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1039 ( .a ({signal_2551, signal_2550, signal_1013}), .b ({signal_2633, signal_2632, signal_1054}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1041 ( .a ({signal_2555, signal_2554, signal_1015}), .b ({signal_2637, signal_2636, signal_1056}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1042 ( .a ({signal_2557, signal_2556, signal_1016}), .b ({signal_2639, signal_2638, signal_1057}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1043 ( .a ({signal_2559, signal_2558, signal_1017}), .b ({signal_2641, signal_2640, signal_1058}) ) ;
    buf_clk cell_2386 ( .C ( clk ), .D ( signal_7977 ), .Q ( signal_7978 ) ) ;
    buf_clk cell_2388 ( .C ( clk ), .D ( signal_7979 ), .Q ( signal_7980 ) ) ;
    buf_clk cell_2390 ( .C ( clk ), .D ( signal_7981 ), .Q ( signal_7982 ) ) ;
    buf_clk cell_2392 ( .C ( clk ), .D ( signal_7983 ), .Q ( signal_7984 ) ) ;
    buf_clk cell_2394 ( .C ( clk ), .D ( signal_7985 ), .Q ( signal_7986 ) ) ;
    buf_clk cell_2396 ( .C ( clk ), .D ( signal_7987 ), .Q ( signal_7988 ) ) ;
    buf_clk cell_2398 ( .C ( clk ), .D ( signal_7989 ), .Q ( signal_7990 ) ) ;
    buf_clk cell_2400 ( .C ( clk ), .D ( signal_7991 ), .Q ( signal_7992 ) ) ;
    buf_clk cell_2402 ( .C ( clk ), .D ( signal_7993 ), .Q ( signal_7994 ) ) ;
    buf_clk cell_2404 ( .C ( clk ), .D ( signal_7995 ), .Q ( signal_7996 ) ) ;
    buf_clk cell_2406 ( .C ( clk ), .D ( signal_7997 ), .Q ( signal_7998 ) ) ;
    buf_clk cell_2408 ( .C ( clk ), .D ( signal_7999 ), .Q ( signal_8000 ) ) ;
    buf_clk cell_2410 ( .C ( clk ), .D ( signal_8001 ), .Q ( signal_8002 ) ) ;
    buf_clk cell_2412 ( .C ( clk ), .D ( signal_8003 ), .Q ( signal_8004 ) ) ;
    buf_clk cell_2414 ( .C ( clk ), .D ( signal_8005 ), .Q ( signal_8006 ) ) ;
    buf_clk cell_2416 ( .C ( clk ), .D ( signal_8007 ), .Q ( signal_8008 ) ) ;
    buf_clk cell_2418 ( .C ( clk ), .D ( signal_8009 ), .Q ( signal_8010 ) ) ;
    buf_clk cell_2420 ( .C ( clk ), .D ( signal_8011 ), .Q ( signal_8012 ) ) ;
    buf_clk cell_2422 ( .C ( clk ), .D ( signal_8013 ), .Q ( signal_8014 ) ) ;
    buf_clk cell_2424 ( .C ( clk ), .D ( signal_8015 ), .Q ( signal_8016 ) ) ;
    buf_clk cell_2426 ( .C ( clk ), .D ( signal_8017 ), .Q ( signal_8018 ) ) ;
    buf_clk cell_2428 ( .C ( clk ), .D ( signal_8019 ), .Q ( signal_8020 ) ) ;
    buf_clk cell_2430 ( .C ( clk ), .D ( signal_8021 ), .Q ( signal_8022 ) ) ;
    buf_clk cell_2432 ( .C ( clk ), .D ( signal_8023 ), .Q ( signal_8024 ) ) ;
    buf_clk cell_2434 ( .C ( clk ), .D ( signal_8025 ), .Q ( signal_8026 ) ) ;
    buf_clk cell_2436 ( .C ( clk ), .D ( signal_8027 ), .Q ( signal_8028 ) ) ;
    buf_clk cell_2438 ( .C ( clk ), .D ( signal_8029 ), .Q ( signal_8030 ) ) ;
    buf_clk cell_2440 ( .C ( clk ), .D ( signal_8031 ), .Q ( signal_8032 ) ) ;
    buf_clk cell_2442 ( .C ( clk ), .D ( signal_8033 ), .Q ( signal_8034 ) ) ;
    buf_clk cell_2444 ( .C ( clk ), .D ( signal_8035 ), .Q ( signal_8036 ) ) ;
    buf_clk cell_2446 ( .C ( clk ), .D ( signal_8037 ), .Q ( signal_8038 ) ) ;
    buf_clk cell_2448 ( .C ( clk ), .D ( signal_8039 ), .Q ( signal_8040 ) ) ;
    buf_clk cell_2450 ( .C ( clk ), .D ( signal_8041 ), .Q ( signal_8042 ) ) ;
    buf_clk cell_2452 ( .C ( clk ), .D ( signal_8043 ), .Q ( signal_8044 ) ) ;
    buf_clk cell_2454 ( .C ( clk ), .D ( signal_8045 ), .Q ( signal_8046 ) ) ;
    buf_clk cell_2456 ( .C ( clk ), .D ( signal_8047 ), .Q ( signal_8048 ) ) ;
    buf_clk cell_2458 ( .C ( clk ), .D ( signal_8049 ), .Q ( signal_8050 ) ) ;
    buf_clk cell_2460 ( .C ( clk ), .D ( signal_8051 ), .Q ( signal_8052 ) ) ;
    buf_clk cell_2462 ( .C ( clk ), .D ( signal_8053 ), .Q ( signal_8054 ) ) ;
    buf_clk cell_2464 ( .C ( clk ), .D ( signal_8055 ), .Q ( signal_8056 ) ) ;
    buf_clk cell_2468 ( .C ( clk ), .D ( signal_8059 ), .Q ( signal_8060 ) ) ;
    buf_clk cell_2472 ( .C ( clk ), .D ( signal_8063 ), .Q ( signal_8064 ) ) ;
    buf_clk cell_2680 ( .C ( clk ), .D ( signal_8271 ), .Q ( signal_8272 ) ) ;
    buf_clk cell_2684 ( .C ( clk ), .D ( signal_8275 ), .Q ( signal_8276 ) ) ;
    buf_clk cell_2688 ( .C ( clk ), .D ( signal_8279 ), .Q ( signal_8280 ) ) ;
    buf_clk cell_2890 ( .C ( clk ), .D ( signal_8481 ), .Q ( signal_8482 ) ) ;
    buf_clk cell_2896 ( .C ( clk ), .D ( signal_8487 ), .Q ( signal_8488 ) ) ;
    buf_clk cell_2902 ( .C ( clk ), .D ( signal_8493 ), .Q ( signal_8494 ) ) ;
    buf_clk cell_3178 ( .C ( clk ), .D ( signal_8769 ), .Q ( signal_8770 ) ) ;
    buf_clk cell_3184 ( .C ( clk ), .D ( signal_8775 ), .Q ( signal_8776 ) ) ;
    buf_clk cell_3190 ( .C ( clk ), .D ( signal_8781 ), .Q ( signal_8782 ) ) ;
    buf_clk cell_3400 ( .C ( clk ), .D ( signal_8991 ), .Q ( signal_8992 ) ) ;
    buf_clk cell_3408 ( .C ( clk ), .D ( signal_8999 ), .Q ( signal_9000 ) ) ;
    buf_clk cell_3416 ( .C ( clk ), .D ( signal_9007 ), .Q ( signal_9008 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_2465 ( .C ( clk ), .D ( signal_8056 ), .Q ( signal_8057 ) ) ;
    buf_clk cell_2469 ( .C ( clk ), .D ( signal_8060 ), .Q ( signal_8061 ) ) ;
    buf_clk cell_2473 ( .C ( clk ), .D ( signal_8064 ), .Q ( signal_8065 ) ) ;
    buf_clk cell_2475 ( .C ( clk ), .D ( signal_8026 ), .Q ( signal_8067 ) ) ;
    buf_clk cell_2477 ( .C ( clk ), .D ( signal_8028 ), .Q ( signal_8069 ) ) ;
    buf_clk cell_2479 ( .C ( clk ), .D ( signal_8030 ), .Q ( signal_8071 ) ) ;
    buf_clk cell_2481 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_8073 ) ) ;
    buf_clk cell_2483 ( .C ( clk ), .D ( signal_2514 ), .Q ( signal_8075 ) ) ;
    buf_clk cell_2485 ( .C ( clk ), .D ( signal_2515 ), .Q ( signal_8077 ) ) ;
    buf_clk cell_2487 ( .C ( clk ), .D ( signal_1010 ), .Q ( signal_8079 ) ) ;
    buf_clk cell_2489 ( .C ( clk ), .D ( signal_2544 ), .Q ( signal_8081 ) ) ;
    buf_clk cell_2491 ( .C ( clk ), .D ( signal_2545 ), .Q ( signal_8083 ) ) ;
    buf_clk cell_2493 ( .C ( clk ), .D ( signal_992 ), .Q ( signal_8085 ) ) ;
    buf_clk cell_2495 ( .C ( clk ), .D ( signal_2508 ), .Q ( signal_8087 ) ) ;
    buf_clk cell_2497 ( .C ( clk ), .D ( signal_2509 ), .Q ( signal_8089 ) ) ;
    buf_clk cell_2499 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_8091 ) ) ;
    buf_clk cell_2501 ( .C ( clk ), .D ( signal_2510 ), .Q ( signal_8093 ) ) ;
    buf_clk cell_2503 ( .C ( clk ), .D ( signal_2511 ), .Q ( signal_8095 ) ) ;
    buf_clk cell_2505 ( .C ( clk ), .D ( signal_1008 ), .Q ( signal_8097 ) ) ;
    buf_clk cell_2507 ( .C ( clk ), .D ( signal_2540 ), .Q ( signal_8099 ) ) ;
    buf_clk cell_2509 ( .C ( clk ), .D ( signal_2541 ), .Q ( signal_8101 ) ) ;
    buf_clk cell_2511 ( .C ( clk ), .D ( signal_991 ), .Q ( signal_8103 ) ) ;
    buf_clk cell_2513 ( .C ( clk ), .D ( signal_2506 ), .Q ( signal_8105 ) ) ;
    buf_clk cell_2515 ( .C ( clk ), .D ( signal_2507 ), .Q ( signal_8107 ) ) ;
    buf_clk cell_2517 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_8109 ) ) ;
    buf_clk cell_2519 ( .C ( clk ), .D ( signal_2442 ), .Q ( signal_8111 ) ) ;
    buf_clk cell_2521 ( .C ( clk ), .D ( signal_2443 ), .Q ( signal_8113 ) ) ;
    buf_clk cell_2523 ( .C ( clk ), .D ( signal_987 ), .Q ( signal_8115 ) ) ;
    buf_clk cell_2525 ( .C ( clk ), .D ( signal_2498 ), .Q ( signal_8117 ) ) ;
    buf_clk cell_2527 ( .C ( clk ), .D ( signal_2499 ), .Q ( signal_8119 ) ) ;
    buf_clk cell_2529 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_8121 ) ) ;
    buf_clk cell_2531 ( .C ( clk ), .D ( signal_2446 ), .Q ( signal_8123 ) ) ;
    buf_clk cell_2533 ( .C ( clk ), .D ( signal_2447 ), .Q ( signal_8125 ) ) ;
    buf_clk cell_2535 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_8127 ) ) ;
    buf_clk cell_2537 ( .C ( clk ), .D ( signal_2482 ), .Q ( signal_8129 ) ) ;
    buf_clk cell_2539 ( .C ( clk ), .D ( signal_2483 ), .Q ( signal_8131 ) ) ;
    buf_clk cell_2541 ( .C ( clk ), .D ( signal_8014 ), .Q ( signal_8133 ) ) ;
    buf_clk cell_2543 ( .C ( clk ), .D ( signal_8016 ), .Q ( signal_8135 ) ) ;
    buf_clk cell_2545 ( .C ( clk ), .D ( signal_8018 ), .Q ( signal_8137 ) ) ;
    buf_clk cell_2547 ( .C ( clk ), .D ( signal_960 ), .Q ( signal_8139 ) ) ;
    buf_clk cell_2549 ( .C ( clk ), .D ( signal_2444 ), .Q ( signal_8141 ) ) ;
    buf_clk cell_2551 ( .C ( clk ), .D ( signal_2445 ), .Q ( signal_8143 ) ) ;
    buf_clk cell_2553 ( .C ( clk ), .D ( signal_8050 ), .Q ( signal_8145 ) ) ;
    buf_clk cell_2555 ( .C ( clk ), .D ( signal_8052 ), .Q ( signal_8147 ) ) ;
    buf_clk cell_2557 ( .C ( clk ), .D ( signal_8054 ), .Q ( signal_8149 ) ) ;
    buf_clk cell_2559 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_8151 ) ) ;
    buf_clk cell_2561 ( .C ( clk ), .D ( signal_2424 ), .Q ( signal_8153 ) ) ;
    buf_clk cell_2563 ( .C ( clk ), .D ( signal_2425 ), .Q ( signal_8155 ) ) ;
    buf_clk cell_2565 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_8157 ) ) ;
    buf_clk cell_2567 ( .C ( clk ), .D ( signal_2524 ), .Q ( signal_8159 ) ) ;
    buf_clk cell_2569 ( .C ( clk ), .D ( signal_2525 ), .Q ( signal_8161 ) ) ;
    buf_clk cell_2571 ( .C ( clk ), .D ( signal_7984 ), .Q ( signal_8163 ) ) ;
    buf_clk cell_2573 ( .C ( clk ), .D ( signal_7986 ), .Q ( signal_8165 ) ) ;
    buf_clk cell_2575 ( .C ( clk ), .D ( signal_7988 ), .Q ( signal_8167 ) ) ;
    buf_clk cell_2577 ( .C ( clk ), .D ( signal_8008 ), .Q ( signal_8169 ) ) ;
    buf_clk cell_2579 ( .C ( clk ), .D ( signal_8010 ), .Q ( signal_8171 ) ) ;
    buf_clk cell_2581 ( .C ( clk ), .D ( signal_8012 ), .Q ( signal_8173 ) ) ;
    buf_clk cell_2583 ( .C ( clk ), .D ( signal_989 ), .Q ( signal_8175 ) ) ;
    buf_clk cell_2585 ( .C ( clk ), .D ( signal_2502 ), .Q ( signal_8177 ) ) ;
    buf_clk cell_2587 ( .C ( clk ), .D ( signal_2503 ), .Q ( signal_8179 ) ) ;
    buf_clk cell_2589 ( .C ( clk ), .D ( signal_8032 ), .Q ( signal_8181 ) ) ;
    buf_clk cell_2591 ( .C ( clk ), .D ( signal_8034 ), .Q ( signal_8183 ) ) ;
    buf_clk cell_2593 ( .C ( clk ), .D ( signal_8036 ), .Q ( signal_8185 ) ) ;
    buf_clk cell_2595 ( .C ( clk ), .D ( signal_986 ), .Q ( signal_8187 ) ) ;
    buf_clk cell_2597 ( .C ( clk ), .D ( signal_2496 ), .Q ( signal_8189 ) ) ;
    buf_clk cell_2599 ( .C ( clk ), .D ( signal_2497 ), .Q ( signal_8191 ) ) ;
    buf_clk cell_2601 ( .C ( clk ), .D ( signal_1032 ), .Q ( signal_8193 ) ) ;
    buf_clk cell_2603 ( .C ( clk ), .D ( signal_2588 ), .Q ( signal_8195 ) ) ;
    buf_clk cell_2605 ( .C ( clk ), .D ( signal_2589 ), .Q ( signal_8197 ) ) ;
    buf_clk cell_2607 ( .C ( clk ), .D ( signal_1016 ), .Q ( signal_8199 ) ) ;
    buf_clk cell_2609 ( .C ( clk ), .D ( signal_2556 ), .Q ( signal_8201 ) ) ;
    buf_clk cell_2611 ( .C ( clk ), .D ( signal_2557 ), .Q ( signal_8203 ) ) ;
    buf_clk cell_2613 ( .C ( clk ), .D ( signal_8020 ), .Q ( signal_8205 ) ) ;
    buf_clk cell_2615 ( .C ( clk ), .D ( signal_8022 ), .Q ( signal_8207 ) ) ;
    buf_clk cell_2617 ( .C ( clk ), .D ( signal_8024 ), .Q ( signal_8209 ) ) ;
    buf_clk cell_2619 ( .C ( clk ), .D ( signal_8038 ), .Q ( signal_8211 ) ) ;
    buf_clk cell_2621 ( .C ( clk ), .D ( signal_8040 ), .Q ( signal_8213 ) ) ;
    buf_clk cell_2623 ( .C ( clk ), .D ( signal_8042 ), .Q ( signal_8215 ) ) ;
    buf_clk cell_2625 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_8217 ) ) ;
    buf_clk cell_2627 ( .C ( clk ), .D ( signal_2448 ), .Q ( signal_8219 ) ) ;
    buf_clk cell_2629 ( .C ( clk ), .D ( signal_2449 ), .Q ( signal_8221 ) ) ;
    buf_clk cell_2631 ( .C ( clk ), .D ( signal_998 ), .Q ( signal_8223 ) ) ;
    buf_clk cell_2633 ( .C ( clk ), .D ( signal_2520 ), .Q ( signal_8225 ) ) ;
    buf_clk cell_2635 ( .C ( clk ), .D ( signal_2521 ), .Q ( signal_8227 ) ) ;
    buf_clk cell_2637 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_8229 ) ) ;
    buf_clk cell_2639 ( .C ( clk ), .D ( signal_2526 ), .Q ( signal_8231 ) ) ;
    buf_clk cell_2641 ( .C ( clk ), .D ( signal_2527 ), .Q ( signal_8233 ) ) ;
    buf_clk cell_2643 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_8235 ) ) ;
    buf_clk cell_2645 ( .C ( clk ), .D ( signal_2542 ), .Q ( signal_8237 ) ) ;
    buf_clk cell_2647 ( .C ( clk ), .D ( signal_2543 ), .Q ( signal_8239 ) ) ;
    buf_clk cell_2649 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_8241 ) ) ;
    buf_clk cell_2651 ( .C ( clk ), .D ( signal_2430 ), .Q ( signal_8243 ) ) ;
    buf_clk cell_2653 ( .C ( clk ), .D ( signal_2431 ), .Q ( signal_8245 ) ) ;
    buf_clk cell_2655 ( .C ( clk ), .D ( signal_988 ), .Q ( signal_8247 ) ) ;
    buf_clk cell_2657 ( .C ( clk ), .D ( signal_2500 ), .Q ( signal_8249 ) ) ;
    buf_clk cell_2659 ( .C ( clk ), .D ( signal_2501 ), .Q ( signal_8251 ) ) ;
    buf_clk cell_2661 ( .C ( clk ), .D ( signal_7990 ), .Q ( signal_8253 ) ) ;
    buf_clk cell_2663 ( .C ( clk ), .D ( signal_7992 ), .Q ( signal_8255 ) ) ;
    buf_clk cell_2665 ( .C ( clk ), .D ( signal_7994 ), .Q ( signal_8257 ) ) ;
    buf_clk cell_2667 ( .C ( clk ), .D ( signal_1004 ), .Q ( signal_8259 ) ) ;
    buf_clk cell_2669 ( .C ( clk ), .D ( signal_2532 ), .Q ( signal_8261 ) ) ;
    buf_clk cell_2671 ( .C ( clk ), .D ( signal_2533 ), .Q ( signal_8263 ) ) ;
    buf_clk cell_2673 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_8265 ) ) ;
    buf_clk cell_2675 ( .C ( clk ), .D ( signal_2438 ), .Q ( signal_8267 ) ) ;
    buf_clk cell_2677 ( .C ( clk ), .D ( signal_2439 ), .Q ( signal_8269 ) ) ;
    buf_clk cell_2681 ( .C ( clk ), .D ( signal_8272 ), .Q ( signal_8273 ) ) ;
    buf_clk cell_2685 ( .C ( clk ), .D ( signal_8276 ), .Q ( signal_8277 ) ) ;
    buf_clk cell_2689 ( .C ( clk ), .D ( signal_8280 ), .Q ( signal_8281 ) ) ;
    buf_clk cell_2691 ( .C ( clk ), .D ( signal_984 ), .Q ( signal_8283 ) ) ;
    buf_clk cell_2693 ( .C ( clk ), .D ( signal_2492 ), .Q ( signal_8285 ) ) ;
    buf_clk cell_2695 ( .C ( clk ), .D ( signal_2493 ), .Q ( signal_8287 ) ) ;
    buf_clk cell_2697 ( .C ( clk ), .D ( signal_997 ), .Q ( signal_8289 ) ) ;
    buf_clk cell_2699 ( .C ( clk ), .D ( signal_2518 ), .Q ( signal_8291 ) ) ;
    buf_clk cell_2701 ( .C ( clk ), .D ( signal_2519 ), .Q ( signal_8293 ) ) ;
    buf_clk cell_2703 ( .C ( clk ), .D ( signal_1007 ), .Q ( signal_8295 ) ) ;
    buf_clk cell_2705 ( .C ( clk ), .D ( signal_2538 ), .Q ( signal_8297 ) ) ;
    buf_clk cell_2707 ( .C ( clk ), .D ( signal_2539 ), .Q ( signal_8299 ) ) ;
    buf_clk cell_2709 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_8301 ) ) ;
    buf_clk cell_2711 ( .C ( clk ), .D ( signal_2426 ), .Q ( signal_8303 ) ) ;
    buf_clk cell_2713 ( .C ( clk ), .D ( signal_2427 ), .Q ( signal_8305 ) ) ;
    buf_clk cell_2715 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_8307 ) ) ;
    buf_clk cell_2717 ( .C ( clk ), .D ( signal_2486 ), .Q ( signal_8309 ) ) ;
    buf_clk cell_2719 ( .C ( clk ), .D ( signal_2487 ), .Q ( signal_8311 ) ) ;
    buf_clk cell_2721 ( .C ( clk ), .D ( signal_7978 ), .Q ( signal_8313 ) ) ;
    buf_clk cell_2723 ( .C ( clk ), .D ( signal_7980 ), .Q ( signal_8315 ) ) ;
    buf_clk cell_2725 ( .C ( clk ), .D ( signal_7982 ), .Q ( signal_8317 ) ) ;
    buf_clk cell_2727 ( .C ( clk ), .D ( signal_990 ), .Q ( signal_8319 ) ) ;
    buf_clk cell_2729 ( .C ( clk ), .D ( signal_2504 ), .Q ( signal_8321 ) ) ;
    buf_clk cell_2731 ( .C ( clk ), .D ( signal_2505 ), .Q ( signal_8323 ) ) ;
    buf_clk cell_2733 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_8325 ) ) ;
    buf_clk cell_2735 ( .C ( clk ), .D ( signal_2536 ), .Q ( signal_8327 ) ) ;
    buf_clk cell_2737 ( .C ( clk ), .D ( signal_2537 ), .Q ( signal_8329 ) ) ;
    buf_clk cell_2739 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_8331 ) ) ;
    buf_clk cell_2741 ( .C ( clk ), .D ( signal_2490 ), .Q ( signal_8333 ) ) ;
    buf_clk cell_2743 ( .C ( clk ), .D ( signal_2491 ), .Q ( signal_8335 ) ) ;
    buf_clk cell_2745 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_8337 ) ) ;
    buf_clk cell_2747 ( .C ( clk ), .D ( signal_2484 ), .Q ( signal_8339 ) ) ;
    buf_clk cell_2749 ( .C ( clk ), .D ( signal_2485 ), .Q ( signal_8341 ) ) ;
    buf_clk cell_2751 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_8343 ) ) ;
    buf_clk cell_2753 ( .C ( clk ), .D ( signal_2522 ), .Q ( signal_8345 ) ) ;
    buf_clk cell_2755 ( .C ( clk ), .D ( signal_2523 ), .Q ( signal_8347 ) ) ;
    buf_clk cell_2757 ( .C ( clk ), .D ( signal_972 ), .Q ( signal_8349 ) ) ;
    buf_clk cell_2759 ( .C ( clk ), .D ( signal_2468 ), .Q ( signal_8351 ) ) ;
    buf_clk cell_2761 ( .C ( clk ), .D ( signal_2469 ), .Q ( signal_8353 ) ) ;
    buf_clk cell_2763 ( .C ( clk ), .D ( signal_976 ), .Q ( signal_8355 ) ) ;
    buf_clk cell_2765 ( .C ( clk ), .D ( signal_2476 ), .Q ( signal_8357 ) ) ;
    buf_clk cell_2767 ( .C ( clk ), .D ( signal_2477 ), .Q ( signal_8359 ) ) ;
    buf_clk cell_2769 ( .C ( clk ), .D ( signal_1057 ), .Q ( signal_8361 ) ) ;
    buf_clk cell_2771 ( .C ( clk ), .D ( signal_2638 ), .Q ( signal_8363 ) ) ;
    buf_clk cell_2773 ( .C ( clk ), .D ( signal_2639 ), .Q ( signal_8365 ) ) ;
    buf_clk cell_2775 ( .C ( clk ), .D ( signal_1039 ), .Q ( signal_8367 ) ) ;
    buf_clk cell_2777 ( .C ( clk ), .D ( signal_2602 ), .Q ( signal_8369 ) ) ;
    buf_clk cell_2779 ( .C ( clk ), .D ( signal_2603 ), .Q ( signal_8371 ) ) ;
    buf_clk cell_2781 ( .C ( clk ), .D ( signal_1046 ), .Q ( signal_8373 ) ) ;
    buf_clk cell_2783 ( .C ( clk ), .D ( signal_2616 ), .Q ( signal_8375 ) ) ;
    buf_clk cell_2785 ( .C ( clk ), .D ( signal_2617 ), .Q ( signal_8377 ) ) ;
    buf_clk cell_2787 ( .C ( clk ), .D ( signal_1005 ), .Q ( signal_8379 ) ) ;
    buf_clk cell_2789 ( .C ( clk ), .D ( signal_2534 ), .Q ( signal_8381 ) ) ;
    buf_clk cell_2791 ( .C ( clk ), .D ( signal_2535 ), .Q ( signal_8383 ) ) ;
    buf_clk cell_2793 ( .C ( clk ), .D ( signal_1041 ), .Q ( signal_8385 ) ) ;
    buf_clk cell_2795 ( .C ( clk ), .D ( signal_2606 ), .Q ( signal_8387 ) ) ;
    buf_clk cell_2797 ( .C ( clk ), .D ( signal_2607 ), .Q ( signal_8389 ) ) ;
    buf_clk cell_2799 ( .C ( clk ), .D ( signal_1034 ), .Q ( signal_8391 ) ) ;
    buf_clk cell_2801 ( .C ( clk ), .D ( signal_2592 ), .Q ( signal_8393 ) ) ;
    buf_clk cell_2803 ( .C ( clk ), .D ( signal_2593 ), .Q ( signal_8395 ) ) ;
    buf_clk cell_2805 ( .C ( clk ), .D ( signal_996 ), .Q ( signal_8397 ) ) ;
    buf_clk cell_2807 ( .C ( clk ), .D ( signal_2516 ), .Q ( signal_8399 ) ) ;
    buf_clk cell_2809 ( .C ( clk ), .D ( signal_2517 ), .Q ( signal_8401 ) ) ;
    buf_clk cell_2811 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_8403 ) ) ;
    buf_clk cell_2813 ( .C ( clk ), .D ( signal_2512 ), .Q ( signal_8405 ) ) ;
    buf_clk cell_2815 ( .C ( clk ), .D ( signal_2513 ), .Q ( signal_8407 ) ) ;
    buf_clk cell_2817 ( .C ( clk ), .D ( signal_985 ), .Q ( signal_8409 ) ) ;
    buf_clk cell_2819 ( .C ( clk ), .D ( signal_2494 ), .Q ( signal_8411 ) ) ;
    buf_clk cell_2821 ( .C ( clk ), .D ( signal_2495 ), .Q ( signal_8413 ) ) ;
    buf_clk cell_2891 ( .C ( clk ), .D ( signal_8482 ), .Q ( signal_8483 ) ) ;
    buf_clk cell_2897 ( .C ( clk ), .D ( signal_8488 ), .Q ( signal_8489 ) ) ;
    buf_clk cell_2903 ( .C ( clk ), .D ( signal_8494 ), .Q ( signal_8495 ) ) ;
    buf_clk cell_3027 ( .C ( clk ), .D ( signal_1054 ), .Q ( signal_8619 ) ) ;
    buf_clk cell_3031 ( .C ( clk ), .D ( signal_2632 ), .Q ( signal_8623 ) ) ;
    buf_clk cell_3035 ( .C ( clk ), .D ( signal_2633 ), .Q ( signal_8627 ) ) ;
    buf_clk cell_3051 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_8643 ) ) ;
    buf_clk cell_3055 ( .C ( clk ), .D ( signal_2428 ), .Q ( signal_8647 ) ) ;
    buf_clk cell_3059 ( .C ( clk ), .D ( signal_2429 ), .Q ( signal_8651 ) ) ;
    buf_clk cell_3129 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_8721 ) ) ;
    buf_clk cell_3133 ( .C ( clk ), .D ( signal_2440 ), .Q ( signal_8725 ) ) ;
    buf_clk cell_3137 ( .C ( clk ), .D ( signal_2441 ), .Q ( signal_8729 ) ) ;
    buf_clk cell_3147 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_8739 ) ) ;
    buf_clk cell_3151 ( .C ( clk ), .D ( signal_2432 ), .Q ( signal_8743 ) ) ;
    buf_clk cell_3155 ( .C ( clk ), .D ( signal_2433 ), .Q ( signal_8747 ) ) ;
    buf_clk cell_3179 ( .C ( clk ), .D ( signal_8770 ), .Q ( signal_8771 ) ) ;
    buf_clk cell_3185 ( .C ( clk ), .D ( signal_8776 ), .Q ( signal_8777 ) ) ;
    buf_clk cell_3191 ( .C ( clk ), .D ( signal_8782 ), .Q ( signal_8783 ) ) ;
    buf_clk cell_3219 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_8811 ) ) ;
    buf_clk cell_3223 ( .C ( clk ), .D ( signal_2450 ), .Q ( signal_8815 ) ) ;
    buf_clk cell_3227 ( .C ( clk ), .D ( signal_2451 ), .Q ( signal_8819 ) ) ;
    buf_clk cell_3285 ( .C ( clk ), .D ( signal_8002 ), .Q ( signal_8877 ) ) ;
    buf_clk cell_3289 ( .C ( clk ), .D ( signal_8004 ), .Q ( signal_8881 ) ) ;
    buf_clk cell_3293 ( .C ( clk ), .D ( signal_8006 ), .Q ( signal_8885 ) ) ;
    buf_clk cell_3401 ( .C ( clk ), .D ( signal_8992 ), .Q ( signal_8993 ) ) ;
    buf_clk cell_3409 ( .C ( clk ), .D ( signal_9000 ), .Q ( signal_9001 ) ) ;
    buf_clk cell_3417 ( .C ( clk ), .D ( signal_9008 ), .Q ( signal_9009 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_988 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2431, signal_2430, signal_953}), .clk ( clk ), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_2531, signal_2530, signal_1003}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_999 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2435, signal_2434, signal_955}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({signal_2553, signal_2552, signal_1014}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1004 ( .a ({signal_7982, signal_7980, signal_7978}), .b ({signal_2431, signal_2430, signal_953}), .clk ( clk ), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_2563, signal_2562, signal_1019}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1005 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2441, signal_2440, signal_958}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({signal_2565, signal_2564, signal_1020}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1006 ( .a ({signal_7988, signal_7986, signal_7984}), .b ({signal_2431, signal_2430, signal_953}), .clk ( clk ), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_2567, signal_2566, signal_1021}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1007 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2445, signal_2444, signal_960}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({signal_2569, signal_2568, signal_1022}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1008 ( .a ({signal_2439, signal_2438, signal_957}), .b ({signal_2443, signal_2442, signal_959}), .clk ( clk ), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_2571, signal_2570, signal_1023}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1009 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({signal_2573, signal_2572, signal_1024}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1010 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_2575, signal_2574, signal_1025}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1011 ( .a ({signal_2435, signal_2434, signal_955}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({signal_2577, signal_2576, signal_1026}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1012 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_2579, signal_2578, signal_1027}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1013 ( .a ({signal_2425, signal_2424, signal_950}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({signal_2581, signal_2580, signal_1028}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1014 ( .a ({signal_8000, signal_7998, signal_7996}), .b ({signal_2445, signal_2444, signal_960}), .clk ( clk ), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_2583, signal_2582, signal_1029}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1015 ( .a ({signal_2437, signal_2436, signal_956}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({signal_2585, signal_2584, signal_1030}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1033 ( .a ({signal_2531, signal_2530, signal_1003}), .b ({signal_2621, signal_2620, signal_1048}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1040 ( .a ({signal_2553, signal_2552, signal_1014}), .b ({signal_2635, signal_2634, signal_1055}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1044 ( .a ({signal_2565, signal_2564, signal_1020}), .b ({signal_2643, signal_2642, signal_1059}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1045 ( .a ({signal_2571, signal_2570, signal_1023}), .b ({signal_2645, signal_2644, signal_1060}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1046 ( .a ({signal_2575, signal_2574, signal_1025}), .b ({signal_2647, signal_2646, signal_1061}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1047 ( .a ({signal_2577, signal_2576, signal_1026}), .b ({signal_2649, signal_2648, signal_1062}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1048 ( .a ({signal_2579, signal_2578, signal_1027}), .b ({signal_2651, signal_2650, signal_1063}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1049 ( .a ({signal_2581, signal_2580, signal_1028}), .b ({signal_2653, signal_2652, signal_1064}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1050 ( .a ({signal_2583, signal_2582, signal_1029}), .b ({signal_2655, signal_2654, signal_1065}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1051 ( .a ({signal_2585, signal_2584, signal_1030}), .b ({signal_2657, signal_2656, signal_1066}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1052 ( .a ({signal_7988, signal_7986, signal_7984}), .b ({signal_2483, signal_2482, signal_979}), .clk ( clk ), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_2659, signal_2658, signal_1067}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1053 ( .a ({signal_8006, signal_8004, signal_8002}), .b ({signal_2491, signal_2490, signal_983}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({signal_2661, signal_2660, signal_1068}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1054 ( .a ({signal_2459, signal_2458, signal_967}), .b ({signal_2461, signal_2460, signal_968}), .clk ( clk ), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_2663, signal_2662, signal_1069}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1055 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2457, signal_2456, signal_966}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({signal_2665, signal_2664, signal_1070}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1056 ( .a ({signal_8012, signal_8010, signal_8008}), .b ({signal_2485, signal_2484, signal_980}), .clk ( clk ), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_2667, signal_2666, signal_1071}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1057 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2485, signal_2484, signal_980}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({signal_2669, signal_2668, signal_1072}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1058 ( .a ({signal_2495, signal_2494, signal_985}), .b ({signal_2441, signal_2440, signal_958}), .clk ( clk ), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_2671, signal_2670, signal_1073}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1059 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2487, signal_2486, signal_981}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({signal_2673, signal_2672, signal_1074}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1060 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2517, signal_2516, signal_996}), .clk ( clk ), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_2675, signal_2674, signal_1075}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1061 ( .a ({signal_2513, signal_2512, signal_994}), .b ({signal_2523, signal_2522, signal_999}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({signal_2677, signal_2676, signal_1076}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1062 ( .a ({signal_8006, signal_8004, signal_8002}), .b ({signal_2483, signal_2482, signal_979}), .clk ( clk ), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_2679, signal_2678, signal_1077}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1063 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({signal_2681, signal_2680, signal_1078}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1064 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2529, signal_2528, signal_1002}), .clk ( clk ), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_2683, signal_2682, signal_1079}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1065 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({signal_2685, signal_2684, signal_1080}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1066 ( .a ({signal_8018, signal_8016, signal_8014}), .b ({signal_2533, signal_2532, signal_1004}), .clk ( clk ), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_2687, signal_2686, signal_1081}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1067 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2495, signal_2494, signal_985}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({signal_2689, signal_2688, signal_1082}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1068 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_2691, signal_2690, signal_1083}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1069 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2491, signal_2490, signal_983}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({signal_2693, signal_2692, signal_1084}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1070 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2521, signal_2520, signal_998}), .clk ( clk ), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_2695, signal_2694, signal_1085}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1071 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({signal_2697, signal_2696, signal_1086}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1072 ( .a ({signal_2525, signal_2524, signal_1000}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_2699, signal_2698, signal_1087}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1073 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2493, signal_2492, signal_984}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({signal_2701, signal_2700, signal_1088}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1074 ( .a ({signal_7982, signal_7980, signal_7978}), .b ({signal_2511, signal_2510, signal_993}), .clk ( clk ), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_2703, signal_2702, signal_1089}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1075 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2517, signal_2516, signal_996}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({signal_2705, signal_2704, signal_1090}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1076 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_2707, signal_2706, signal_1091}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1077 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({signal_2709, signal_2708, signal_1092}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1078 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_2711, signal_2710, signal_1093}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1079 ( .a ({signal_2425, signal_2424, signal_950}), .b ({signal_2509, signal_2508, signal_992}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({signal_2713, signal_2712, signal_1094}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1080 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2441, signal_2440, signal_958}), .clk ( clk ), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_2715, signal_2714, signal_1095}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1081 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_2549, signal_2548, signal_1012}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({signal_2717, signal_2716, signal_1096}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1082 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_2719, signal_2718, signal_1097}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1083 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2487, signal_2486, signal_981}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({signal_2721, signal_2720, signal_1098}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1084 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_2723, signal_2722, signal_1099}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1086 ( .a ({signal_2489, signal_2488, signal_982}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({signal_2727, signal_2726, signal_1101}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1087 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2489, signal_2488, signal_982}), .clk ( clk ), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_2729, signal_2728, signal_1102}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1088 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({signal_2731, signal_2730, signal_1103}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1089 ( .a ({signal_7988, signal_7986, signal_7984}), .b ({signal_2501, signal_2500, signal_988}), .clk ( clk ), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_2733, signal_2732, signal_1104}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1090 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2445, signal_2444, signal_960}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({signal_2735, signal_2734, signal_1105}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1091 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2557, signal_2556, signal_1016}), .clk ( clk ), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_2737, signal_2736, signal_1106}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1092 ( .a ({signal_8006, signal_8004, signal_8002}), .b ({signal_2533, signal_2532, signal_1004}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({signal_2739, signal_2738, signal_1107}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1093 ( .a ({signal_8024, signal_8022, signal_8020}), .b ({signal_2485, signal_2484, signal_980}), .clk ( clk ), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_2741, signal_2740, signal_1108}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1094 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2549, signal_2548, signal_1012}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({signal_2743, signal_2742, signal_1109}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1095 ( .a ({signal_2505, signal_2504, signal_990}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_2745, signal_2744, signal_1110}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1096 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2509, signal_2508, signal_992}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({signal_2747, signal_2746, signal_1111}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1097 ( .a ({signal_2447, signal_2446, signal_961}), .b ({signal_2551, signal_2550, signal_1013}), .clk ( clk ), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_2749, signal_2748, signal_1112}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1098 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({signal_2751, signal_2750, signal_1113}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1099 ( .a ({signal_8030, signal_8028, signal_8026}), .b ({signal_2545, signal_2544, signal_1010}), .clk ( clk ), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_2753, signal_2752, signal_1114}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1100 ( .a ({signal_8012, signal_8010, signal_8008}), .b ({signal_2517, signal_2516, signal_996}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({signal_2755, signal_2754, signal_1115}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1101 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2545, signal_2544, signal_1010}), .clk ( clk ), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_2757, signal_2756, signal_1116}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1102 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({signal_2759, signal_2758, signal_1117}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1103 ( .a ({signal_8018, signal_8016, signal_8014}), .b ({signal_2529, signal_2528, signal_1002}), .clk ( clk ), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_2761, signal_2760, signal_1118}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1104 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2511, signal_2510, signal_993}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({signal_2763, signal_2762, signal_1119}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1105 ( .a ({signal_8036, signal_8034, signal_8032}), .b ({signal_2491, signal_2490, signal_983}), .clk ( clk ), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_2765, signal_2764, signal_1120}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1106 ( .a ({signal_2503, signal_2502, signal_989}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({signal_2767, signal_2766, signal_1121}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1107 ( .a ({signal_2445, signal_2444, signal_960}), .b ({signal_2561, signal_2560, signal_1018}), .clk ( clk ), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_2769, signal_2768, signal_1122}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1108 ( .a ({signal_2535, signal_2534, signal_1005}), .b ({signal_2541, signal_2540, signal_1008}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({signal_2771, signal_2770, signal_1123}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1109 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2523, signal_2522, signal_999}), .clk ( clk ), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_2773, signal_2772, signal_1124}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1110 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({signal_2775, signal_2774, signal_1125}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1111 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2541, signal_2540, signal_1008}), .clk ( clk ), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_2777, signal_2776, signal_1126}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1112 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2437, signal_2436, signal_956}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({signal_2779, signal_2778, signal_1127}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1113 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_2451, signal_2450, signal_963}), .clk ( clk ), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_2781, signal_2780, signal_1128}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1114 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2557, signal_2556, signal_1016}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({signal_2783, signal_2782, signal_1129}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1115 ( .a ({signal_2433, signal_2432, signal_954}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_2785, signal_2784, signal_1130}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1116 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({signal_2787, signal_2786, signal_1131}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1117 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2497, signal_2496, signal_986}), .clk ( clk ), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_2789, signal_2788, signal_1132}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1118 ( .a ({signal_2503, signal_2502, signal_989}), .b ({signal_2505, signal_2504, signal_990}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({signal_2791, signal_2790, signal_1133}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1119 ( .a ({signal_2505, signal_2504, signal_990}), .b ({signal_2509, signal_2508, signal_992}), .clk ( clk ), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_2793, signal_2792, signal_1134}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1120 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2511, signal_2510, signal_993}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({signal_2795, signal_2794, signal_1135}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1121 ( .a ({signal_2505, signal_2504, signal_990}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_2797, signal_2796, signal_1136}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1122 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2515, signal_2514, signal_995}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({signal_2799, signal_2798, signal_1137}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1123 ( .a ({signal_8024, signal_8022, signal_8020}), .b ({signal_2519, signal_2518, signal_997}), .clk ( clk ), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_2801, signal_2800, signal_1138}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1125 ( .a ({signal_2489, signal_2488, signal_982}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({signal_2805, signal_2804, signal_1140}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1126 ( .a ({signal_2439, signal_2438, signal_957}), .b ({signal_2511, signal_2510, signal_993}), .clk ( clk ), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_2807, signal_2806, signal_1141}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1127 ( .a ({signal_2441, signal_2440, signal_958}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({signal_2809, signal_2808, signal_1142}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1128 ( .a ({signal_2527, signal_2526, signal_1001}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_2811, signal_2810, signal_1143}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1129 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2517, signal_2516, signal_996}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({signal_2813, signal_2812, signal_1144}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1130 ( .a ({signal_8018, signal_8016, signal_8014}), .b ({signal_2519, signal_2518, signal_997}), .clk ( clk ), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_2815, signal_2814, signal_1145}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1131 ( .a ({signal_2509, signal_2508, signal_992}), .b ({signal_2537, signal_2536, signal_1006}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({signal_2817, signal_2816, signal_1146}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1133 ( .a ({signal_2433, signal_2432, signal_954}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_2821, signal_2820, signal_1148}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1134 ( .a ({signal_2503, signal_2502, signal_989}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({signal_2823, signal_2822, signal_1149}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1135 ( .a ({signal_2533, signal_2532, signal_1004}), .b ({signal_2449, signal_2448, signal_962}), .clk ( clk ), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_2825, signal_2824, signal_1150}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1136 ( .a ({signal_8042, signal_8040, signal_8038}), .b ({signal_2541, signal_2540, signal_1008}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({signal_2827, signal_2826, signal_1151}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1137 ( .a ({signal_2535, signal_2534, signal_1005}), .b ({signal_2543, signal_2542, signal_1009}), .clk ( clk ), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_2829, signal_2828, signal_1152}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1138 ( .a ({signal_7988, signal_7986, signal_7984}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({signal_2831, signal_2830, signal_1153}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1139 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_2833, signal_2832, signal_1154}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1141 ( .a ({signal_2525, signal_2524, signal_1000}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({signal_2837, signal_2836, signal_1156}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1142 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_2839, signal_2838, signal_1157}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1143 ( .a ({signal_7994, signal_7992, signal_7990}), .b ({signal_2501, signal_2500, signal_988}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({signal_2841, signal_2840, signal_1158}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1144 ( .a ({signal_2495, signal_2494, signal_985}), .b ({signal_2439, signal_2438, signal_957}), .clk ( clk ), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_2843, signal_2842, signal_1159}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1145 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2511, signal_2510, signal_993}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({signal_2845, signal_2844, signal_1160}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1146 ( .a ({signal_2429, signal_2428, signal_952}), .b ({signal_2507, signal_2506, signal_991}), .clk ( clk ), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_2847, signal_2846, signal_1161}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1147 ( .a ({signal_2495, signal_2494, signal_985}), .b ({signal_2517, signal_2516, signal_996}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({signal_2849, signal_2848, signal_1162}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1148 ( .a ({signal_2457, signal_2456, signal_966}), .b ({signal_2471, signal_2470, signal_973}), .clk ( clk ), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_2851, signal_2850, signal_1163}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1149 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({signal_2853, signal_2852, signal_1164}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1150 ( .a ({signal_2509, signal_2508, signal_992}), .b ({signal_2547, signal_2546, signal_1011}), .clk ( clk ), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_2855, signal_2854, signal_1165}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1151 ( .a ({signal_2489, signal_2488, signal_982}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({signal_2857, signal_2856, signal_1166}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1152 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2519, signal_2518, signal_997}), .clk ( clk ), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_2859, signal_2858, signal_1167}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1153 ( .a ({signal_8042, signal_8040, signal_8038}), .b ({signal_2513, signal_2512, signal_994}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({signal_2861, signal_2860, signal_1168}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1154 ( .a ({signal_2439, signal_2438, signal_957}), .b ({signal_2545, signal_2544, signal_1010}), .clk ( clk ), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_2863, signal_2862, signal_1169}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1156 ( .a ({signal_2537, signal_2536, signal_1006}), .b ({signal_2545, signal_2544, signal_1010}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({signal_2867, signal_2866, signal_1171}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1157 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2507, signal_2506, signal_991}), .clk ( clk ), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_2869, signal_2868, signal_1172}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1158 ( .a ({signal_2519, signal_2518, signal_997}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({signal_2871, signal_2870, signal_1173}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1159 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2541, signal_2540, signal_1008}), .clk ( clk ), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_2873, signal_2872, signal_1174}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1160 ( .a ({signal_8024, signal_8022, signal_8020}), .b ({signal_2501, signal_2500, signal_988}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({signal_2875, signal_2874, signal_1175}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1161 ( .a ({signal_8012, signal_8010, signal_8008}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_2877, signal_2876, signal_1176}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1162 ( .a ({signal_8006, signal_8004, signal_8002}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({signal_2879, signal_2878, signal_1177}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1163 ( .a ({signal_2515, signal_2514, signal_995}), .b ({signal_2555, signal_2554, signal_1015}), .clk ( clk ), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_2881, signal_2880, signal_1178}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1164 ( .a ({signal_2457, signal_2456, signal_966}), .b ({signal_2469, signal_2468, signal_972}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({signal_2883, signal_2882, signal_1179}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1165 ( .a ({signal_2467, signal_2466, signal_971}), .b ({signal_2469, signal_2468, signal_972}), .clk ( clk ), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_2885, signal_2884, signal_1180}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1166 ( .a ({signal_2449, signal_2448, signal_962}), .b ({signal_2549, signal_2548, signal_1012}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({signal_2887, signal_2886, signal_1181}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1167 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2507, signal_2506, signal_991}), .clk ( clk ), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_2889, signal_2888, signal_1182}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1168 ( .a ({signal_2435, signal_2434, signal_955}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({signal_2891, signal_2890, signal_1183}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1169 ( .a ({signal_8000, signal_7998, signal_7996}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_2893, signal_2892, signal_1184}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1170 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2525, signal_2524, signal_1000}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({signal_2895, signal_2894, signal_1185}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1171 ( .a ({signal_2449, signal_2448, signal_962}), .b ({signal_2555, signal_2554, signal_1015}), .clk ( clk ), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_2897, signal_2896, signal_1186}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1172 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2515, signal_2514, signal_995}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({signal_2899, signal_2898, signal_1187}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1174 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2493, signal_2492, signal_984}), .clk ( clk ), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_2903, signal_2902, signal_1189}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1175 ( .a ({signal_2491, signal_2490, signal_983}), .b ({signal_2533, signal_2532, signal_1004}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({signal_2905, signal_2904, signal_1190}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1176 ( .a ({signal_2427, signal_2426, signal_951}), .b ({signal_2507, signal_2506, signal_991}), .clk ( clk ), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_2907, signal_2906, signal_1191}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1177 ( .a ({signal_2517, signal_2516, signal_996}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({signal_2909, signal_2908, signal_1192}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1178 ( .a ({signal_2463, signal_2462, signal_969}), .b ({signal_2477, signal_2476, signal_976}), .clk ( clk ), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_2911, signal_2910, signal_1193}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1179 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2507, signal_2506, signal_991}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({signal_2913, signal_2912, signal_1194}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1180 ( .a ({signal_2499, signal_2498, signal_987}), .b ({signal_2439, signal_2438, signal_957}), .clk ( clk ), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_2915, signal_2914, signal_1195}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1181 ( .a ({signal_2449, signal_2448, signal_962}), .b ({signal_2543, signal_2542, signal_1009}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({signal_2917, signal_2916, signal_1196}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1182 ( .a ({signal_8018, signal_8016, signal_8014}), .b ({signal_2543, signal_2542, signal_1009}), .clk ( clk ), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_2919, signal_2918, signal_1197}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1183 ( .a ({signal_2485, signal_2484, signal_980}), .b ({signal_2447, signal_2446, signal_961}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({signal_2921, signal_2920, signal_1198}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1185 ( .a ({signal_2493, signal_2492, signal_984}), .b ({signal_2555, signal_2554, signal_1015}), .clk ( clk ), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_2925, signal_2924, signal_1200}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1186 ( .a ({signal_2521, signal_2520, signal_998}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({signal_2927, signal_2926, signal_1201}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1187 ( .a ({signal_8042, signal_8040, signal_8038}), .b ({signal_2495, signal_2494, signal_985}), .clk ( clk ), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_2929, signal_2928, signal_1202}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1188 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2443, signal_2442, signal_959}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({signal_2931, signal_2930, signal_1203}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1191 ( .a ({signal_2487, signal_2486, signal_981}), .b ({signal_2499, signal_2498, signal_987}), .clk ( clk ), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_2937, signal_2936, signal_1206}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1192 ( .a ({signal_2521, signal_2520, signal_998}), .b ({signal_2543, signal_2542, signal_1009}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({signal_2939, signal_2938, signal_1207}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1193 ( .a ({signal_2439, signal_2438, signal_957}), .b ({signal_2509, signal_2508, signal_992}), .clk ( clk ), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_2941, signal_2940, signal_1208}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1194 ( .a ({signal_2497, signal_2496, signal_986}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({signal_2943, signal_2942, signal_1209}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1195 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_2945, signal_2944, signal_1210}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1196 ( .a ({signal_2503, signal_2502, signal_989}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({signal_2947, signal_2946, signal_1211}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1197 ( .a ({signal_2495, signal_2494, signal_985}), .b ({signal_2497, signal_2496, signal_986}), .clk ( clk ), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_2949, signal_2948, signal_1212}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1199 ( .a ({signal_2507, signal_2506, signal_991}), .b ({signal_2509, signal_2508, signal_992}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({signal_2953, signal_2952, signal_1214}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1200 ( .a ({signal_2431, signal_2430, signal_953}), .b ({signal_2539, signal_2538, signal_1007}), .clk ( clk ), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_2955, signal_2954, signal_1215}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1201 ( .a ({signal_2511, signal_2510, signal_993}), .b ({signal_2521, signal_2520, signal_998}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({signal_2957, signal_2956, signal_1216}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1202 ( .a ({signal_2501, signal_2500, signal_988}), .b ({signal_2527, signal_2526, signal_1001}), .clk ( clk ), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_2959, signal_2958, signal_1217}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1203 ( .a ({signal_2515, signal_2514, signal_995}), .b ({signal_2519, signal_2518, signal_997}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({signal_2961, signal_2960, signal_1218}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1204 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_2503, signal_2502, signal_989}), .clk ( clk ), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_2963, signal_2962, signal_1219}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1205 ( .a ({signal_8030, signal_8028, signal_8026}), .b ({signal_2519, signal_2518, signal_997}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({signal_2965, signal_2964, signal_1220}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1206 ( .a ({signal_8000, signal_7998, signal_7996}), .b ({signal_2543, signal_2542, signal_1009}), .clk ( clk ), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_2967, signal_2966, signal_1221}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1208 ( .a ({signal_2533, signal_2532, signal_1004}), .b ({signal_2535, signal_2534, signal_1005}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({signal_2971, signal_2970, signal_1223}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1210 ( .a ({signal_8036, signal_8034, signal_8032}), .b ({signal_2465, signal_2464, signal_970}), .clk ( clk ), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_2975, signal_2974, signal_1225}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1213 ( .a ({signal_2483, signal_2482, signal_979}), .b ({signal_8048, signal_8046, signal_8044}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({signal_2981, signal_2980, signal_1228}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1214 ( .a ({signal_8036, signal_8034, signal_8032}), .b ({signal_2469, signal_2468, signal_972}), .clk ( clk ), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_2983, signal_2982, signal_1229}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1215 ( .a ({signal_2663, signal_2662, signal_1069}), .b ({signal_2985, signal_2984, signal_1230}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1216 ( .a ({signal_2665, signal_2664, signal_1070}), .b ({signal_2987, signal_2986, signal_1231}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1217 ( .a ({signal_2669, signal_2668, signal_1072}), .b ({signal_2989, signal_2988, signal_1232}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1218 ( .a ({signal_2671, signal_2670, signal_1073}), .b ({signal_2991, signal_2990, signal_1233}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1219 ( .a ({signal_2673, signal_2672, signal_1074}), .b ({signal_2993, signal_2992, signal_1234}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1220 ( .a ({signal_2675, signal_2674, signal_1075}), .b ({signal_2995, signal_2994, signal_1235}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1221 ( .a ({signal_2677, signal_2676, signal_1076}), .b ({signal_2997, signal_2996, signal_1236}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1222 ( .a ({signal_2679, signal_2678, signal_1077}), .b ({signal_2999, signal_2998, signal_1237}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1223 ( .a ({signal_2681, signal_2680, signal_1078}), .b ({signal_3001, signal_3000, signal_1238}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1224 ( .a ({signal_2683, signal_2682, signal_1079}), .b ({signal_3003, signal_3002, signal_1239}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1225 ( .a ({signal_2685, signal_2684, signal_1080}), .b ({signal_3005, signal_3004, signal_1240}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1226 ( .a ({signal_2687, signal_2686, signal_1081}), .b ({signal_3007, signal_3006, signal_1241}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1227 ( .a ({signal_2689, signal_2688, signal_1082}), .b ({signal_3009, signal_3008, signal_1242}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1228 ( .a ({signal_2691, signal_2690, signal_1083}), .b ({signal_3011, signal_3010, signal_1243}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1229 ( .a ({signal_2693, signal_2692, signal_1084}), .b ({signal_3013, signal_3012, signal_1244}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1230 ( .a ({signal_2697, signal_2696, signal_1086}), .b ({signal_3015, signal_3014, signal_1245}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1231 ( .a ({signal_2699, signal_2698, signal_1087}), .b ({signal_3017, signal_3016, signal_1246}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1232 ( .a ({signal_2701, signal_2700, signal_1088}), .b ({signal_3019, signal_3018, signal_1247}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1233 ( .a ({signal_2705, signal_2704, signal_1090}), .b ({signal_3021, signal_3020, signal_1248}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1234 ( .a ({signal_2707, signal_2706, signal_1091}), .b ({signal_3023, signal_3022, signal_1249}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1235 ( .a ({signal_2709, signal_2708, signal_1092}), .b ({signal_3025, signal_3024, signal_1250}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1236 ( .a ({signal_2711, signal_2710, signal_1093}), .b ({signal_3027, signal_3026, signal_1251}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1237 ( .a ({signal_2713, signal_2712, signal_1094}), .b ({signal_3029, signal_3028, signal_1252}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1238 ( .a ({signal_2715, signal_2714, signal_1095}), .b ({signal_3031, signal_3030, signal_1253}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1239 ( .a ({signal_2717, signal_2716, signal_1096}), .b ({signal_3033, signal_3032, signal_1254}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1240 ( .a ({signal_2719, signal_2718, signal_1097}), .b ({signal_3035, signal_3034, signal_1255}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1241 ( .a ({signal_2721, signal_2720, signal_1098}), .b ({signal_3037, signal_3036, signal_1256}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1242 ( .a ({signal_2723, signal_2722, signal_1099}), .b ({signal_3039, signal_3038, signal_1257}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1244 ( .a ({signal_2727, signal_2726, signal_1101}), .b ({signal_3043, signal_3042, signal_1259}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1245 ( .a ({signal_2731, signal_2730, signal_1103}), .b ({signal_3045, signal_3044, signal_1260}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1246 ( .a ({signal_2735, signal_2734, signal_1105}), .b ({signal_3047, signal_3046, signal_1261}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1247 ( .a ({signal_2737, signal_2736, signal_1106}), .b ({signal_3049, signal_3048, signal_1262}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1248 ( .a ({signal_2741, signal_2740, signal_1108}), .b ({signal_3051, signal_3050, signal_1263}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1249 ( .a ({signal_2743, signal_2742, signal_1109}), .b ({signal_3053, signal_3052, signal_1264}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1250 ( .a ({signal_2745, signal_2744, signal_1110}), .b ({signal_3055, signal_3054, signal_1265}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1251 ( .a ({signal_2747, signal_2746, signal_1111}), .b ({signal_3057, signal_3056, signal_1266}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1252 ( .a ({signal_2749, signal_2748, signal_1112}), .b ({signal_3059, signal_3058, signal_1267}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1253 ( .a ({signal_2751, signal_2750, signal_1113}), .b ({signal_3061, signal_3060, signal_1268}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1254 ( .a ({signal_2755, signal_2754, signal_1115}), .b ({signal_3063, signal_3062, signal_1269}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1255 ( .a ({signal_2757, signal_2756, signal_1116}), .b ({signal_3065, signal_3064, signal_1270}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1256 ( .a ({signal_2759, signal_2758, signal_1117}), .b ({signal_3067, signal_3066, signal_1271}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1257 ( .a ({signal_2761, signal_2760, signal_1118}), .b ({signal_3069, signal_3068, signal_1272}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1258 ( .a ({signal_2765, signal_2764, signal_1120}), .b ({signal_3071, signal_3070, signal_1273}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1259 ( .a ({signal_2767, signal_2766, signal_1121}), .b ({signal_3073, signal_3072, signal_1274}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1260 ( .a ({signal_2769, signal_2768, signal_1122}), .b ({signal_3075, signal_3074, signal_1275}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1261 ( .a ({signal_2773, signal_2772, signal_1124}), .b ({signal_3077, signal_3076, signal_1276}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1262 ( .a ({signal_2775, signal_2774, signal_1125}), .b ({signal_3079, signal_3078, signal_1277}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1263 ( .a ({signal_2777, signal_2776, signal_1126}), .b ({signal_3081, signal_3080, signal_1278}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1264 ( .a ({signal_2779, signal_2778, signal_1127}), .b ({signal_3083, signal_3082, signal_1279}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1265 ( .a ({signal_2783, signal_2782, signal_1129}), .b ({signal_3085, signal_3084, signal_1280}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1266 ( .a ({signal_2785, signal_2784, signal_1130}), .b ({signal_3087, signal_3086, signal_1281}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1267 ( .a ({signal_2787, signal_2786, signal_1131}), .b ({signal_3089, signal_3088, signal_1282}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1268 ( .a ({signal_2793, signal_2792, signal_1134}), .b ({signal_3091, signal_3090, signal_1283}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1269 ( .a ({signal_2795, signal_2794, signal_1135}), .b ({signal_3093, signal_3092, signal_1284}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1270 ( .a ({signal_2797, signal_2796, signal_1136}), .b ({signal_3095, signal_3094, signal_1285}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1271 ( .a ({signal_2799, signal_2798, signal_1137}), .b ({signal_3097, signal_3096, signal_1286}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1273 ( .a ({signal_2807, signal_2806, signal_1141}), .b ({signal_3101, signal_3100, signal_1288}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1274 ( .a ({signal_2811, signal_2810, signal_1143}), .b ({signal_3103, signal_3102, signal_1289}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1275 ( .a ({signal_2813, signal_2812, signal_1144}), .b ({signal_3105, signal_3104, signal_1290}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1276 ( .a ({signal_2817, signal_2816, signal_1146}), .b ({signal_3107, signal_3106, signal_1291}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1278 ( .a ({signal_2821, signal_2820, signal_1148}), .b ({signal_3111, signal_3110, signal_1293}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1279 ( .a ({signal_2823, signal_2822, signal_1149}), .b ({signal_3113, signal_3112, signal_1294}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1280 ( .a ({signal_2825, signal_2824, signal_1150}), .b ({signal_3115, signal_3114, signal_1295}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1281 ( .a ({signal_2829, signal_2828, signal_1152}), .b ({signal_3117, signal_3116, signal_1296}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1282 ( .a ({signal_2831, signal_2830, signal_1153}), .b ({signal_3119, signal_3118, signal_1297}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1283 ( .a ({signal_2833, signal_2832, signal_1154}), .b ({signal_3121, signal_3120, signal_1298}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1285 ( .a ({signal_2837, signal_2836, signal_1156}), .b ({signal_3125, signal_3124, signal_1300}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1286 ( .a ({signal_2839, signal_2838, signal_1157}), .b ({signal_3127, signal_3126, signal_1301}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1287 ( .a ({signal_2843, signal_2842, signal_1159}), .b ({signal_3129, signal_3128, signal_1302}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1288 ( .a ({signal_2845, signal_2844, signal_1160}), .b ({signal_3131, signal_3130, signal_1303}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1289 ( .a ({signal_2847, signal_2846, signal_1161}), .b ({signal_3133, signal_3132, signal_1304}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1290 ( .a ({signal_2849, signal_2848, signal_1162}), .b ({signal_3135, signal_3134, signal_1305}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1291 ( .a ({signal_2851, signal_2850, signal_1163}), .b ({signal_3137, signal_3136, signal_1306}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1292 ( .a ({signal_2853, signal_2852, signal_1164}), .b ({signal_3139, signal_3138, signal_1307}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1293 ( .a ({signal_2855, signal_2854, signal_1165}), .b ({signal_3141, signal_3140, signal_1308}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1294 ( .a ({signal_2857, signal_2856, signal_1166}), .b ({signal_3143, signal_3142, signal_1309}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1295 ( .a ({signal_2859, signal_2858, signal_1167}), .b ({signal_3145, signal_3144, signal_1310}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1296 ( .a ({signal_2863, signal_2862, signal_1169}), .b ({signal_3147, signal_3146, signal_1311}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1298 ( .a ({signal_2867, signal_2866, signal_1171}), .b ({signal_3151, signal_3150, signal_1313}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1299 ( .a ({signal_2869, signal_2868, signal_1172}), .b ({signal_3153, signal_3152, signal_1314}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1300 ( .a ({signal_2871, signal_2870, signal_1173}), .b ({signal_3155, signal_3154, signal_1315}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1301 ( .a ({signal_2873, signal_2872, signal_1174}), .b ({signal_3157, signal_3156, signal_1316}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1302 ( .a ({signal_2875, signal_2874, signal_1175}), .b ({signal_3159, signal_3158, signal_1317}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1303 ( .a ({signal_2877, signal_2876, signal_1176}), .b ({signal_3161, signal_3160, signal_1318}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1304 ( .a ({signal_2879, signal_2878, signal_1177}), .b ({signal_3163, signal_3162, signal_1319}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1305 ( .a ({signal_2883, signal_2882, signal_1179}), .b ({signal_3165, signal_3164, signal_1320}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1306 ( .a ({signal_2885, signal_2884, signal_1180}), .b ({signal_3167, signal_3166, signal_1321}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1307 ( .a ({signal_2887, signal_2886, signal_1181}), .b ({signal_3169, signal_3168, signal_1322}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1308 ( .a ({signal_2889, signal_2888, signal_1182}), .b ({signal_3171, signal_3170, signal_1323}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1309 ( .a ({signal_2891, signal_2890, signal_1183}), .b ({signal_3173, signal_3172, signal_1324}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1310 ( .a ({signal_2893, signal_2892, signal_1184}), .b ({signal_3175, signal_3174, signal_1325}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1311 ( .a ({signal_2895, signal_2894, signal_1185}), .b ({signal_3177, signal_3176, signal_1326}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1312 ( .a ({signal_2897, signal_2896, signal_1186}), .b ({signal_3179, signal_3178, signal_1327}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1313 ( .a ({signal_2899, signal_2898, signal_1187}), .b ({signal_3181, signal_3180, signal_1328}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1315 ( .a ({signal_2903, signal_2902, signal_1189}), .b ({signal_3185, signal_3184, signal_1330}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1316 ( .a ({signal_2907, signal_2906, signal_1191}), .b ({signal_3187, signal_3186, signal_1331}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1317 ( .a ({signal_2909, signal_2908, signal_1192}), .b ({signal_3189, signal_3188, signal_1332}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1318 ( .a ({signal_2911, signal_2910, signal_1193}), .b ({signal_3191, signal_3190, signal_1333}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1319 ( .a ({signal_2913, signal_2912, signal_1194}), .b ({signal_3193, signal_3192, signal_1334}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1320 ( .a ({signal_2915, signal_2914, signal_1195}), .b ({signal_3195, signal_3194, signal_1335}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1321 ( .a ({signal_2917, signal_2916, signal_1196}), .b ({signal_3197, signal_3196, signal_1336}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1322 ( .a ({signal_2919, signal_2918, signal_1197}), .b ({signal_3199, signal_3198, signal_1337}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1324 ( .a ({signal_2925, signal_2924, signal_1200}), .b ({signal_3203, signal_3202, signal_1339}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1325 ( .a ({signal_2927, signal_2926, signal_1201}), .b ({signal_3205, signal_3204, signal_1340}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1326 ( .a ({signal_2929, signal_2928, signal_1202}), .b ({signal_3207, signal_3206, signal_1341}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1327 ( .a ({signal_2931, signal_2930, signal_1203}), .b ({signal_3209, signal_3208, signal_1342}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1330 ( .a ({signal_2939, signal_2938, signal_1207}), .b ({signal_3215, signal_3214, signal_1345}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1331 ( .a ({signal_2943, signal_2942, signal_1209}), .b ({signal_3217, signal_3216, signal_1346}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1332 ( .a ({signal_2945, signal_2944, signal_1210}), .b ({signal_3219, signal_3218, signal_1347}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1333 ( .a ({signal_2947, signal_2946, signal_1211}), .b ({signal_3221, signal_3220, signal_1348}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1334 ( .a ({signal_2949, signal_2948, signal_1212}), .b ({signal_3223, signal_3222, signal_1349}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1336 ( .a ({signal_2953, signal_2952, signal_1214}), .b ({signal_3227, signal_3226, signal_1351}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1337 ( .a ({signal_2955, signal_2954, signal_1215}), .b ({signal_3229, signal_3228, signal_1352}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1338 ( .a ({signal_2957, signal_2956, signal_1216}), .b ({signal_3231, signal_3230, signal_1353}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1339 ( .a ({signal_2961, signal_2960, signal_1218}), .b ({signal_3233, signal_3232, signal_1354}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1340 ( .a ({signal_2963, signal_2962, signal_1219}), .b ({signal_3235, signal_3234, signal_1355}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1341 ( .a ({signal_2965, signal_2964, signal_1220}), .b ({signal_3237, signal_3236, signal_1356}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1342 ( .a ({signal_2967, signal_2966, signal_1221}), .b ({signal_3239, signal_3238, signal_1357}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1344 ( .a ({signal_2971, signal_2970, signal_1223}), .b ({signal_3243, signal_3242, signal_1359}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1346 ( .a ({signal_2975, signal_2974, signal_1225}), .b ({signal_3247, signal_3246, signal_1361}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1349 ( .a ({signal_2981, signal_2980, signal_1228}), .b ({signal_3253, signal_3252, signal_1364}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1350 ( .a ({signal_2983, signal_2982, signal_1229}), .b ({signal_3255, signal_3254, signal_1365}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1353 ( .a ({signal_8054, signal_8052, signal_8050}), .b ({signal_2617, signal_2616, signal_1046}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({signal_3261, signal_3260, signal_1368}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1354 ( .a ({signal_8024, signal_8022, signal_8020}), .b ({signal_2609, signal_2608, signal_1042}), .clk ( clk ), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_3263, signal_3262, signal_1369}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1355 ( .a ({signal_2587, signal_2586, signal_1031}), .b ({signal_2641, signal_2640, signal_1058}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({signal_3265, signal_3264, signal_1370}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1356 ( .a ({signal_2615, signal_2614, signal_1045}), .b ({signal_2639, signal_2638, signal_1057}), .clk ( clk ), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_3267, signal_3266, signal_1371}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1357 ( .a ({signal_2597, signal_2596, signal_1036}), .b ({signal_2599, signal_2598, signal_1037}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({signal_3269, signal_3268, signal_1372}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1360 ( .a ({signal_2597, signal_2596, signal_1036}), .b ({signal_2615, signal_2614, signal_1045}), .clk ( clk ), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_3275, signal_3274, signal_1375}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1361 ( .a ({signal_2607, signal_2606, signal_1041}), .b ({signal_2629, signal_2628, signal_1052}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({signal_3277, signal_3276, signal_1376}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1362 ( .a ({signal_2627, signal_2626, signal_1051}), .b ({signal_2631, signal_2630, signal_1053}), .clk ( clk ), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_3279, signal_3278, signal_1377}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1365 ( .a ({signal_2587, signal_2586, signal_1031}), .b ({signal_2613, signal_2612, signal_1044}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({signal_3285, signal_3284, signal_1380}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1366 ( .a ({signal_2589, signal_2588, signal_1032}), .b ({signal_2629, signal_2628, signal_1052}), .clk ( clk ), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_3287, signal_3286, signal_1381}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1367 ( .a ({signal_2609, signal_2608, signal_1042}), .b ({signal_2611, signal_2610, signal_1043}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({signal_3289, signal_3288, signal_1382}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1368 ( .a ({signal_2599, signal_2598, signal_1037}), .b ({signal_2615, signal_2614, signal_1045}), .clk ( clk ), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_3291, signal_3290, signal_1383}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1369 ( .a ({signal_2473, signal_2472, signal_974}), .b ({signal_2631, signal_2630, signal_1053}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({signal_3293, signal_3292, signal_1384}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1375 ( .a ({signal_2605, signal_2604, signal_1040}), .b ({signal_2637, signal_2636, signal_1056}), .clk ( clk ), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_3305, signal_3304, signal_1390}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1376 ( .a ({signal_2615, signal_2614, signal_1045}), .b ({signal_2625, signal_2624, signal_1050}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({signal_3307, signal_3306, signal_1391}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1383 ( .a ({signal_2591, signal_2590, signal_1033}), .b ({signal_2595, signal_2594, signal_1035}), .clk ( clk ), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_3321, signal_3320, signal_1398}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1395 ( .a ({signal_2467, signal_2466, signal_971}), .b ({signal_2623, signal_2622, signal_1049}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({signal_3345, signal_3344, signal_1410}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1396 ( .a ({signal_2589, signal_2588, signal_1032}), .b ({signal_2619, signal_2618, signal_1047}), .clk ( clk ), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_3347, signal_3346, signal_1411}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1401 ( .a ({signal_2459, signal_2458, signal_967}), .b ({signal_2611, signal_2610, signal_1043}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({signal_3357, signal_3356, signal_1416}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1402 ( .a ({signal_2625, signal_2624, signal_1050}), .b ({signal_2475, signal_2474, signal_975}), .clk ( clk ), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_3359, signal_3358, signal_1417}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1403 ( .a ({signal_2469, signal_2468, signal_972}), .b ({signal_2615, signal_2614, signal_1045}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({signal_3361, signal_3360, signal_1418}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1407 ( .a ({signal_2601, signal_2600, signal_1038}), .b ({signal_2617, signal_2616, signal_1046}), .clk ( clk ), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_3369, signal_3368, signal_1422}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1408 ( .a ({signal_2605, signal_2604, signal_1040}), .b ({signal_2475, signal_2474, signal_975}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({signal_3371, signal_3370, signal_1423}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1492 ( .a ({signal_3261, signal_3260, signal_1368}), .b ({signal_3539, signal_3538, signal_1507}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1493 ( .a ({signal_3263, signal_3262, signal_1369}), .b ({signal_3541, signal_3540, signal_1508}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1494 ( .a ({signal_3265, signal_3264, signal_1370}), .b ({signal_3543, signal_3542, signal_1509}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1495 ( .a ({signal_3267, signal_3266, signal_1371}), .b ({signal_3545, signal_3544, signal_1510}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1496 ( .a ({signal_3269, signal_3268, signal_1372}), .b ({signal_3547, signal_3546, signal_1511}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1499 ( .a ({signal_3275, signal_3274, signal_1375}), .b ({signal_3553, signal_3552, signal_1514}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1500 ( .a ({signal_3277, signal_3276, signal_1376}), .b ({signal_3555, signal_3554, signal_1515}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1501 ( .a ({signal_3279, signal_3278, signal_1377}), .b ({signal_3557, signal_3556, signal_1516}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1504 ( .a ({signal_3285, signal_3284, signal_1380}), .b ({signal_3563, signal_3562, signal_1519}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1505 ( .a ({signal_3287, signal_3286, signal_1381}), .b ({signal_3565, signal_3564, signal_1520}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1506 ( .a ({signal_3289, signal_3288, signal_1382}), .b ({signal_3567, signal_3566, signal_1521}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1507 ( .a ({signal_3293, signal_3292, signal_1384}), .b ({signal_3569, signal_3568, signal_1522}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1513 ( .a ({signal_3307, signal_3306, signal_1391}), .b ({signal_3581, signal_3580, signal_1528}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1520 ( .a ({signal_3321, signal_3320, signal_1398}), .b ({signal_3595, signal_3594, signal_1535}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1532 ( .a ({signal_3345, signal_3344, signal_1410}), .b ({signal_3619, signal_3618, signal_1547}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1533 ( .a ({signal_3347, signal_3346, signal_1411}), .b ({signal_3621, signal_3620, signal_1548}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1538 ( .a ({signal_3357, signal_3356, signal_1416}), .b ({signal_3631, signal_3630, signal_1553}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1539 ( .a ({signal_3359, signal_3358, signal_1417}), .b ({signal_3633, signal_3632, signal_1554}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1543 ( .a ({signal_3369, signal_3368, signal_1422}), .b ({signal_3641, signal_3640, signal_1558}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1544 ( .a ({signal_3371, signal_3370, signal_1423}), .b ({signal_3643, signal_3642, signal_1559}) ) ;
    buf_clk cell_2466 ( .C ( clk ), .D ( signal_8057 ), .Q ( signal_8058 ) ) ;
    buf_clk cell_2470 ( .C ( clk ), .D ( signal_8061 ), .Q ( signal_8062 ) ) ;
    buf_clk cell_2474 ( .C ( clk ), .D ( signal_8065 ), .Q ( signal_8066 ) ) ;
    buf_clk cell_2476 ( .C ( clk ), .D ( signal_8067 ), .Q ( signal_8068 ) ) ;
    buf_clk cell_2478 ( .C ( clk ), .D ( signal_8069 ), .Q ( signal_8070 ) ) ;
    buf_clk cell_2480 ( .C ( clk ), .D ( signal_8071 ), .Q ( signal_8072 ) ) ;
    buf_clk cell_2482 ( .C ( clk ), .D ( signal_8073 ), .Q ( signal_8074 ) ) ;
    buf_clk cell_2484 ( .C ( clk ), .D ( signal_8075 ), .Q ( signal_8076 ) ) ;
    buf_clk cell_2486 ( .C ( clk ), .D ( signal_8077 ), .Q ( signal_8078 ) ) ;
    buf_clk cell_2488 ( .C ( clk ), .D ( signal_8079 ), .Q ( signal_8080 ) ) ;
    buf_clk cell_2490 ( .C ( clk ), .D ( signal_8081 ), .Q ( signal_8082 ) ) ;
    buf_clk cell_2492 ( .C ( clk ), .D ( signal_8083 ), .Q ( signal_8084 ) ) ;
    buf_clk cell_2494 ( .C ( clk ), .D ( signal_8085 ), .Q ( signal_8086 ) ) ;
    buf_clk cell_2496 ( .C ( clk ), .D ( signal_8087 ), .Q ( signal_8088 ) ) ;
    buf_clk cell_2498 ( .C ( clk ), .D ( signal_8089 ), .Q ( signal_8090 ) ) ;
    buf_clk cell_2500 ( .C ( clk ), .D ( signal_8091 ), .Q ( signal_8092 ) ) ;
    buf_clk cell_2502 ( .C ( clk ), .D ( signal_8093 ), .Q ( signal_8094 ) ) ;
    buf_clk cell_2504 ( .C ( clk ), .D ( signal_8095 ), .Q ( signal_8096 ) ) ;
    buf_clk cell_2506 ( .C ( clk ), .D ( signal_8097 ), .Q ( signal_8098 ) ) ;
    buf_clk cell_2508 ( .C ( clk ), .D ( signal_8099 ), .Q ( signal_8100 ) ) ;
    buf_clk cell_2510 ( .C ( clk ), .D ( signal_8101 ), .Q ( signal_8102 ) ) ;
    buf_clk cell_2512 ( .C ( clk ), .D ( signal_8103 ), .Q ( signal_8104 ) ) ;
    buf_clk cell_2514 ( .C ( clk ), .D ( signal_8105 ), .Q ( signal_8106 ) ) ;
    buf_clk cell_2516 ( .C ( clk ), .D ( signal_8107 ), .Q ( signal_8108 ) ) ;
    buf_clk cell_2518 ( .C ( clk ), .D ( signal_8109 ), .Q ( signal_8110 ) ) ;
    buf_clk cell_2520 ( .C ( clk ), .D ( signal_8111 ), .Q ( signal_8112 ) ) ;
    buf_clk cell_2522 ( .C ( clk ), .D ( signal_8113 ), .Q ( signal_8114 ) ) ;
    buf_clk cell_2524 ( .C ( clk ), .D ( signal_8115 ), .Q ( signal_8116 ) ) ;
    buf_clk cell_2526 ( .C ( clk ), .D ( signal_8117 ), .Q ( signal_8118 ) ) ;
    buf_clk cell_2528 ( .C ( clk ), .D ( signal_8119 ), .Q ( signal_8120 ) ) ;
    buf_clk cell_2530 ( .C ( clk ), .D ( signal_8121 ), .Q ( signal_8122 ) ) ;
    buf_clk cell_2532 ( .C ( clk ), .D ( signal_8123 ), .Q ( signal_8124 ) ) ;
    buf_clk cell_2534 ( .C ( clk ), .D ( signal_8125 ), .Q ( signal_8126 ) ) ;
    buf_clk cell_2536 ( .C ( clk ), .D ( signal_8127 ), .Q ( signal_8128 ) ) ;
    buf_clk cell_2538 ( .C ( clk ), .D ( signal_8129 ), .Q ( signal_8130 ) ) ;
    buf_clk cell_2540 ( .C ( clk ), .D ( signal_8131 ), .Q ( signal_8132 ) ) ;
    buf_clk cell_2542 ( .C ( clk ), .D ( signal_8133 ), .Q ( signal_8134 ) ) ;
    buf_clk cell_2544 ( .C ( clk ), .D ( signal_8135 ), .Q ( signal_8136 ) ) ;
    buf_clk cell_2546 ( .C ( clk ), .D ( signal_8137 ), .Q ( signal_8138 ) ) ;
    buf_clk cell_2548 ( .C ( clk ), .D ( signal_8139 ), .Q ( signal_8140 ) ) ;
    buf_clk cell_2550 ( .C ( clk ), .D ( signal_8141 ), .Q ( signal_8142 ) ) ;
    buf_clk cell_2552 ( .C ( clk ), .D ( signal_8143 ), .Q ( signal_8144 ) ) ;
    buf_clk cell_2554 ( .C ( clk ), .D ( signal_8145 ), .Q ( signal_8146 ) ) ;
    buf_clk cell_2556 ( .C ( clk ), .D ( signal_8147 ), .Q ( signal_8148 ) ) ;
    buf_clk cell_2558 ( .C ( clk ), .D ( signal_8149 ), .Q ( signal_8150 ) ) ;
    buf_clk cell_2560 ( .C ( clk ), .D ( signal_8151 ), .Q ( signal_8152 ) ) ;
    buf_clk cell_2562 ( .C ( clk ), .D ( signal_8153 ), .Q ( signal_8154 ) ) ;
    buf_clk cell_2564 ( .C ( clk ), .D ( signal_8155 ), .Q ( signal_8156 ) ) ;
    buf_clk cell_2566 ( .C ( clk ), .D ( signal_8157 ), .Q ( signal_8158 ) ) ;
    buf_clk cell_2568 ( .C ( clk ), .D ( signal_8159 ), .Q ( signal_8160 ) ) ;
    buf_clk cell_2570 ( .C ( clk ), .D ( signal_8161 ), .Q ( signal_8162 ) ) ;
    buf_clk cell_2572 ( .C ( clk ), .D ( signal_8163 ), .Q ( signal_8164 ) ) ;
    buf_clk cell_2574 ( .C ( clk ), .D ( signal_8165 ), .Q ( signal_8166 ) ) ;
    buf_clk cell_2576 ( .C ( clk ), .D ( signal_8167 ), .Q ( signal_8168 ) ) ;
    buf_clk cell_2578 ( .C ( clk ), .D ( signal_8169 ), .Q ( signal_8170 ) ) ;
    buf_clk cell_2580 ( .C ( clk ), .D ( signal_8171 ), .Q ( signal_8172 ) ) ;
    buf_clk cell_2582 ( .C ( clk ), .D ( signal_8173 ), .Q ( signal_8174 ) ) ;
    buf_clk cell_2584 ( .C ( clk ), .D ( signal_8175 ), .Q ( signal_8176 ) ) ;
    buf_clk cell_2586 ( .C ( clk ), .D ( signal_8177 ), .Q ( signal_8178 ) ) ;
    buf_clk cell_2588 ( .C ( clk ), .D ( signal_8179 ), .Q ( signal_8180 ) ) ;
    buf_clk cell_2590 ( .C ( clk ), .D ( signal_8181 ), .Q ( signal_8182 ) ) ;
    buf_clk cell_2592 ( .C ( clk ), .D ( signal_8183 ), .Q ( signal_8184 ) ) ;
    buf_clk cell_2594 ( .C ( clk ), .D ( signal_8185 ), .Q ( signal_8186 ) ) ;
    buf_clk cell_2596 ( .C ( clk ), .D ( signal_8187 ), .Q ( signal_8188 ) ) ;
    buf_clk cell_2598 ( .C ( clk ), .D ( signal_8189 ), .Q ( signal_8190 ) ) ;
    buf_clk cell_2600 ( .C ( clk ), .D ( signal_8191 ), .Q ( signal_8192 ) ) ;
    buf_clk cell_2602 ( .C ( clk ), .D ( signal_8193 ), .Q ( signal_8194 ) ) ;
    buf_clk cell_2604 ( .C ( clk ), .D ( signal_8195 ), .Q ( signal_8196 ) ) ;
    buf_clk cell_2606 ( .C ( clk ), .D ( signal_8197 ), .Q ( signal_8198 ) ) ;
    buf_clk cell_2608 ( .C ( clk ), .D ( signal_8199 ), .Q ( signal_8200 ) ) ;
    buf_clk cell_2610 ( .C ( clk ), .D ( signal_8201 ), .Q ( signal_8202 ) ) ;
    buf_clk cell_2612 ( .C ( clk ), .D ( signal_8203 ), .Q ( signal_8204 ) ) ;
    buf_clk cell_2614 ( .C ( clk ), .D ( signal_8205 ), .Q ( signal_8206 ) ) ;
    buf_clk cell_2616 ( .C ( clk ), .D ( signal_8207 ), .Q ( signal_8208 ) ) ;
    buf_clk cell_2618 ( .C ( clk ), .D ( signal_8209 ), .Q ( signal_8210 ) ) ;
    buf_clk cell_2620 ( .C ( clk ), .D ( signal_8211 ), .Q ( signal_8212 ) ) ;
    buf_clk cell_2622 ( .C ( clk ), .D ( signal_8213 ), .Q ( signal_8214 ) ) ;
    buf_clk cell_2624 ( .C ( clk ), .D ( signal_8215 ), .Q ( signal_8216 ) ) ;
    buf_clk cell_2626 ( .C ( clk ), .D ( signal_8217 ), .Q ( signal_8218 ) ) ;
    buf_clk cell_2628 ( .C ( clk ), .D ( signal_8219 ), .Q ( signal_8220 ) ) ;
    buf_clk cell_2630 ( .C ( clk ), .D ( signal_8221 ), .Q ( signal_8222 ) ) ;
    buf_clk cell_2632 ( .C ( clk ), .D ( signal_8223 ), .Q ( signal_8224 ) ) ;
    buf_clk cell_2634 ( .C ( clk ), .D ( signal_8225 ), .Q ( signal_8226 ) ) ;
    buf_clk cell_2636 ( .C ( clk ), .D ( signal_8227 ), .Q ( signal_8228 ) ) ;
    buf_clk cell_2638 ( .C ( clk ), .D ( signal_8229 ), .Q ( signal_8230 ) ) ;
    buf_clk cell_2640 ( .C ( clk ), .D ( signal_8231 ), .Q ( signal_8232 ) ) ;
    buf_clk cell_2642 ( .C ( clk ), .D ( signal_8233 ), .Q ( signal_8234 ) ) ;
    buf_clk cell_2644 ( .C ( clk ), .D ( signal_8235 ), .Q ( signal_8236 ) ) ;
    buf_clk cell_2646 ( .C ( clk ), .D ( signal_8237 ), .Q ( signal_8238 ) ) ;
    buf_clk cell_2648 ( .C ( clk ), .D ( signal_8239 ), .Q ( signal_8240 ) ) ;
    buf_clk cell_2650 ( .C ( clk ), .D ( signal_8241 ), .Q ( signal_8242 ) ) ;
    buf_clk cell_2652 ( .C ( clk ), .D ( signal_8243 ), .Q ( signal_8244 ) ) ;
    buf_clk cell_2654 ( .C ( clk ), .D ( signal_8245 ), .Q ( signal_8246 ) ) ;
    buf_clk cell_2656 ( .C ( clk ), .D ( signal_8247 ), .Q ( signal_8248 ) ) ;
    buf_clk cell_2658 ( .C ( clk ), .D ( signal_8249 ), .Q ( signal_8250 ) ) ;
    buf_clk cell_2660 ( .C ( clk ), .D ( signal_8251 ), .Q ( signal_8252 ) ) ;
    buf_clk cell_2662 ( .C ( clk ), .D ( signal_8253 ), .Q ( signal_8254 ) ) ;
    buf_clk cell_2664 ( .C ( clk ), .D ( signal_8255 ), .Q ( signal_8256 ) ) ;
    buf_clk cell_2666 ( .C ( clk ), .D ( signal_8257 ), .Q ( signal_8258 ) ) ;
    buf_clk cell_2668 ( .C ( clk ), .D ( signal_8259 ), .Q ( signal_8260 ) ) ;
    buf_clk cell_2670 ( .C ( clk ), .D ( signal_8261 ), .Q ( signal_8262 ) ) ;
    buf_clk cell_2672 ( .C ( clk ), .D ( signal_8263 ), .Q ( signal_8264 ) ) ;
    buf_clk cell_2674 ( .C ( clk ), .D ( signal_8265 ), .Q ( signal_8266 ) ) ;
    buf_clk cell_2676 ( .C ( clk ), .D ( signal_8267 ), .Q ( signal_8268 ) ) ;
    buf_clk cell_2678 ( .C ( clk ), .D ( signal_8269 ), .Q ( signal_8270 ) ) ;
    buf_clk cell_2682 ( .C ( clk ), .D ( signal_8273 ), .Q ( signal_8274 ) ) ;
    buf_clk cell_2686 ( .C ( clk ), .D ( signal_8277 ), .Q ( signal_8278 ) ) ;
    buf_clk cell_2690 ( .C ( clk ), .D ( signal_8281 ), .Q ( signal_8282 ) ) ;
    buf_clk cell_2692 ( .C ( clk ), .D ( signal_8283 ), .Q ( signal_8284 ) ) ;
    buf_clk cell_2694 ( .C ( clk ), .D ( signal_8285 ), .Q ( signal_8286 ) ) ;
    buf_clk cell_2696 ( .C ( clk ), .D ( signal_8287 ), .Q ( signal_8288 ) ) ;
    buf_clk cell_2698 ( .C ( clk ), .D ( signal_8289 ), .Q ( signal_8290 ) ) ;
    buf_clk cell_2700 ( .C ( clk ), .D ( signal_8291 ), .Q ( signal_8292 ) ) ;
    buf_clk cell_2702 ( .C ( clk ), .D ( signal_8293 ), .Q ( signal_8294 ) ) ;
    buf_clk cell_2704 ( .C ( clk ), .D ( signal_8295 ), .Q ( signal_8296 ) ) ;
    buf_clk cell_2706 ( .C ( clk ), .D ( signal_8297 ), .Q ( signal_8298 ) ) ;
    buf_clk cell_2708 ( .C ( clk ), .D ( signal_8299 ), .Q ( signal_8300 ) ) ;
    buf_clk cell_2710 ( .C ( clk ), .D ( signal_8301 ), .Q ( signal_8302 ) ) ;
    buf_clk cell_2712 ( .C ( clk ), .D ( signal_8303 ), .Q ( signal_8304 ) ) ;
    buf_clk cell_2714 ( .C ( clk ), .D ( signal_8305 ), .Q ( signal_8306 ) ) ;
    buf_clk cell_2716 ( .C ( clk ), .D ( signal_8307 ), .Q ( signal_8308 ) ) ;
    buf_clk cell_2718 ( .C ( clk ), .D ( signal_8309 ), .Q ( signal_8310 ) ) ;
    buf_clk cell_2720 ( .C ( clk ), .D ( signal_8311 ), .Q ( signal_8312 ) ) ;
    buf_clk cell_2722 ( .C ( clk ), .D ( signal_8313 ), .Q ( signal_8314 ) ) ;
    buf_clk cell_2724 ( .C ( clk ), .D ( signal_8315 ), .Q ( signal_8316 ) ) ;
    buf_clk cell_2726 ( .C ( clk ), .D ( signal_8317 ), .Q ( signal_8318 ) ) ;
    buf_clk cell_2728 ( .C ( clk ), .D ( signal_8319 ), .Q ( signal_8320 ) ) ;
    buf_clk cell_2730 ( .C ( clk ), .D ( signal_8321 ), .Q ( signal_8322 ) ) ;
    buf_clk cell_2732 ( .C ( clk ), .D ( signal_8323 ), .Q ( signal_8324 ) ) ;
    buf_clk cell_2734 ( .C ( clk ), .D ( signal_8325 ), .Q ( signal_8326 ) ) ;
    buf_clk cell_2736 ( .C ( clk ), .D ( signal_8327 ), .Q ( signal_8328 ) ) ;
    buf_clk cell_2738 ( .C ( clk ), .D ( signal_8329 ), .Q ( signal_8330 ) ) ;
    buf_clk cell_2740 ( .C ( clk ), .D ( signal_8331 ), .Q ( signal_8332 ) ) ;
    buf_clk cell_2742 ( .C ( clk ), .D ( signal_8333 ), .Q ( signal_8334 ) ) ;
    buf_clk cell_2744 ( .C ( clk ), .D ( signal_8335 ), .Q ( signal_8336 ) ) ;
    buf_clk cell_2746 ( .C ( clk ), .D ( signal_8337 ), .Q ( signal_8338 ) ) ;
    buf_clk cell_2748 ( .C ( clk ), .D ( signal_8339 ), .Q ( signal_8340 ) ) ;
    buf_clk cell_2750 ( .C ( clk ), .D ( signal_8341 ), .Q ( signal_8342 ) ) ;
    buf_clk cell_2752 ( .C ( clk ), .D ( signal_8343 ), .Q ( signal_8344 ) ) ;
    buf_clk cell_2754 ( .C ( clk ), .D ( signal_8345 ), .Q ( signal_8346 ) ) ;
    buf_clk cell_2756 ( .C ( clk ), .D ( signal_8347 ), .Q ( signal_8348 ) ) ;
    buf_clk cell_2758 ( .C ( clk ), .D ( signal_8349 ), .Q ( signal_8350 ) ) ;
    buf_clk cell_2760 ( .C ( clk ), .D ( signal_8351 ), .Q ( signal_8352 ) ) ;
    buf_clk cell_2762 ( .C ( clk ), .D ( signal_8353 ), .Q ( signal_8354 ) ) ;
    buf_clk cell_2764 ( .C ( clk ), .D ( signal_8355 ), .Q ( signal_8356 ) ) ;
    buf_clk cell_2766 ( .C ( clk ), .D ( signal_8357 ), .Q ( signal_8358 ) ) ;
    buf_clk cell_2768 ( .C ( clk ), .D ( signal_8359 ), .Q ( signal_8360 ) ) ;
    buf_clk cell_2770 ( .C ( clk ), .D ( signal_8361 ), .Q ( signal_8362 ) ) ;
    buf_clk cell_2772 ( .C ( clk ), .D ( signal_8363 ), .Q ( signal_8364 ) ) ;
    buf_clk cell_2774 ( .C ( clk ), .D ( signal_8365 ), .Q ( signal_8366 ) ) ;
    buf_clk cell_2776 ( .C ( clk ), .D ( signal_8367 ), .Q ( signal_8368 ) ) ;
    buf_clk cell_2778 ( .C ( clk ), .D ( signal_8369 ), .Q ( signal_8370 ) ) ;
    buf_clk cell_2780 ( .C ( clk ), .D ( signal_8371 ), .Q ( signal_8372 ) ) ;
    buf_clk cell_2782 ( .C ( clk ), .D ( signal_8373 ), .Q ( signal_8374 ) ) ;
    buf_clk cell_2784 ( .C ( clk ), .D ( signal_8375 ), .Q ( signal_8376 ) ) ;
    buf_clk cell_2786 ( .C ( clk ), .D ( signal_8377 ), .Q ( signal_8378 ) ) ;
    buf_clk cell_2788 ( .C ( clk ), .D ( signal_8379 ), .Q ( signal_8380 ) ) ;
    buf_clk cell_2790 ( .C ( clk ), .D ( signal_8381 ), .Q ( signal_8382 ) ) ;
    buf_clk cell_2792 ( .C ( clk ), .D ( signal_8383 ), .Q ( signal_8384 ) ) ;
    buf_clk cell_2794 ( .C ( clk ), .D ( signal_8385 ), .Q ( signal_8386 ) ) ;
    buf_clk cell_2796 ( .C ( clk ), .D ( signal_8387 ), .Q ( signal_8388 ) ) ;
    buf_clk cell_2798 ( .C ( clk ), .D ( signal_8389 ), .Q ( signal_8390 ) ) ;
    buf_clk cell_2800 ( .C ( clk ), .D ( signal_8391 ), .Q ( signal_8392 ) ) ;
    buf_clk cell_2802 ( .C ( clk ), .D ( signal_8393 ), .Q ( signal_8394 ) ) ;
    buf_clk cell_2804 ( .C ( clk ), .D ( signal_8395 ), .Q ( signal_8396 ) ) ;
    buf_clk cell_2806 ( .C ( clk ), .D ( signal_8397 ), .Q ( signal_8398 ) ) ;
    buf_clk cell_2808 ( .C ( clk ), .D ( signal_8399 ), .Q ( signal_8400 ) ) ;
    buf_clk cell_2810 ( .C ( clk ), .D ( signal_8401 ), .Q ( signal_8402 ) ) ;
    buf_clk cell_2812 ( .C ( clk ), .D ( signal_8403 ), .Q ( signal_8404 ) ) ;
    buf_clk cell_2814 ( .C ( clk ), .D ( signal_8405 ), .Q ( signal_8406 ) ) ;
    buf_clk cell_2816 ( .C ( clk ), .D ( signal_8407 ), .Q ( signal_8408 ) ) ;
    buf_clk cell_2818 ( .C ( clk ), .D ( signal_8409 ), .Q ( signal_8410 ) ) ;
    buf_clk cell_2820 ( .C ( clk ), .D ( signal_8411 ), .Q ( signal_8412 ) ) ;
    buf_clk cell_2822 ( .C ( clk ), .D ( signal_8413 ), .Q ( signal_8414 ) ) ;
    buf_clk cell_2892 ( .C ( clk ), .D ( signal_8483 ), .Q ( signal_8484 ) ) ;
    buf_clk cell_2898 ( .C ( clk ), .D ( signal_8489 ), .Q ( signal_8490 ) ) ;
    buf_clk cell_2904 ( .C ( clk ), .D ( signal_8495 ), .Q ( signal_8496 ) ) ;
    buf_clk cell_3028 ( .C ( clk ), .D ( signal_8619 ), .Q ( signal_8620 ) ) ;
    buf_clk cell_3032 ( .C ( clk ), .D ( signal_8623 ), .Q ( signal_8624 ) ) ;
    buf_clk cell_3036 ( .C ( clk ), .D ( signal_8627 ), .Q ( signal_8628 ) ) ;
    buf_clk cell_3052 ( .C ( clk ), .D ( signal_8643 ), .Q ( signal_8644 ) ) ;
    buf_clk cell_3056 ( .C ( clk ), .D ( signal_8647 ), .Q ( signal_8648 ) ) ;
    buf_clk cell_3060 ( .C ( clk ), .D ( signal_8651 ), .Q ( signal_8652 ) ) ;
    buf_clk cell_3130 ( .C ( clk ), .D ( signal_8721 ), .Q ( signal_8722 ) ) ;
    buf_clk cell_3134 ( .C ( clk ), .D ( signal_8725 ), .Q ( signal_8726 ) ) ;
    buf_clk cell_3138 ( .C ( clk ), .D ( signal_8729 ), .Q ( signal_8730 ) ) ;
    buf_clk cell_3148 ( .C ( clk ), .D ( signal_8739 ), .Q ( signal_8740 ) ) ;
    buf_clk cell_3152 ( .C ( clk ), .D ( signal_8743 ), .Q ( signal_8744 ) ) ;
    buf_clk cell_3156 ( .C ( clk ), .D ( signal_8747 ), .Q ( signal_8748 ) ) ;
    buf_clk cell_3180 ( .C ( clk ), .D ( signal_8771 ), .Q ( signal_8772 ) ) ;
    buf_clk cell_3186 ( .C ( clk ), .D ( signal_8777 ), .Q ( signal_8778 ) ) ;
    buf_clk cell_3192 ( .C ( clk ), .D ( signal_8783 ), .Q ( signal_8784 ) ) ;
    buf_clk cell_3220 ( .C ( clk ), .D ( signal_8811 ), .Q ( signal_8812 ) ) ;
    buf_clk cell_3224 ( .C ( clk ), .D ( signal_8815 ), .Q ( signal_8816 ) ) ;
    buf_clk cell_3228 ( .C ( clk ), .D ( signal_8819 ), .Q ( signal_8820 ) ) ;
    buf_clk cell_3286 ( .C ( clk ), .D ( signal_8877 ), .Q ( signal_8878 ) ) ;
    buf_clk cell_3290 ( .C ( clk ), .D ( signal_8881 ), .Q ( signal_8882 ) ) ;
    buf_clk cell_3294 ( .C ( clk ), .D ( signal_8885 ), .Q ( signal_8886 ) ) ;
    buf_clk cell_3402 ( .C ( clk ), .D ( signal_8993 ), .Q ( signal_8994 ) ) ;
    buf_clk cell_3410 ( .C ( clk ), .D ( signal_9001 ), .Q ( signal_9002 ) ) ;
    buf_clk cell_3418 ( .C ( clk ), .D ( signal_9009 ), .Q ( signal_9010 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_2823 ( .C ( clk ), .D ( signal_1293 ), .Q ( signal_8415 ) ) ;
    buf_clk cell_2825 ( .C ( clk ), .D ( signal_3110 ), .Q ( signal_8417 ) ) ;
    buf_clk cell_2827 ( .C ( clk ), .D ( signal_3111 ), .Q ( signal_8419 ) ) ;
    buf_clk cell_2829 ( .C ( clk ), .D ( signal_8260 ), .Q ( signal_8421 ) ) ;
    buf_clk cell_2831 ( .C ( clk ), .D ( signal_8262 ), .Q ( signal_8423 ) ) ;
    buf_clk cell_2833 ( .C ( clk ), .D ( signal_8264 ), .Q ( signal_8425 ) ) ;
    buf_clk cell_2835 ( .C ( clk ), .D ( signal_1328 ), .Q ( signal_8427 ) ) ;
    buf_clk cell_2837 ( .C ( clk ), .D ( signal_3180 ), .Q ( signal_8429 ) ) ;
    buf_clk cell_2839 ( .C ( clk ), .D ( signal_3181 ), .Q ( signal_8431 ) ) ;
    buf_clk cell_2841 ( .C ( clk ), .D ( signal_1342 ), .Q ( signal_8433 ) ) ;
    buf_clk cell_2843 ( .C ( clk ), .D ( signal_3208 ), .Q ( signal_8435 ) ) ;
    buf_clk cell_2845 ( .C ( clk ), .D ( signal_3209 ), .Q ( signal_8437 ) ) ;
    buf_clk cell_2847 ( .C ( clk ), .D ( signal_1282 ), .Q ( signal_8439 ) ) ;
    buf_clk cell_2849 ( .C ( clk ), .D ( signal_3088 ), .Q ( signal_8441 ) ) ;
    buf_clk cell_2851 ( .C ( clk ), .D ( signal_3089 ), .Q ( signal_8443 ) ) ;
    buf_clk cell_2853 ( .C ( clk ), .D ( signal_1291 ), .Q ( signal_8445 ) ) ;
    buf_clk cell_2855 ( .C ( clk ), .D ( signal_3106 ), .Q ( signal_8447 ) ) ;
    buf_clk cell_2857 ( .C ( clk ), .D ( signal_3107 ), .Q ( signal_8449 ) ) ;
    buf_clk cell_2859 ( .C ( clk ), .D ( signal_8110 ), .Q ( signal_8451 ) ) ;
    buf_clk cell_2861 ( .C ( clk ), .D ( signal_8112 ), .Q ( signal_8453 ) ) ;
    buf_clk cell_2863 ( .C ( clk ), .D ( signal_8114 ), .Q ( signal_8455 ) ) ;
    buf_clk cell_2865 ( .C ( clk ), .D ( signal_8158 ), .Q ( signal_8457 ) ) ;
    buf_clk cell_2867 ( .C ( clk ), .D ( signal_8160 ), .Q ( signal_8459 ) ) ;
    buf_clk cell_2869 ( .C ( clk ), .D ( signal_8162 ), .Q ( signal_8461 ) ) ;
    buf_clk cell_2871 ( .C ( clk ), .D ( signal_8164 ), .Q ( signal_8463 ) ) ;
    buf_clk cell_2873 ( .C ( clk ), .D ( signal_8166 ), .Q ( signal_8465 ) ) ;
    buf_clk cell_2875 ( .C ( clk ), .D ( signal_8168 ), .Q ( signal_8467 ) ) ;
    buf_clk cell_2877 ( .C ( clk ), .D ( signal_8356 ), .Q ( signal_8469 ) ) ;
    buf_clk cell_2879 ( .C ( clk ), .D ( signal_8358 ), .Q ( signal_8471 ) ) ;
    buf_clk cell_2881 ( .C ( clk ), .D ( signal_8360 ), .Q ( signal_8473 ) ) ;
    buf_clk cell_2883 ( .C ( clk ), .D ( signal_8218 ), .Q ( signal_8475 ) ) ;
    buf_clk cell_2885 ( .C ( clk ), .D ( signal_8220 ), .Q ( signal_8477 ) ) ;
    buf_clk cell_2887 ( .C ( clk ), .D ( signal_8222 ), .Q ( signal_8479 ) ) ;
    buf_clk cell_2893 ( .C ( clk ), .D ( signal_8484 ), .Q ( signal_8485 ) ) ;
    buf_clk cell_2899 ( .C ( clk ), .D ( signal_8490 ), .Q ( signal_8491 ) ) ;
    buf_clk cell_2905 ( .C ( clk ), .D ( signal_8496 ), .Q ( signal_8497 ) ) ;
    buf_clk cell_2907 ( .C ( clk ), .D ( signal_8254 ), .Q ( signal_8499 ) ) ;
    buf_clk cell_2909 ( .C ( clk ), .D ( signal_8256 ), .Q ( signal_8501 ) ) ;
    buf_clk cell_2911 ( .C ( clk ), .D ( signal_8258 ), .Q ( signal_8503 ) ) ;
    buf_clk cell_2913 ( .C ( clk ), .D ( signal_8374 ), .Q ( signal_8505 ) ) ;
    buf_clk cell_2915 ( .C ( clk ), .D ( signal_8376 ), .Q ( signal_8507 ) ) ;
    buf_clk cell_2917 ( .C ( clk ), .D ( signal_8378 ), .Q ( signal_8509 ) ) ;
    buf_clk cell_2919 ( .C ( clk ), .D ( signal_8086 ), .Q ( signal_8511 ) ) ;
    buf_clk cell_2921 ( .C ( clk ), .D ( signal_8088 ), .Q ( signal_8513 ) ) ;
    buf_clk cell_2923 ( .C ( clk ), .D ( signal_8090 ), .Q ( signal_8515 ) ) ;
    buf_clk cell_2925 ( .C ( clk ), .D ( signal_8152 ), .Q ( signal_8517 ) ) ;
    buf_clk cell_2927 ( .C ( clk ), .D ( signal_8154 ), .Q ( signal_8519 ) ) ;
    buf_clk cell_2929 ( .C ( clk ), .D ( signal_8156 ), .Q ( signal_8521 ) ) ;
    buf_clk cell_2931 ( .C ( clk ), .D ( signal_1048 ), .Q ( signal_8523 ) ) ;
    buf_clk cell_2933 ( .C ( clk ), .D ( signal_2620 ), .Q ( signal_8525 ) ) ;
    buf_clk cell_2935 ( .C ( clk ), .D ( signal_2621 ), .Q ( signal_8527 ) ) ;
    buf_clk cell_2937 ( .C ( clk ), .D ( signal_8134 ), .Q ( signal_8529 ) ) ;
    buf_clk cell_2939 ( .C ( clk ), .D ( signal_8136 ), .Q ( signal_8531 ) ) ;
    buf_clk cell_2941 ( .C ( clk ), .D ( signal_8138 ), .Q ( signal_8533 ) ) ;
    buf_clk cell_2943 ( .C ( clk ), .D ( signal_1262 ), .Q ( signal_8535 ) ) ;
    buf_clk cell_2945 ( .C ( clk ), .D ( signal_3048 ), .Q ( signal_8537 ) ) ;
    buf_clk cell_2947 ( .C ( clk ), .D ( signal_3049 ), .Q ( signal_8539 ) ) ;
    buf_clk cell_2949 ( .C ( clk ), .D ( signal_1244 ), .Q ( signal_8541 ) ) ;
    buf_clk cell_2951 ( .C ( clk ), .D ( signal_3012 ), .Q ( signal_8543 ) ) ;
    buf_clk cell_2953 ( .C ( clk ), .D ( signal_3013 ), .Q ( signal_8545 ) ) ;
    buf_clk cell_2955 ( .C ( clk ), .D ( signal_1275 ), .Q ( signal_8547 ) ) ;
    buf_clk cell_2957 ( .C ( clk ), .D ( signal_3074 ), .Q ( signal_8549 ) ) ;
    buf_clk cell_2959 ( .C ( clk ), .D ( signal_3075 ), .Q ( signal_8551 ) ) ;
    buf_clk cell_2961 ( .C ( clk ), .D ( signal_1255 ), .Q ( signal_8553 ) ) ;
    buf_clk cell_2963 ( .C ( clk ), .D ( signal_3034 ), .Q ( signal_8555 ) ) ;
    buf_clk cell_2965 ( .C ( clk ), .D ( signal_3035 ), .Q ( signal_8557 ) ) ;
    buf_clk cell_2967 ( .C ( clk ), .D ( signal_1353 ), .Q ( signal_8559 ) ) ;
    buf_clk cell_2969 ( .C ( clk ), .D ( signal_3230 ), .Q ( signal_8561 ) ) ;
    buf_clk cell_2971 ( .C ( clk ), .D ( signal_3231 ), .Q ( signal_8563 ) ) ;
    buf_clk cell_2973 ( .C ( clk ), .D ( signal_1349 ), .Q ( signal_8565 ) ) ;
    buf_clk cell_2975 ( .C ( clk ), .D ( signal_3222 ), .Q ( signal_8567 ) ) ;
    buf_clk cell_2977 ( .C ( clk ), .D ( signal_3223 ), .Q ( signal_8569 ) ) ;
    buf_clk cell_2979 ( .C ( clk ), .D ( signal_1232 ), .Q ( signal_8571 ) ) ;
    buf_clk cell_2981 ( .C ( clk ), .D ( signal_2988 ), .Q ( signal_8573 ) ) ;
    buf_clk cell_2983 ( .C ( clk ), .D ( signal_2989 ), .Q ( signal_8575 ) ) ;
    buf_clk cell_2985 ( .C ( clk ), .D ( signal_1285 ), .Q ( signal_8577 ) ) ;
    buf_clk cell_2987 ( .C ( clk ), .D ( signal_3094 ), .Q ( signal_8579 ) ) ;
    buf_clk cell_2989 ( .C ( clk ), .D ( signal_3095 ), .Q ( signal_8581 ) ) ;
    buf_clk cell_2991 ( .C ( clk ), .D ( signal_1245 ), .Q ( signal_8583 ) ) ;
    buf_clk cell_2993 ( .C ( clk ), .D ( signal_3014 ), .Q ( signal_8585 ) ) ;
    buf_clk cell_2995 ( .C ( clk ), .D ( signal_3015 ), .Q ( signal_8587 ) ) ;
    buf_clk cell_2997 ( .C ( clk ), .D ( signal_1246 ), .Q ( signal_8589 ) ) ;
    buf_clk cell_2999 ( .C ( clk ), .D ( signal_3016 ), .Q ( signal_8591 ) ) ;
    buf_clk cell_3001 ( .C ( clk ), .D ( signal_3017 ), .Q ( signal_8593 ) ) ;
    buf_clk cell_3003 ( .C ( clk ), .D ( signal_1063 ), .Q ( signal_8595 ) ) ;
    buf_clk cell_3005 ( .C ( clk ), .D ( signal_2650 ), .Q ( signal_8597 ) ) ;
    buf_clk cell_3007 ( .C ( clk ), .D ( signal_2651 ), .Q ( signal_8599 ) ) ;
    buf_clk cell_3009 ( .C ( clk ), .D ( signal_1301 ), .Q ( signal_8601 ) ) ;
    buf_clk cell_3011 ( .C ( clk ), .D ( signal_3126 ), .Q ( signal_8603 ) ) ;
    buf_clk cell_3013 ( .C ( clk ), .D ( signal_3127 ), .Q ( signal_8605 ) ) ;
    buf_clk cell_3015 ( .C ( clk ), .D ( signal_1249 ), .Q ( signal_8607 ) ) ;
    buf_clk cell_3017 ( .C ( clk ), .D ( signal_3022 ), .Q ( signal_8609 ) ) ;
    buf_clk cell_3019 ( .C ( clk ), .D ( signal_3023 ), .Q ( signal_8611 ) ) ;
    buf_clk cell_3021 ( .C ( clk ), .D ( signal_1303 ), .Q ( signal_8613 ) ) ;
    buf_clk cell_3023 ( .C ( clk ), .D ( signal_3130 ), .Q ( signal_8615 ) ) ;
    buf_clk cell_3025 ( .C ( clk ), .D ( signal_3131 ), .Q ( signal_8617 ) ) ;
    buf_clk cell_3029 ( .C ( clk ), .D ( signal_8620 ), .Q ( signal_8621 ) ) ;
    buf_clk cell_3033 ( .C ( clk ), .D ( signal_8624 ), .Q ( signal_8625 ) ) ;
    buf_clk cell_3037 ( .C ( clk ), .D ( signal_8628 ), .Q ( signal_8629 ) ) ;
    buf_clk cell_3039 ( .C ( clk ), .D ( signal_1253 ), .Q ( signal_8631 ) ) ;
    buf_clk cell_3041 ( .C ( clk ), .D ( signal_3030 ), .Q ( signal_8633 ) ) ;
    buf_clk cell_3043 ( .C ( clk ), .D ( signal_3031 ), .Q ( signal_8635 ) ) ;
    buf_clk cell_3045 ( .C ( clk ), .D ( signal_1259 ), .Q ( signal_8637 ) ) ;
    buf_clk cell_3047 ( .C ( clk ), .D ( signal_3042 ), .Q ( signal_8639 ) ) ;
    buf_clk cell_3049 ( .C ( clk ), .D ( signal_3043 ), .Q ( signal_8641 ) ) ;
    buf_clk cell_3053 ( .C ( clk ), .D ( signal_8644 ), .Q ( signal_8645 ) ) ;
    buf_clk cell_3057 ( .C ( clk ), .D ( signal_8648 ), .Q ( signal_8649 ) ) ;
    buf_clk cell_3061 ( .C ( clk ), .D ( signal_8652 ), .Q ( signal_8653 ) ) ;
    buf_clk cell_3063 ( .C ( clk ), .D ( signal_1339 ), .Q ( signal_8655 ) ) ;
    buf_clk cell_3065 ( .C ( clk ), .D ( signal_3202 ), .Q ( signal_8657 ) ) ;
    buf_clk cell_3067 ( .C ( clk ), .D ( signal_3203 ), .Q ( signal_8659 ) ) ;
    buf_clk cell_3069 ( .C ( clk ), .D ( signal_8182 ), .Q ( signal_8661 ) ) ;
    buf_clk cell_3071 ( .C ( clk ), .D ( signal_8184 ), .Q ( signal_8663 ) ) ;
    buf_clk cell_3073 ( .C ( clk ), .D ( signal_8186 ), .Q ( signal_8665 ) ) ;
    buf_clk cell_3075 ( .C ( clk ), .D ( signal_1272 ), .Q ( signal_8667 ) ) ;
    buf_clk cell_3077 ( .C ( clk ), .D ( signal_3068 ), .Q ( signal_8669 ) ) ;
    buf_clk cell_3079 ( .C ( clk ), .D ( signal_3069 ), .Q ( signal_8671 ) ) ;
    buf_clk cell_3081 ( .C ( clk ), .D ( signal_1062 ), .Q ( signal_8673 ) ) ;
    buf_clk cell_3083 ( .C ( clk ), .D ( signal_2648 ), .Q ( signal_8675 ) ) ;
    buf_clk cell_3085 ( .C ( clk ), .D ( signal_2649 ), .Q ( signal_8677 ) ) ;
    buf_clk cell_3087 ( .C ( clk ), .D ( signal_1345 ), .Q ( signal_8679 ) ) ;
    buf_clk cell_3089 ( .C ( clk ), .D ( signal_3214 ), .Q ( signal_8681 ) ) ;
    buf_clk cell_3091 ( .C ( clk ), .D ( signal_3215 ), .Q ( signal_8683 ) ) ;
    buf_clk cell_3093 ( .C ( clk ), .D ( signal_1278 ), .Q ( signal_8685 ) ) ;
    buf_clk cell_3095 ( .C ( clk ), .D ( signal_3080 ), .Q ( signal_8687 ) ) ;
    buf_clk cell_3097 ( .C ( clk ), .D ( signal_3081 ), .Q ( signal_8689 ) ) ;
    buf_clk cell_3099 ( .C ( clk ), .D ( signal_1238 ), .Q ( signal_8691 ) ) ;
    buf_clk cell_3101 ( .C ( clk ), .D ( signal_3000 ), .Q ( signal_8693 ) ) ;
    buf_clk cell_3103 ( .C ( clk ), .D ( signal_3001 ), .Q ( signal_8695 ) ) ;
    buf_clk cell_3105 ( .C ( clk ), .D ( signal_1279 ), .Q ( signal_8697 ) ) ;
    buf_clk cell_3107 ( .C ( clk ), .D ( signal_3082 ), .Q ( signal_8699 ) ) ;
    buf_clk cell_3109 ( .C ( clk ), .D ( signal_3083 ), .Q ( signal_8701 ) ) ;
    buf_clk cell_3111 ( .C ( clk ), .D ( signal_1233 ), .Q ( signal_8703 ) ) ;
    buf_clk cell_3113 ( .C ( clk ), .D ( signal_2990 ), .Q ( signal_8705 ) ) ;
    buf_clk cell_3115 ( .C ( clk ), .D ( signal_2991 ), .Q ( signal_8707 ) ) ;
    buf_clk cell_3117 ( .C ( clk ), .D ( signal_1286 ), .Q ( signal_8709 ) ) ;
    buf_clk cell_3119 ( .C ( clk ), .D ( signal_3096 ), .Q ( signal_8711 ) ) ;
    buf_clk cell_3121 ( .C ( clk ), .D ( signal_3097 ), .Q ( signal_8713 ) ) ;
    buf_clk cell_3123 ( .C ( clk ), .D ( signal_1265 ), .Q ( signal_8715 ) ) ;
    buf_clk cell_3125 ( .C ( clk ), .D ( signal_3054 ), .Q ( signal_8717 ) ) ;
    buf_clk cell_3127 ( .C ( clk ), .D ( signal_3055 ), .Q ( signal_8719 ) ) ;
    buf_clk cell_3131 ( .C ( clk ), .D ( signal_8722 ), .Q ( signal_8723 ) ) ;
    buf_clk cell_3135 ( .C ( clk ), .D ( signal_8726 ), .Q ( signal_8727 ) ) ;
    buf_clk cell_3139 ( .C ( clk ), .D ( signal_8730 ), .Q ( signal_8731 ) ) ;
    buf_clk cell_3141 ( .C ( clk ), .D ( signal_8248 ), .Q ( signal_8733 ) ) ;
    buf_clk cell_3143 ( .C ( clk ), .D ( signal_8250 ), .Q ( signal_8735 ) ) ;
    buf_clk cell_3145 ( .C ( clk ), .D ( signal_8252 ), .Q ( signal_8737 ) ) ;
    buf_clk cell_3149 ( .C ( clk ), .D ( signal_8740 ), .Q ( signal_8741 ) ) ;
    buf_clk cell_3153 ( .C ( clk ), .D ( signal_8744 ), .Q ( signal_8745 ) ) ;
    buf_clk cell_3157 ( .C ( clk ), .D ( signal_8748 ), .Q ( signal_8749 ) ) ;
    buf_clk cell_3159 ( .C ( clk ), .D ( signal_1333 ), .Q ( signal_8751 ) ) ;
    buf_clk cell_3161 ( .C ( clk ), .D ( signal_3190 ), .Q ( signal_8753 ) ) ;
    buf_clk cell_3163 ( .C ( clk ), .D ( signal_3191 ), .Q ( signal_8755 ) ) ;
    buf_clk cell_3165 ( .C ( clk ), .D ( signal_8296 ), .Q ( signal_8757 ) ) ;
    buf_clk cell_3167 ( .C ( clk ), .D ( signal_8298 ), .Q ( signal_8759 ) ) ;
    buf_clk cell_3169 ( .C ( clk ), .D ( signal_8300 ), .Q ( signal_8761 ) ) ;
    buf_clk cell_3171 ( .C ( clk ), .D ( signal_8274 ), .Q ( signal_8763 ) ) ;
    buf_clk cell_3173 ( .C ( clk ), .D ( signal_8278 ), .Q ( signal_8765 ) ) ;
    buf_clk cell_3175 ( .C ( clk ), .D ( signal_8282 ), .Q ( signal_8767 ) ) ;
    buf_clk cell_3181 ( .C ( clk ), .D ( signal_8772 ), .Q ( signal_8773 ) ) ;
    buf_clk cell_3187 ( .C ( clk ), .D ( signal_8778 ), .Q ( signal_8779 ) ) ;
    buf_clk cell_3193 ( .C ( clk ), .D ( signal_8784 ), .Q ( signal_8785 ) ) ;
    buf_clk cell_3195 ( .C ( clk ), .D ( signal_8224 ), .Q ( signal_8787 ) ) ;
    buf_clk cell_3197 ( .C ( clk ), .D ( signal_8226 ), .Q ( signal_8789 ) ) ;
    buf_clk cell_3199 ( .C ( clk ), .D ( signal_8228 ), .Q ( signal_8791 ) ) ;
    buf_clk cell_3201 ( .C ( clk ), .D ( signal_8098 ), .Q ( signal_8793 ) ) ;
    buf_clk cell_3203 ( .C ( clk ), .D ( signal_8100 ), .Q ( signal_8795 ) ) ;
    buf_clk cell_3205 ( .C ( clk ), .D ( signal_8102 ), .Q ( signal_8797 ) ) ;
    buf_clk cell_3207 ( .C ( clk ), .D ( signal_8302 ), .Q ( signal_8799 ) ) ;
    buf_clk cell_3209 ( .C ( clk ), .D ( signal_8304 ), .Q ( signal_8801 ) ) ;
    buf_clk cell_3211 ( .C ( clk ), .D ( signal_8306 ), .Q ( signal_8803 ) ) ;
    buf_clk cell_3213 ( .C ( clk ), .D ( signal_1145 ), .Q ( signal_8805 ) ) ;
    buf_clk cell_3215 ( .C ( clk ), .D ( signal_2814 ), .Q ( signal_8807 ) ) ;
    buf_clk cell_3217 ( .C ( clk ), .D ( signal_2815 ), .Q ( signal_8809 ) ) ;
    buf_clk cell_3221 ( .C ( clk ), .D ( signal_8812 ), .Q ( signal_8813 ) ) ;
    buf_clk cell_3225 ( .C ( clk ), .D ( signal_8816 ), .Q ( signal_8817 ) ) ;
    buf_clk cell_3229 ( .C ( clk ), .D ( signal_8820 ), .Q ( signal_8821 ) ) ;
    buf_clk cell_3231 ( .C ( clk ), .D ( signal_1095 ), .Q ( signal_8823 ) ) ;
    buf_clk cell_3233 ( .C ( clk ), .D ( signal_2714 ), .Q ( signal_8825 ) ) ;
    buf_clk cell_3235 ( .C ( clk ), .D ( signal_2715 ), .Q ( signal_8827 ) ) ;
    buf_clk cell_3237 ( .C ( clk ), .D ( signal_1078 ), .Q ( signal_8829 ) ) ;
    buf_clk cell_3239 ( .C ( clk ), .D ( signal_2680 ), .Q ( signal_8831 ) ) ;
    buf_clk cell_3241 ( .C ( clk ), .D ( signal_2681 ), .Q ( signal_8833 ) ) ;
    buf_clk cell_3243 ( .C ( clk ), .D ( signal_1073 ), .Q ( signal_8835 ) ) ;
    buf_clk cell_3245 ( .C ( clk ), .D ( signal_2670 ), .Q ( signal_8837 ) ) ;
    buf_clk cell_3247 ( .C ( clk ), .D ( signal_2671 ), .Q ( signal_8839 ) ) ;
    buf_clk cell_3249 ( .C ( clk ), .D ( signal_1158 ), .Q ( signal_8841 ) ) ;
    buf_clk cell_3251 ( .C ( clk ), .D ( signal_2840 ), .Q ( signal_8843 ) ) ;
    buf_clk cell_3253 ( .C ( clk ), .D ( signal_2841 ), .Q ( signal_8845 ) ) ;
    buf_clk cell_3255 ( .C ( clk ), .D ( signal_1020 ), .Q ( signal_8847 ) ) ;
    buf_clk cell_3257 ( .C ( clk ), .D ( signal_2564 ), .Q ( signal_8849 ) ) ;
    buf_clk cell_3259 ( .C ( clk ), .D ( signal_2565 ), .Q ( signal_8851 ) ) ;
    buf_clk cell_3261 ( .C ( clk ), .D ( signal_8380 ), .Q ( signal_8853 ) ) ;
    buf_clk cell_3263 ( .C ( clk ), .D ( signal_8382 ), .Q ( signal_8855 ) ) ;
    buf_clk cell_3265 ( .C ( clk ), .D ( signal_8384 ), .Q ( signal_8857 ) ) ;
    buf_clk cell_3267 ( .C ( clk ), .D ( signal_8266 ), .Q ( signal_8859 ) ) ;
    buf_clk cell_3269 ( .C ( clk ), .D ( signal_8268 ), .Q ( signal_8861 ) ) ;
    buf_clk cell_3271 ( .C ( clk ), .D ( signal_8270 ), .Q ( signal_8863 ) ) ;
    buf_clk cell_3273 ( .C ( clk ), .D ( signal_1162 ), .Q ( signal_8865 ) ) ;
    buf_clk cell_3275 ( .C ( clk ), .D ( signal_2848 ), .Q ( signal_8867 ) ) ;
    buf_clk cell_3277 ( .C ( clk ), .D ( signal_2849 ), .Q ( signal_8869 ) ) ;
    buf_clk cell_3279 ( .C ( clk ), .D ( signal_1071 ), .Q ( signal_8871 ) ) ;
    buf_clk cell_3281 ( .C ( clk ), .D ( signal_2666 ), .Q ( signal_8873 ) ) ;
    buf_clk cell_3283 ( .C ( clk ), .D ( signal_2667 ), .Q ( signal_8875 ) ) ;
    buf_clk cell_3287 ( .C ( clk ), .D ( signal_8878 ), .Q ( signal_8879 ) ) ;
    buf_clk cell_3291 ( .C ( clk ), .D ( signal_8882 ), .Q ( signal_8883 ) ) ;
    buf_clk cell_3295 ( .C ( clk ), .D ( signal_8886 ), .Q ( signal_8887 ) ) ;
    buf_clk cell_3297 ( .C ( clk ), .D ( signal_1081 ), .Q ( signal_8889 ) ) ;
    buf_clk cell_3299 ( .C ( clk ), .D ( signal_2686 ), .Q ( signal_8891 ) ) ;
    buf_clk cell_3301 ( .C ( clk ), .D ( signal_2687 ), .Q ( signal_8893 ) ) ;
    buf_clk cell_3303 ( .C ( clk ), .D ( signal_8338 ), .Q ( signal_8895 ) ) ;
    buf_clk cell_3305 ( .C ( clk ), .D ( signal_8340 ), .Q ( signal_8897 ) ) ;
    buf_clk cell_3307 ( .C ( clk ), .D ( signal_8342 ), .Q ( signal_8899 ) ) ;
    buf_clk cell_3309 ( .C ( clk ), .D ( signal_8308 ), .Q ( signal_8901 ) ) ;
    buf_clk cell_3311 ( .C ( clk ), .D ( signal_8310 ), .Q ( signal_8903 ) ) ;
    buf_clk cell_3313 ( .C ( clk ), .D ( signal_8312 ), .Q ( signal_8905 ) ) ;
    buf_clk cell_3315 ( .C ( clk ), .D ( signal_1304 ), .Q ( signal_8907 ) ) ;
    buf_clk cell_3317 ( .C ( clk ), .D ( signal_3132 ), .Q ( signal_8909 ) ) ;
    buf_clk cell_3319 ( .C ( clk ), .D ( signal_3133 ), .Q ( signal_8911 ) ) ;
    buf_clk cell_3321 ( .C ( clk ), .D ( signal_1250 ), .Q ( signal_8913 ) ) ;
    buf_clk cell_3323 ( .C ( clk ), .D ( signal_3024 ), .Q ( signal_8915 ) ) ;
    buf_clk cell_3325 ( .C ( clk ), .D ( signal_3025 ), .Q ( signal_8917 ) ) ;
    buf_clk cell_3327 ( .C ( clk ), .D ( signal_1327 ), .Q ( signal_8919 ) ) ;
    buf_clk cell_3329 ( .C ( clk ), .D ( signal_3178 ), .Q ( signal_8921 ) ) ;
    buf_clk cell_3331 ( .C ( clk ), .D ( signal_3179 ), .Q ( signal_8923 ) ) ;
    buf_clk cell_3345 ( .C ( clk ), .D ( signal_8404 ), .Q ( signal_8937 ) ) ;
    buf_clk cell_3349 ( .C ( clk ), .D ( signal_8406 ), .Q ( signal_8941 ) ) ;
    buf_clk cell_3353 ( .C ( clk ), .D ( signal_8408 ), .Q ( signal_8945 ) ) ;
    buf_clk cell_3363 ( .C ( clk ), .D ( signal_1290 ), .Q ( signal_8955 ) ) ;
    buf_clk cell_3367 ( .C ( clk ), .D ( signal_3104 ), .Q ( signal_8959 ) ) ;
    buf_clk cell_3371 ( .C ( clk ), .D ( signal_3105 ), .Q ( signal_8963 ) ) ;
    buf_clk cell_3375 ( .C ( clk ), .D ( signal_1354 ), .Q ( signal_8967 ) ) ;
    buf_clk cell_3379 ( .C ( clk ), .D ( signal_3232 ), .Q ( signal_8971 ) ) ;
    buf_clk cell_3383 ( .C ( clk ), .D ( signal_3233 ), .Q ( signal_8975 ) ) ;
    buf_clk cell_3387 ( .C ( clk ), .D ( signal_1234 ), .Q ( signal_8979 ) ) ;
    buf_clk cell_3391 ( .C ( clk ), .D ( signal_2992 ), .Q ( signal_8983 ) ) ;
    buf_clk cell_3395 ( .C ( clk ), .D ( signal_2993 ), .Q ( signal_8987 ) ) ;
    buf_clk cell_3403 ( .C ( clk ), .D ( signal_8994 ), .Q ( signal_8995 ) ) ;
    buf_clk cell_3411 ( .C ( clk ), .D ( signal_9002 ), .Q ( signal_9003 ) ) ;
    buf_clk cell_3419 ( .C ( clk ), .D ( signal_9010 ), .Q ( signal_9011 ) ) ;
    buf_clk cell_3435 ( .C ( clk ), .D ( signal_1313 ), .Q ( signal_9027 ) ) ;
    buf_clk cell_3439 ( .C ( clk ), .D ( signal_3150 ), .Q ( signal_9031 ) ) ;
    buf_clk cell_3443 ( .C ( clk ), .D ( signal_3151 ), .Q ( signal_9035 ) ) ;
    buf_clk cell_3459 ( .C ( clk ), .D ( signal_1335 ), .Q ( signal_9051 ) ) ;
    buf_clk cell_3463 ( .C ( clk ), .D ( signal_3194 ), .Q ( signal_9055 ) ) ;
    buf_clk cell_3467 ( .C ( clk ), .D ( signal_3195 ), .Q ( signal_9059 ) ) ;
    buf_clk cell_3501 ( .C ( clk ), .D ( signal_1061 ), .Q ( signal_9093 ) ) ;
    buf_clk cell_3505 ( .C ( clk ), .D ( signal_2646 ), .Q ( signal_9097 ) ) ;
    buf_clk cell_3509 ( .C ( clk ), .D ( signal_2647 ), .Q ( signal_9101 ) ) ;
    buf_clk cell_3537 ( .C ( clk ), .D ( signal_1361 ), .Q ( signal_9129 ) ) ;
    buf_clk cell_3541 ( .C ( clk ), .D ( signal_3246 ), .Q ( signal_9133 ) ) ;
    buf_clk cell_3545 ( .C ( clk ), .D ( signal_3247 ), .Q ( signal_9137 ) ) ;
    buf_clk cell_3561 ( .C ( clk ), .D ( signal_8146 ), .Q ( signal_9153 ) ) ;
    buf_clk cell_3565 ( .C ( clk ), .D ( signal_8148 ), .Q ( signal_9157 ) ) ;
    buf_clk cell_3569 ( .C ( clk ), .D ( signal_8150 ), .Q ( signal_9161 ) ) ;
    buf_clk cell_3573 ( .C ( clk ), .D ( signal_8176 ), .Q ( signal_9165 ) ) ;
    buf_clk cell_3577 ( .C ( clk ), .D ( signal_8178 ), .Q ( signal_9169 ) ) ;
    buf_clk cell_3581 ( .C ( clk ), .D ( signal_8180 ), .Q ( signal_9173 ) ) ;
    buf_clk cell_3585 ( .C ( clk ), .D ( signal_8284 ), .Q ( signal_9177 ) ) ;
    buf_clk cell_3589 ( .C ( clk ), .D ( signal_8286 ), .Q ( signal_9181 ) ) ;
    buf_clk cell_3593 ( .C ( clk ), .D ( signal_8288 ), .Q ( signal_9185 ) ) ;
    buf_clk cell_3597 ( .C ( clk ), .D ( signal_8104 ), .Q ( signal_9189 ) ) ;
    buf_clk cell_3601 ( .C ( clk ), .D ( signal_8106 ), .Q ( signal_9193 ) ) ;
    buf_clk cell_3605 ( .C ( clk ), .D ( signal_8108 ), .Q ( signal_9197 ) ) ;
    buf_clk cell_3639 ( .C ( clk ), .D ( signal_8122 ), .Q ( signal_9231 ) ) ;
    buf_clk cell_3643 ( .C ( clk ), .D ( signal_8124 ), .Q ( signal_9235 ) ) ;
    buf_clk cell_3647 ( .C ( clk ), .D ( signal_8126 ), .Q ( signal_9239 ) ) ;
    buf_clk cell_3651 ( .C ( clk ), .D ( signal_8116 ), .Q ( signal_9243 ) ) ;
    buf_clk cell_3655 ( .C ( clk ), .D ( signal_8118 ), .Q ( signal_9247 ) ) ;
    buf_clk cell_3659 ( .C ( clk ), .D ( signal_8120 ), .Q ( signal_9251 ) ) ;
    buf_clk cell_3663 ( .C ( clk ), .D ( signal_8230 ), .Q ( signal_9255 ) ) ;
    buf_clk cell_3667 ( .C ( clk ), .D ( signal_8232 ), .Q ( signal_9259 ) ) ;
    buf_clk cell_3671 ( .C ( clk ), .D ( signal_8234 ), .Q ( signal_9263 ) ) ;
    buf_clk cell_3681 ( .C ( clk ), .D ( signal_8170 ), .Q ( signal_9273 ) ) ;
    buf_clk cell_3685 ( .C ( clk ), .D ( signal_8172 ), .Q ( signal_9277 ) ) ;
    buf_clk cell_3689 ( .C ( clk ), .D ( signal_8174 ), .Q ( signal_9281 ) ) ;
    buf_clk cell_3723 ( .C ( clk ), .D ( signal_1080 ), .Q ( signal_9315 ) ) ;
    buf_clk cell_3727 ( .C ( clk ), .D ( signal_2684 ), .Q ( signal_9319 ) ) ;
    buf_clk cell_3731 ( .C ( clk ), .D ( signal_2685 ), .Q ( signal_9323 ) ) ;
    buf_clk cell_3735 ( .C ( clk ), .D ( signal_1365 ), .Q ( signal_9327 ) ) ;
    buf_clk cell_3739 ( .C ( clk ), .D ( signal_3254 ), .Q ( signal_9331 ) ) ;
    buf_clk cell_3743 ( .C ( clk ), .D ( signal_3255 ), .Q ( signal_9335 ) ) ;
    buf_clk cell_3753 ( .C ( clk ), .D ( signal_1242 ), .Q ( signal_9345 ) ) ;
    buf_clk cell_3757 ( .C ( clk ), .D ( signal_3008 ), .Q ( signal_9349 ) ) ;
    buf_clk cell_3761 ( .C ( clk ), .D ( signal_3009 ), .Q ( signal_9353 ) ) ;
    buf_clk cell_3777 ( .C ( clk ), .D ( signal_1296 ), .Q ( signal_9369 ) ) ;
    buf_clk cell_3781 ( .C ( clk ), .D ( signal_3116 ), .Q ( signal_9373 ) ) ;
    buf_clk cell_3785 ( .C ( clk ), .D ( signal_3117 ), .Q ( signal_9377 ) ) ;
    buf_clk cell_3789 ( .C ( clk ), .D ( signal_1308 ), .Q ( signal_9381 ) ) ;
    buf_clk cell_3793 ( .C ( clk ), .D ( signal_3140 ), .Q ( signal_9385 ) ) ;
    buf_clk cell_3797 ( .C ( clk ), .D ( signal_3141 ), .Q ( signal_9389 ) ) ;
    buf_clk cell_3801 ( .C ( clk ), .D ( signal_1251 ), .Q ( signal_9393 ) ) ;
    buf_clk cell_3805 ( .C ( clk ), .D ( signal_3026 ), .Q ( signal_9397 ) ) ;
    buf_clk cell_3809 ( .C ( clk ), .D ( signal_3027 ), .Q ( signal_9401 ) ) ;
    buf_clk cell_3819 ( .C ( clk ), .D ( signal_1326 ), .Q ( signal_9411 ) ) ;
    buf_clk cell_3823 ( .C ( clk ), .D ( signal_3176 ), .Q ( signal_9415 ) ) ;
    buf_clk cell_3827 ( .C ( clk ), .D ( signal_3177 ), .Q ( signal_9419 ) ) ;
    buf_clk cell_3831 ( .C ( clk ), .D ( signal_1261 ), .Q ( signal_9423 ) ) ;
    buf_clk cell_3835 ( .C ( clk ), .D ( signal_3046 ), .Q ( signal_9427 ) ) ;
    buf_clk cell_3839 ( .C ( clk ), .D ( signal_3047 ), .Q ( signal_9431 ) ) ;
    buf_clk cell_3849 ( .C ( clk ), .D ( signal_1271 ), .Q ( signal_9441 ) ) ;
    buf_clk cell_3853 ( .C ( clk ), .D ( signal_3066 ), .Q ( signal_9445 ) ) ;
    buf_clk cell_3857 ( .C ( clk ), .D ( signal_3067 ), .Q ( signal_9449 ) ) ;
    buf_clk cell_3879 ( .C ( clk ), .D ( signal_8092 ), .Q ( signal_9471 ) ) ;
    buf_clk cell_3883 ( .C ( clk ), .D ( signal_8094 ), .Q ( signal_9475 ) ) ;
    buf_clk cell_3887 ( .C ( clk ), .D ( signal_8096 ), .Q ( signal_9479 ) ) ;
    buf_clk cell_3897 ( .C ( clk ), .D ( signal_8410 ), .Q ( signal_9489 ) ) ;
    buf_clk cell_3903 ( .C ( clk ), .D ( signal_8412 ), .Q ( signal_9495 ) ) ;
    buf_clk cell_3909 ( .C ( clk ), .D ( signal_8414 ), .Q ( signal_9501 ) ) ;
    buf_clk cell_3915 ( .C ( clk ), .D ( signal_1248 ), .Q ( signal_9507 ) ) ;
    buf_clk cell_3921 ( .C ( clk ), .D ( signal_3020 ), .Q ( signal_9513 ) ) ;
    buf_clk cell_3927 ( .C ( clk ), .D ( signal_3021 ), .Q ( signal_9519 ) ) ;
    buf_clk cell_3933 ( .C ( clk ), .D ( signal_1314 ), .Q ( signal_9525 ) ) ;
    buf_clk cell_3939 ( .C ( clk ), .D ( signal_3152 ), .Q ( signal_9531 ) ) ;
    buf_clk cell_3945 ( .C ( clk ), .D ( signal_3153 ), .Q ( signal_9537 ) ) ;
    buf_clk cell_3963 ( .C ( clk ), .D ( signal_1336 ), .Q ( signal_9555 ) ) ;
    buf_clk cell_3969 ( .C ( clk ), .D ( signal_3196 ), .Q ( signal_9561 ) ) ;
    buf_clk cell_3975 ( .C ( clk ), .D ( signal_3197 ), .Q ( signal_9567 ) ) ;
    buf_clk cell_4041 ( .C ( clk ), .D ( signal_8236 ), .Q ( signal_9633 ) ) ;
    buf_clk cell_4047 ( .C ( clk ), .D ( signal_8238 ), .Q ( signal_9639 ) ) ;
    buf_clk cell_4053 ( .C ( clk ), .D ( signal_8240 ), .Q ( signal_9645 ) ) ;
    buf_clk cell_4131 ( .C ( clk ), .D ( signal_8074 ), .Q ( signal_9723 ) ) ;
    buf_clk cell_4137 ( .C ( clk ), .D ( signal_8076 ), .Q ( signal_9729 ) ) ;
    buf_clk cell_4143 ( .C ( clk ), .D ( signal_8078 ), .Q ( signal_9735 ) ) ;
    buf_clk cell_4179 ( .C ( clk ), .D ( signal_1298 ), .Q ( signal_9771 ) ) ;
    buf_clk cell_4185 ( .C ( clk ), .D ( signal_3120 ), .Q ( signal_9777 ) ) ;
    buf_clk cell_4191 ( .C ( clk ), .D ( signal_3121 ), .Q ( signal_9783 ) ) ;
    buf_clk cell_4263 ( .C ( clk ), .D ( signal_1064 ), .Q ( signal_9855 ) ) ;
    buf_clk cell_4269 ( .C ( clk ), .D ( signal_2652 ), .Q ( signal_9861 ) ) ;
    buf_clk cell_4275 ( .C ( clk ), .D ( signal_2653 ), .Q ( signal_9867 ) ) ;
    buf_clk cell_4293 ( .C ( clk ), .D ( signal_1316 ), .Q ( signal_9885 ) ) ;
    buf_clk cell_4299 ( .C ( clk ), .D ( signal_3156 ), .Q ( signal_9891 ) ) ;
    buf_clk cell_4305 ( .C ( clk ), .D ( signal_3157 ), .Q ( signal_9897 ) ) ;
    buf_clk cell_4377 ( .C ( clk ), .D ( signal_1289 ), .Q ( signal_9969 ) ) ;
    buf_clk cell_4383 ( .C ( clk ), .D ( signal_3102 ), .Q ( signal_9975 ) ) ;
    buf_clk cell_4389 ( .C ( clk ), .D ( signal_3103 ), .Q ( signal_9981 ) ) ;
    buf_clk cell_4419 ( .C ( clk ), .D ( signal_1359 ), .Q ( signal_10011 ) ) ;
    buf_clk cell_4425 ( .C ( clk ), .D ( signal_3242 ), .Q ( signal_10017 ) ) ;
    buf_clk cell_4431 ( .C ( clk ), .D ( signal_3243 ), .Q ( signal_10023 ) ) ;
    buf_clk cell_4437 ( .C ( clk ), .D ( signal_1307 ), .Q ( signal_10029 ) ) ;
    buf_clk cell_4443 ( .C ( clk ), .D ( signal_3138 ), .Q ( signal_10035 ) ) ;
    buf_clk cell_4449 ( .C ( clk ), .D ( signal_3139 ), .Q ( signal_10041 ) ) ;
    buf_clk cell_4455 ( .C ( clk ), .D ( signal_8290 ), .Q ( signal_10047 ) ) ;
    buf_clk cell_4461 ( .C ( clk ), .D ( signal_8292 ), .Q ( signal_10053 ) ) ;
    buf_clk cell_4467 ( .C ( clk ), .D ( signal_8294 ), .Q ( signal_10059 ) ) ;
    buf_clk cell_4497 ( .C ( clk ), .D ( signal_1315 ), .Q ( signal_10089 ) ) ;
    buf_clk cell_4505 ( .C ( clk ), .D ( signal_3154 ), .Q ( signal_10097 ) ) ;
    buf_clk cell_4513 ( .C ( clk ), .D ( signal_3155 ), .Q ( signal_10105 ) ) ;
    buf_clk cell_4755 ( .C ( clk ), .D ( signal_1239 ), .Q ( signal_10347 ) ) ;
    buf_clk cell_4763 ( .C ( clk ), .D ( signal_3002 ), .Q ( signal_10355 ) ) ;
    buf_clk cell_4771 ( .C ( clk ), .D ( signal_3003 ), .Q ( signal_10363 ) ) ;
    buf_clk cell_4851 ( .C ( clk ), .D ( signal_1060 ), .Q ( signal_10443 ) ) ;
    buf_clk cell_4859 ( .C ( clk ), .D ( signal_2644 ), .Q ( signal_10451 ) ) ;
    buf_clk cell_4867 ( .C ( clk ), .D ( signal_2645 ), .Q ( signal_10459 ) ) ;
    buf_clk cell_5001 ( .C ( clk ), .D ( signal_1254 ), .Q ( signal_10593 ) ) ;
    buf_clk cell_5011 ( .C ( clk ), .D ( signal_3032 ), .Q ( signal_10603 ) ) ;
    buf_clk cell_5021 ( .C ( clk ), .D ( signal_3033 ), .Q ( signal_10613 ) ) ;
    buf_clk cell_5145 ( .C ( clk ), .D ( signal_1247 ), .Q ( signal_10737 ) ) ;
    buf_clk cell_5155 ( .C ( clk ), .D ( signal_3018 ), .Q ( signal_10747 ) ) ;
    buf_clk cell_5165 ( .C ( clk ), .D ( signal_3019 ), .Q ( signal_10757 ) ) ;
    buf_clk cell_5313 ( .C ( clk ), .D ( signal_1066 ), .Q ( signal_10905 ) ) ;
    buf_clk cell_5323 ( .C ( clk ), .D ( signal_2656 ), .Q ( signal_10915 ) ) ;
    buf_clk cell_5333 ( .C ( clk ), .D ( signal_2657 ), .Q ( signal_10925 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1085 ( .a ({signal_8066, signal_8062, signal_8058}), .b ({signal_2553, signal_2552, signal_1014}), .clk ( clk ), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_2725, signal_2724, signal_1100}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1124 ( .a ({signal_8072, signal_8070, signal_8068}), .b ({signal_2563, signal_2562, signal_1019}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({signal_2803, signal_2802, signal_1139}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1132 ( .a ({signal_8078, signal_8076, signal_8074}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_2819, signal_2818, signal_1147}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1140 ( .a ({signal_8084, signal_8082, signal_8080}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({signal_2835, signal_2834, signal_1155}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1155 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_2565, signal_2564, signal_1020}), .clk ( clk ), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_2865, signal_2864, signal_1170}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1173 ( .a ({signal_8096, signal_8094, signal_8092}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({signal_2901, signal_2900, signal_1188}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1184 ( .a ({signal_8102, signal_8100, signal_8098}), .b ({signal_2573, signal_2572, signal_1024}), .clk ( clk ), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_2923, signal_2922, signal_1199}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1189 ( .a ({signal_8108, signal_8106, signal_8104}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({signal_2933, signal_2932, signal_1204}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1190 ( .a ({signal_8114, signal_8112, signal_8110}), .b ({signal_2573, signal_2572, signal_1024}), .clk ( clk ), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_2935, signal_2934, signal_1205}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1198 ( .a ({signal_8120, signal_8118, signal_8116}), .b ({signal_2573, signal_2572, signal_1024}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({signal_2951, signal_2950, signal_1213}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1207 ( .a ({signal_8126, signal_8124, signal_8122}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_2969, signal_2968, signal_1222}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1209 ( .a ({signal_8132, signal_8130, signal_8128}), .b ({signal_2577, signal_2576, signal_1026}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({signal_2973, signal_2972, signal_1224}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1211 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2565, signal_2564, signal_1020}), .clk ( clk ), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_2977, signal_2976, signal_1226}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1212 ( .a ({signal_8144, signal_8142, signal_8140}), .b ({signal_2565, signal_2564, signal_1020}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({signal_2979, signal_2978, signal_1227}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1243 ( .a ({signal_2725, signal_2724, signal_1100}), .b ({signal_3041, signal_3040, signal_1258}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1272 ( .a ({signal_2803, signal_2802, signal_1139}), .b ({signal_3099, signal_3098, signal_1287}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1277 ( .a ({signal_2819, signal_2818, signal_1147}), .b ({signal_3109, signal_3108, signal_1292}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1284 ( .a ({signal_2835, signal_2834, signal_1155}), .b ({signal_3123, signal_3122, signal_1299}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1297 ( .a ({signal_2865, signal_2864, signal_1170}), .b ({signal_3149, signal_3148, signal_1312}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1314 ( .a ({signal_2901, signal_2900, signal_1188}), .b ({signal_3183, signal_3182, signal_1329}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1323 ( .a ({signal_2923, signal_2922, signal_1199}), .b ({signal_3201, signal_3200, signal_1338}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1328 ( .a ({signal_2933, signal_2932, signal_1204}), .b ({signal_3211, signal_3210, signal_1343}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1329 ( .a ({signal_2935, signal_2934, signal_1205}), .b ({signal_3213, signal_3212, signal_1344}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1335 ( .a ({signal_2951, signal_2950, signal_1213}), .b ({signal_3225, signal_3224, signal_1350}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1343 ( .a ({signal_2969, signal_2968, signal_1222}), .b ({signal_3241, signal_3240, signal_1358}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1345 ( .a ({signal_2973, signal_2972, signal_1224}), .b ({signal_3245, signal_3244, signal_1360}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1347 ( .a ({signal_2977, signal_2976, signal_1226}), .b ({signal_3249, signal_3248, signal_1362}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1348 ( .a ({signal_2979, signal_2978, signal_1227}), .b ({signal_3251, signal_3250, signal_1363}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1351 ( .a ({signal_8150, signal_8148, signal_8146}), .b ({signal_2659, signal_2658, signal_1067}), .clk ( clk ), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_3257, signal_3256, signal_1366}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1352 ( .a ({signal_8156, signal_8154, signal_8152}), .b ({signal_2661, signal_2660, signal_1068}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({signal_3259, signal_3258, signal_1367}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1358 ( .a ({signal_8096, signal_8094, signal_8092}), .b ({signal_2685, signal_2684, signal_1080}), .clk ( clk ), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_3271, signal_3270, signal_1373}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1359 ( .a ({signal_8126, signal_8124, signal_8122}), .b ({signal_2695, signal_2694, signal_1085}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({signal_3273, signal_3272, signal_1374}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1363 ( .a ({signal_8114, signal_8112, signal_8110}), .b ({signal_2703, signal_2702, signal_1089}), .clk ( clk ), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_3281, signal_3280, signal_1378}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1364 ( .a ({signal_8162, signal_8160, signal_8158}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({signal_3283, signal_3282, signal_1379}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1370 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2675, signal_2674, signal_1075}), .clk ( clk ), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_3295, signal_3294, signal_1385}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1371 ( .a ({signal_8174, signal_8172, signal_8170}), .b ({signal_2715, signal_2714, signal_1095}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({signal_3297, signal_3296, signal_1386}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1372 ( .a ({signal_8180, signal_8178, signal_8176}), .b ({signal_2715, signal_2714, signal_1095}), .clk ( clk ), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_3299, signal_3298, signal_1387}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1373 ( .a ({signal_2671, signal_2670, signal_1073}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({signal_3301, signal_3300, signal_1388}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1374 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2719, signal_2718, signal_1097}), .clk ( clk ), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_3303, signal_3302, signal_1389}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1377 ( .a ({signal_8192, signal_8190, signal_8188}), .b ({signal_2733, signal_2732, signal_1104}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({signal_3309, signal_3308, signal_1392}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1378 ( .a ({signal_8198, signal_8196, signal_8194}), .b ({signal_2681, signal_2680, signal_1078}), .clk ( clk ), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_3311, signal_3310, signal_1393}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1379 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({signal_3313, signal_3312, signal_1394}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1380 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2703, signal_2702, signal_1089}), .clk ( clk ), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_3315, signal_3314, signal_1395}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1381 ( .a ({signal_8114, signal_8112, signal_8110}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({signal_3317, signal_3316, signal_1396}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1382 ( .a ({signal_8204, signal_8202, signal_8200}), .b ({signal_2671, signal_2670, signal_1073}), .clk ( clk ), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_3319, signal_3318, signal_1397}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1384 ( .a ({signal_8210, signal_8208, signal_8206}), .b ({signal_2739, signal_2738, signal_1107}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({signal_3323, signal_3322, signal_1399}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1385 ( .a ({signal_8102, signal_8100, signal_8098}), .b ({signal_2709, signal_2708, signal_1092}), .clk ( clk ), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_3325, signal_3324, signal_1400}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1386 ( .a ({signal_8216, signal_8214, signal_8212}), .b ({signal_2685, signal_2684, signal_1080}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({signal_3327, signal_3326, signal_1401}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1387 ( .a ({signal_8222, signal_8220, signal_8218}), .b ({signal_2697, signal_2696, signal_1086}), .clk ( clk ), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_3329, signal_3328, signal_1402}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1388 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_2753, signal_2752, signal_1114}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({signal_3331, signal_3330, signal_1403}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1389 ( .a ({signal_8234, signal_8232, signal_8230}), .b ({signal_2741, signal_2740, signal_1108}), .clk ( clk ), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_3333, signal_3332, signal_1404}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1390 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({signal_3335, signal_3334, signal_1405}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1391 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_2719, signal_2718, signal_1097}), .clk ( clk ), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_3337, signal_3336, signal_1406}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1392 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({signal_3339, signal_3338, signal_1407}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1393 ( .a ({signal_8240, signal_8238, signal_8236}), .b ({signal_2715, signal_2714, signal_1095}), .clk ( clk ), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_3341, signal_3340, signal_1408}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1394 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2753, signal_2752, signal_1114}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({signal_3343, signal_3342, signal_1409}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1397 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2729, signal_2728, signal_1102}), .clk ( clk ), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_3349, signal_3348, signal_1412}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1398 ( .a ({signal_8144, signal_8142, signal_8140}), .b ({signal_2771, signal_2770, signal_1123}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({signal_3351, signal_3350, signal_1413}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1399 ( .a ({signal_8246, signal_8244, signal_8242}), .b ({signal_2675, signal_2674, signal_1075}), .clk ( clk ), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_3353, signal_3352, signal_1414}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1400 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2715, signal_2714, signal_1095}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({signal_3355, signal_3354, signal_1415}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1404 ( .a ({signal_8180, signal_8178, signal_8176}), .b ({signal_2681, signal_2680, signal_1078}), .clk ( clk ), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_3363, signal_3362, signal_1419}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1405 ( .a ({signal_8114, signal_8112, signal_8110}), .b ({signal_2729, signal_2728, signal_1102}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({signal_3365, signal_3364, signal_1420}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1406 ( .a ({signal_8252, signal_8250, signal_8248}), .b ({signal_2755, signal_2754, signal_1115}), .clk ( clk ), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_3367, signal_3366, signal_1421}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1409 ( .a ({signal_8258, signal_8256, signal_8254}), .b ({signal_2671, signal_2670, signal_1073}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({signal_3373, signal_3372, signal_1424}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1410 ( .a ({signal_8072, signal_8070, signal_8068}), .b ({signal_2739, signal_2738, signal_1107}), .clk ( clk ), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_3375, signal_3374, signal_1425}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1411 ( .a ({signal_8180, signal_8178, signal_8176}), .b ({signal_2697, signal_2696, signal_1086}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({signal_3377, signal_3376, signal_1426}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1412 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_2781, signal_2780, signal_1128}), .clk ( clk ), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_3379, signal_3378, signal_1427}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1413 ( .a ({signal_8264, signal_8262, signal_8260}), .b ({signal_2669, signal_2668, signal_1072}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({signal_3381, signal_3380, signal_1428}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1414 ( .a ({signal_8270, signal_8268, signal_8266}), .b ({signal_2791, signal_2790, signal_1133}), .clk ( clk ), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_3383, signal_3382, signal_1429}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1415 ( .a ({signal_8174, signal_8172, signal_8170}), .b ({signal_2675, signal_2674, signal_1075}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({signal_3385, signal_3384, signal_1430}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1416 ( .a ({signal_8282, signal_8278, signal_8274}), .b ({signal_2801, signal_2800, signal_1138}), .clk ( clk ), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_3387, signal_3386, signal_1431}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1417 ( .a ({signal_8144, signal_8142, signal_8140}), .b ({signal_2675, signal_2674, signal_1075}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({signal_3389, signal_3388, signal_1432}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1418 ( .a ({signal_8288, signal_8286, signal_8284}), .b ({signal_2805, signal_2804, signal_1140}), .clk ( clk ), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_3391, signal_3390, signal_1433}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1419 ( .a ({signal_8294, signal_8292, signal_8290}), .b ({signal_2671, signal_2670, signal_1073}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({signal_3393, signal_3392, signal_1434}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1420 ( .a ({signal_8156, signal_8154, signal_8152}), .b ({signal_2809, signal_2808, signal_1142}), .clk ( clk ), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_3395, signal_3394, signal_1435}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1421 ( .a ({signal_8246, signal_8244, signal_8242}), .b ({signal_2693, signal_2692, signal_1084}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({signal_3397, signal_3396, signal_1436}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1422 ( .a ({signal_8156, signal_8154, signal_8152}), .b ({signal_2675, signal_2674, signal_1075}), .clk ( clk ), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_3399, signal_3398, signal_1437}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1423 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2827, signal_2826, signal_1151}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({signal_3401, signal_3400, signal_1438}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1424 ( .a ({signal_8300, signal_8298, signal_8296}), .b ({signal_2831, signal_2830, signal_1153}), .clk ( clk ), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_3403, signal_3402, signal_1439}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1425 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2837, signal_2836, signal_1156}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({signal_3405, signal_3404, signal_1440}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1426 ( .a ({signal_8192, signal_8190, signal_8188}), .b ({signal_2841, signal_2840, signal_1158}), .clk ( clk ), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_3407, signal_3406, signal_1441}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1427 ( .a ({signal_8156, signal_8154, signal_8152}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({signal_3409, signal_3408, signal_1442}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1428 ( .a ({signal_8252, signal_8250, signal_8248}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_3411, signal_3410, signal_1443}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1429 ( .a ({signal_8150, signal_8148, signal_8146}), .b ({signal_2857, signal_2856, signal_1166}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({signal_3413, signal_3412, signal_1444}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1430 ( .a ({signal_2697, signal_2696, signal_1086}), .b ({signal_2567, signal_2566, signal_1021}), .clk ( clk ), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_3415, signal_3414, signal_1445}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1431 ( .a ({signal_8306, signal_8304, signal_8302}), .b ({signal_2861, signal_2860, signal_1168}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({signal_3417, signal_3416, signal_1446}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1432 ( .a ({signal_2569, signal_2568, signal_1022}), .b ({signal_2809, signal_2808, signal_1142}), .clk ( clk ), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_3419, signal_3418, signal_1447}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1433 ( .a ({signal_8102, signal_8100, signal_8098}), .b ({signal_2797, signal_2796, signal_1136}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({signal_3421, signal_3420, signal_1448}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1434 ( .a ({signal_2811, signal_2810, signal_1143}), .b ({signal_2815, signal_2814, signal_1145}), .clk ( clk ), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_3423, signal_3422, signal_1449}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1435 ( .a ({signal_8210, signal_8208, signal_8206}), .b ({signal_2857, signal_2856, signal_1166}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({signal_3425, signal_3424, signal_1450}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1436 ( .a ({signal_8312, signal_8310, signal_8308}), .b ({signal_2831, signal_2830, signal_1153}), .clk ( clk ), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_3427, signal_3426, signal_1451}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1437 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_2877, signal_2876, signal_1176}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({signal_3429, signal_3428, signal_1452}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1438 ( .a ({signal_2797, signal_2796, signal_1136}), .b ({signal_2831, signal_2830, signal_1153}), .clk ( clk ), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_3431, signal_3430, signal_1453}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1439 ( .a ({signal_2707, signal_2706, signal_1091}), .b ({signal_2841, signal_2840, signal_1158}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({signal_3433, signal_3432, signal_1454}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1440 ( .a ({signal_8132, signal_8130, signal_8128}), .b ({signal_2839, signal_2838, signal_1157}), .clk ( clk ), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_3435, signal_3434, signal_1455}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1441 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_2881, signal_2880, signal_1178}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({signal_3437, signal_3436, signal_1456}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1442 ( .a ({signal_8258, signal_8256, signal_8254}), .b ({signal_2689, signal_2688, signal_1082}), .clk ( clk ), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_3439, signal_3438, signal_1457}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1443 ( .a ({signal_8270, signal_8268, signal_8266}), .b ({signal_2841, signal_2840, signal_1158}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({signal_3441, signal_3440, signal_1458}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1444 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2691, signal_2690, signal_1083}), .clk ( clk ), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_3443, signal_3442, signal_1459}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1445 ( .a ({signal_8174, signal_8172, signal_8170}), .b ({signal_2903, signal_2902, signal_1189}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({signal_3445, signal_3444, signal_1460}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1446 ( .a ({signal_8318, signal_8316, signal_8314}), .b ({signal_2905, signal_2904, signal_1190}), .clk ( clk ), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_3447, signal_3446, signal_1461}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1447 ( .a ({signal_8174, signal_8172, signal_8170}), .b ({signal_2811, signal_2810, signal_1143}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({signal_3449, signal_3448, signal_1462}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1448 ( .a ({signal_8324, signal_8322, signal_8320}), .b ({signal_2839, signal_2838, signal_1157}), .clk ( clk ), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_3451, signal_3450, signal_1463}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1449 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_2671, signal_2670, signal_1073}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({signal_3453, signal_3452, signal_1464}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1450 ( .a ({signal_8300, signal_8298, signal_8296}), .b ({signal_2841, signal_2840, signal_1158}), .clk ( clk ), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_3455, signal_3454, signal_1465}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1451 ( .a ({signal_8330, signal_8328, signal_8326}), .b ({signal_2921, signal_2920, signal_1198}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({signal_3457, signal_3456, signal_1466}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1452 ( .a ({signal_8336, signal_8334, signal_8332}), .b ({signal_2815, signal_2814, signal_1145}), .clk ( clk ), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_3459, signal_3458, signal_1467}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1453 ( .a ({signal_8342, signal_8340, signal_8338}), .b ({signal_2909, signal_2908, signal_1192}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({signal_3461, signal_3460, signal_1468}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1454 ( .a ({signal_2729, signal_2728, signal_1102}), .b ({signal_2841, signal_2840, signal_1158}), .clk ( clk ), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_3463, signal_3462, signal_1469}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1455 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_2879, signal_2878, signal_1177}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({signal_3465, signal_3464, signal_1470}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1456 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2689, signal_2688, signal_1082}), .clk ( clk ), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_3467, signal_3466, signal_1471}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1457 ( .a ({signal_8252, signal_8250, signal_8248}), .b ({signal_2907, signal_2906, signal_1191}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({signal_3469, signal_3468, signal_1472}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1458 ( .a ({signal_8204, signal_8202, signal_8200}), .b ({signal_2813, signal_2812, signal_1144}), .clk ( clk ), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_3471, signal_3470, signal_1473}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1459 ( .a ({signal_8174, signal_8172, signal_8170}), .b ({signal_2879, signal_2878, signal_1177}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({signal_3473, signal_3472, signal_1474}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1460 ( .a ({signal_8234, signal_8232, signal_8230}), .b ({signal_2897, signal_2896, signal_1186}), .clk ( clk ), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_3475, signal_3474, signal_1475}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1461 ( .a ({signal_8180, signal_8178, signal_8176}), .b ({signal_2693, signal_2692, signal_1084}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({signal_3477, signal_3476, signal_1476}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1462 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2689, signal_2688, signal_1082}), .clk ( clk ), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_3479, signal_3478, signal_1477}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1463 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2937, signal_2936, signal_1206}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({signal_3481, signal_3480, signal_1478}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1464 ( .a ({signal_8270, signal_8268, signal_8266}), .b ({signal_2831, signal_2830, signal_1153}), .clk ( clk ), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_3483, signal_3482, signal_1479}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1465 ( .a ({signal_8096, signal_8094, signal_8092}), .b ({signal_2897, signal_2896, signal_1186}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({signal_3485, signal_3484, signal_1480}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1466 ( .a ({signal_2675, signal_2674, signal_1075}), .b ({signal_2687, signal_2686, signal_1081}), .clk ( clk ), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_3487, signal_3486, signal_1481}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1467 ( .a ({signal_8120, signal_8118, signal_8116}), .b ({signal_2861, signal_2860, signal_1168}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({signal_3489, signal_3488, signal_1482}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1468 ( .a ({signal_8252, signal_8250, signal_8248}), .b ({signal_2847, signal_2846, signal_1161}), .clk ( clk ), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_3491, signal_3490, signal_1483}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1469 ( .a ({signal_2567, signal_2566, signal_1021}), .b ({signal_2789, signal_2788, signal_1132}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({signal_3493, signal_3492, signal_1484}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1470 ( .a ({signal_8222, signal_8220, signal_8218}), .b ({signal_2693, signal_2692, signal_1084}), .clk ( clk ), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_3495, signal_3494, signal_1485}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1471 ( .a ({signal_8348, signal_8346, signal_8344}), .b ({signal_2941, signal_2940, signal_1208}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({signal_3497, signal_3496, signal_1486}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1472 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2693, signal_2692, signal_1084}), .clk ( clk ), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_3499, signal_3498, signal_1487}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1473 ( .a ({signal_8204, signal_8202, signal_8200}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({signal_3501, signal_3500, signal_1488}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1474 ( .a ({signal_8354, signal_8352, signal_8350}), .b ({signal_2927, signal_2926, signal_1201}), .clk ( clk ), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_3503, signal_3502, signal_1489}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1475 ( .a ({signal_8114, signal_8112, signal_8110}), .b ({signal_2847, signal_2846, signal_1161}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({signal_3505, signal_3504, signal_1490}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1476 ( .a ({signal_8066, signal_8062, signal_8058}), .b ({signal_2811, signal_2810, signal_1143}), .clk ( clk ), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_3507, signal_3506, signal_1491}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1477 ( .a ({signal_8270, signal_8268, signal_8266}), .b ({signal_2959, signal_2958, signal_1217}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({signal_3509, signal_3508, signal_1492}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1478 ( .a ({signal_8264, signal_8262, signal_8260}), .b ({signal_2715, signal_2714, signal_1095}), .clk ( clk ), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_3511, signal_3510, signal_1493}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1479 ( .a ({signal_8066, signal_8062, signal_8058}), .b ({signal_2903, signal_2902, signal_1189}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({signal_3513, signal_3512, signal_1494}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1480 ( .a ({signal_8360, signal_8358, signal_8356}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_3515, signal_3514, signal_1495}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1481 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_2671, signal_2670, signal_1073}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({signal_3517, signal_3516, signal_1496}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1482 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2813, signal_2812, signal_1144}), .clk ( clk ), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_3519, signal_3518, signal_1497}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1483 ( .a ({signal_8180, signal_8178, signal_8176}), .b ({signal_2813, signal_2812, signal_1144}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({signal_3521, signal_3520, signal_1498}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1484 ( .a ({signal_8144, signal_8142, signal_8140}), .b ({signal_2811, signal_2810, signal_1143}), .clk ( clk ), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_3523, signal_3522, signal_1499}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1485 ( .a ({signal_8066, signal_8062, signal_8058}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({signal_3525, signal_3524, signal_1500}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1486 ( .a ({signal_8258, signal_8256, signal_8254}), .b ({signal_2849, signal_2848, signal_1162}), .clk ( clk ), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_3527, signal_3526, signal_1501}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1487 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_2811, signal_2810, signal_1143}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({signal_3529, signal_3528, signal_1502}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1488 ( .a ({signal_8186, signal_8184, signal_8182}), .b ({signal_2811, signal_2810, signal_1143}), .clk ( clk ), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_3531, signal_3530, signal_1503}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1489 ( .a ({signal_8150, signal_8148, signal_8146}), .b ({signal_2763, signal_2762, signal_1119}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({signal_3533, signal_3532, signal_1504}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1490 ( .a ({signal_3257, signal_3256, signal_1366}), .b ({signal_3535, signal_3534, signal_1505}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1491 ( .a ({signal_3259, signal_3258, signal_1367}), .b ({signal_3537, signal_3536, signal_1506}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1497 ( .a ({signal_3271, signal_3270, signal_1373}), .b ({signal_3549, signal_3548, signal_1512}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1498 ( .a ({signal_3273, signal_3272, signal_1374}), .b ({signal_3551, signal_3550, signal_1513}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1502 ( .a ({signal_3281, signal_3280, signal_1378}), .b ({signal_3559, signal_3558, signal_1517}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1503 ( .a ({signal_3283, signal_3282, signal_1379}), .b ({signal_3561, signal_3560, signal_1518}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1508 ( .a ({signal_3295, signal_3294, signal_1385}), .b ({signal_3571, signal_3570, signal_1523}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1509 ( .a ({signal_3297, signal_3296, signal_1386}), .b ({signal_3573, signal_3572, signal_1524}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1510 ( .a ({signal_3299, signal_3298, signal_1387}), .b ({signal_3575, signal_3574, signal_1525}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1511 ( .a ({signal_3301, signal_3300, signal_1388}), .b ({signal_3577, signal_3576, signal_1526}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1512 ( .a ({signal_3303, signal_3302, signal_1389}), .b ({signal_3579, signal_3578, signal_1527}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1514 ( .a ({signal_3309, signal_3308, signal_1392}), .b ({signal_3583, signal_3582, signal_1529}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1515 ( .a ({signal_3311, signal_3310, signal_1393}), .b ({signal_3585, signal_3584, signal_1530}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1516 ( .a ({signal_3313, signal_3312, signal_1394}), .b ({signal_3587, signal_3586, signal_1531}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1517 ( .a ({signal_3315, signal_3314, signal_1395}), .b ({signal_3589, signal_3588, signal_1532}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1518 ( .a ({signal_3317, signal_3316, signal_1396}), .b ({signal_3591, signal_3590, signal_1533}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1519 ( .a ({signal_3319, signal_3318, signal_1397}), .b ({signal_3593, signal_3592, signal_1534}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1521 ( .a ({signal_3323, signal_3322, signal_1399}), .b ({signal_3597, signal_3596, signal_1536}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1522 ( .a ({signal_3325, signal_3324, signal_1400}), .b ({signal_3599, signal_3598, signal_1537}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1523 ( .a ({signal_3327, signal_3326, signal_1401}), .b ({signal_3601, signal_3600, signal_1538}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1524 ( .a ({signal_3329, signal_3328, signal_1402}), .b ({signal_3603, signal_3602, signal_1539}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1525 ( .a ({signal_3331, signal_3330, signal_1403}), .b ({signal_3605, signal_3604, signal_1540}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1526 ( .a ({signal_3333, signal_3332, signal_1404}), .b ({signal_3607, signal_3606, signal_1541}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1527 ( .a ({signal_3335, signal_3334, signal_1405}), .b ({signal_3609, signal_3608, signal_1542}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1528 ( .a ({signal_3337, signal_3336, signal_1406}), .b ({signal_3611, signal_3610, signal_1543}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1529 ( .a ({signal_3339, signal_3338, signal_1407}), .b ({signal_3613, signal_3612, signal_1544}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1530 ( .a ({signal_3341, signal_3340, signal_1408}), .b ({signal_3615, signal_3614, signal_1545}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1531 ( .a ({signal_3343, signal_3342, signal_1409}), .b ({signal_3617, signal_3616, signal_1546}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1534 ( .a ({signal_3349, signal_3348, signal_1412}), .b ({signal_3623, signal_3622, signal_1549}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1535 ( .a ({signal_3351, signal_3350, signal_1413}), .b ({signal_3625, signal_3624, signal_1550}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1536 ( .a ({signal_3353, signal_3352, signal_1414}), .b ({signal_3627, signal_3626, signal_1551}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1537 ( .a ({signal_3355, signal_3354, signal_1415}), .b ({signal_3629, signal_3628, signal_1552}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1540 ( .a ({signal_3363, signal_3362, signal_1419}), .b ({signal_3635, signal_3634, signal_1555}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1541 ( .a ({signal_3365, signal_3364, signal_1420}), .b ({signal_3637, signal_3636, signal_1556}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1542 ( .a ({signal_3367, signal_3366, signal_1421}), .b ({signal_3639, signal_3638, signal_1557}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1545 ( .a ({signal_3373, signal_3372, signal_1424}), .b ({signal_3645, signal_3644, signal_1560}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1546 ( .a ({signal_3375, signal_3374, signal_1425}), .b ({signal_3647, signal_3646, signal_1561}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1547 ( .a ({signal_3377, signal_3376, signal_1426}), .b ({signal_3649, signal_3648, signal_1562}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1548 ( .a ({signal_3379, signal_3378, signal_1427}), .b ({signal_3651, signal_3650, signal_1563}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1549 ( .a ({signal_3381, signal_3380, signal_1428}), .b ({signal_3653, signal_3652, signal_1564}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1550 ( .a ({signal_3383, signal_3382, signal_1429}), .b ({signal_3655, signal_3654, signal_1565}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1551 ( .a ({signal_3385, signal_3384, signal_1430}), .b ({signal_3657, signal_3656, signal_1566}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1552 ( .a ({signal_3387, signal_3386, signal_1431}), .b ({signal_3659, signal_3658, signal_1567}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1553 ( .a ({signal_3389, signal_3388, signal_1432}), .b ({signal_3661, signal_3660, signal_1568}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1554 ( .a ({signal_3391, signal_3390, signal_1433}), .b ({signal_3663, signal_3662, signal_1569}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1555 ( .a ({signal_3393, signal_3392, signal_1434}), .b ({signal_3665, signal_3664, signal_1570}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1556 ( .a ({signal_3395, signal_3394, signal_1435}), .b ({signal_3667, signal_3666, signal_1571}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1557 ( .a ({signal_3397, signal_3396, signal_1436}), .b ({signal_3669, signal_3668, signal_1572}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1558 ( .a ({signal_3399, signal_3398, signal_1437}), .b ({signal_3671, signal_3670, signal_1573}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1559 ( .a ({signal_3401, signal_3400, signal_1438}), .b ({signal_3673, signal_3672, signal_1574}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1560 ( .a ({signal_3403, signal_3402, signal_1439}), .b ({signal_3675, signal_3674, signal_1575}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1561 ( .a ({signal_3405, signal_3404, signal_1440}), .b ({signal_3677, signal_3676, signal_1576}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1562 ( .a ({signal_3407, signal_3406, signal_1441}), .b ({signal_3679, signal_3678, signal_1577}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1563 ( .a ({signal_3409, signal_3408, signal_1442}), .b ({signal_3681, signal_3680, signal_1578}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1564 ( .a ({signal_3411, signal_3410, signal_1443}), .b ({signal_3683, signal_3682, signal_1579}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1565 ( .a ({signal_3413, signal_3412, signal_1444}), .b ({signal_3685, signal_3684, signal_1580}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1566 ( .a ({signal_3415, signal_3414, signal_1445}), .b ({signal_3687, signal_3686, signal_1581}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1567 ( .a ({signal_3419, signal_3418, signal_1447}), .b ({signal_3689, signal_3688, signal_1582}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1568 ( .a ({signal_3421, signal_3420, signal_1448}), .b ({signal_3691, signal_3690, signal_1583}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1569 ( .a ({signal_3423, signal_3422, signal_1449}), .b ({signal_3693, signal_3692, signal_1584}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1570 ( .a ({signal_3425, signal_3424, signal_1450}), .b ({signal_3695, signal_3694, signal_1585}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1571 ( .a ({signal_3427, signal_3426, signal_1451}), .b ({signal_3697, signal_3696, signal_1586}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1572 ( .a ({signal_3429, signal_3428, signal_1452}), .b ({signal_3699, signal_3698, signal_1587}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1573 ( .a ({signal_3431, signal_3430, signal_1453}), .b ({signal_3701, signal_3700, signal_1588}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1574 ( .a ({signal_3433, signal_3432, signal_1454}), .b ({signal_3703, signal_3702, signal_1589}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1575 ( .a ({signal_3435, signal_3434, signal_1455}), .b ({signal_3705, signal_3704, signal_1590}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1576 ( .a ({signal_3437, signal_3436, signal_1456}), .b ({signal_3707, signal_3706, signal_1591}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1577 ( .a ({signal_3439, signal_3438, signal_1457}), .b ({signal_3709, signal_3708, signal_1592}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1578 ( .a ({signal_3441, signal_3440, signal_1458}), .b ({signal_3711, signal_3710, signal_1593}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1579 ( .a ({signal_3443, signal_3442, signal_1459}), .b ({signal_3713, signal_3712, signal_1594}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1580 ( .a ({signal_3445, signal_3444, signal_1460}), .b ({signal_3715, signal_3714, signal_1595}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1581 ( .a ({signal_3449, signal_3448, signal_1462}), .b ({signal_3717, signal_3716, signal_1596}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1582 ( .a ({signal_3451, signal_3450, signal_1463}), .b ({signal_3719, signal_3718, signal_1597}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1583 ( .a ({signal_3453, signal_3452, signal_1464}), .b ({signal_3721, signal_3720, signal_1598}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1584 ( .a ({signal_3455, signal_3454, signal_1465}), .b ({signal_3723, signal_3722, signal_1599}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1585 ( .a ({signal_3457, signal_3456, signal_1466}), .b ({signal_3725, signal_3724, signal_1600}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1586 ( .a ({signal_3459, signal_3458, signal_1467}), .b ({signal_3727, signal_3726, signal_1601}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1587 ( .a ({signal_3461, signal_3460, signal_1468}), .b ({signal_3729, signal_3728, signal_1602}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1588 ( .a ({signal_3463, signal_3462, signal_1469}), .b ({signal_3731, signal_3730, signal_1603}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1589 ( .a ({signal_3465, signal_3464, signal_1470}), .b ({signal_3733, signal_3732, signal_1604}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1590 ( .a ({signal_3467, signal_3466, signal_1471}), .b ({signal_3735, signal_3734, signal_1605}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1591 ( .a ({signal_3469, signal_3468, signal_1472}), .b ({signal_3737, signal_3736, signal_1606}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1592 ( .a ({signal_3471, signal_3470, signal_1473}), .b ({signal_3739, signal_3738, signal_1607}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1593 ( .a ({signal_3473, signal_3472, signal_1474}), .b ({signal_3741, signal_3740, signal_1608}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1594 ( .a ({signal_3475, signal_3474, signal_1475}), .b ({signal_3743, signal_3742, signal_1609}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1595 ( .a ({signal_3477, signal_3476, signal_1476}), .b ({signal_3745, signal_3744, signal_1610}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1596 ( .a ({signal_3479, signal_3478, signal_1477}), .b ({signal_3747, signal_3746, signal_1611}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1597 ( .a ({signal_3483, signal_3482, signal_1479}), .b ({signal_3749, signal_3748, signal_1612}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1598 ( .a ({signal_3485, signal_3484, signal_1480}), .b ({signal_3751, signal_3750, signal_1613}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1599 ( .a ({signal_3487, signal_3486, signal_1481}), .b ({signal_3753, signal_3752, signal_1614}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1600 ( .a ({signal_3489, signal_3488, signal_1482}), .b ({signal_3755, signal_3754, signal_1615}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1601 ( .a ({signal_3491, signal_3490, signal_1483}), .b ({signal_3757, signal_3756, signal_1616}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1602 ( .a ({signal_3493, signal_3492, signal_1484}), .b ({signal_3759, signal_3758, signal_1617}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1603 ( .a ({signal_3495, signal_3494, signal_1485}), .b ({signal_3761, signal_3760, signal_1618}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1604 ( .a ({signal_3497, signal_3496, signal_1486}), .b ({signal_3763, signal_3762, signal_1619}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1605 ( .a ({signal_3499, signal_3498, signal_1487}), .b ({signal_3765, signal_3764, signal_1620}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1606 ( .a ({signal_3501, signal_3500, signal_1488}), .b ({signal_3767, signal_3766, signal_1621}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1607 ( .a ({signal_3503, signal_3502, signal_1489}), .b ({signal_3769, signal_3768, signal_1622}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1608 ( .a ({signal_3505, signal_3504, signal_1490}), .b ({signal_3771, signal_3770, signal_1623}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1609 ( .a ({signal_3507, signal_3506, signal_1491}), .b ({signal_3773, signal_3772, signal_1624}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1610 ( .a ({signal_3509, signal_3508, signal_1492}), .b ({signal_3775, signal_3774, signal_1625}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1611 ( .a ({signal_3511, signal_3510, signal_1493}), .b ({signal_3777, signal_3776, signal_1626}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1612 ( .a ({signal_3513, signal_3512, signal_1494}), .b ({signal_3779, signal_3778, signal_1627}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1613 ( .a ({signal_3515, signal_3514, signal_1495}), .b ({signal_3781, signal_3780, signal_1628}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1614 ( .a ({signal_3517, signal_3516, signal_1496}), .b ({signal_3783, signal_3782, signal_1629}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1615 ( .a ({signal_3519, signal_3518, signal_1497}), .b ({signal_3785, signal_3784, signal_1630}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1616 ( .a ({signal_3521, signal_3520, signal_1498}), .b ({signal_3787, signal_3786, signal_1631}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1617 ( .a ({signal_3523, signal_3522, signal_1499}), .b ({signal_3789, signal_3788, signal_1632}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1618 ( .a ({signal_3525, signal_3524, signal_1500}), .b ({signal_3791, signal_3790, signal_1633}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1619 ( .a ({signal_3527, signal_3526, signal_1501}), .b ({signal_3793, signal_3792, signal_1634}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1620 ( .a ({signal_3529, signal_3528, signal_1502}), .b ({signal_3795, signal_3794, signal_1635}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1621 ( .a ({signal_3531, signal_3530, signal_1503}), .b ({signal_3797, signal_3796, signal_1636}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1622 ( .a ({signal_3533, signal_3532, signal_1504}), .b ({signal_3799, signal_3798, signal_1637}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1623 ( .a ({signal_8342, signal_8340, signal_8338}), .b ({signal_2985, signal_2984, signal_1230}), .clk ( clk ), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_3801, signal_3800, signal_1638}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1624 ( .a ({signal_8366, signal_8364, signal_8362}), .b ({signal_2987, signal_2986, signal_1231}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({signal_3803, signal_3802, signal_1639}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1625 ( .a ({signal_8258, signal_8256, signal_8254}), .b ({signal_2997, signal_2996, signal_1236}), .clk ( clk ), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_3805, signal_3804, signal_1640}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1626 ( .a ({signal_2995, signal_2994, signal_1235}), .b ({signal_3037, signal_3036, signal_1256}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({signal_3807, signal_3806, signal_1641}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1627 ( .a ({signal_8372, signal_8370, signal_8368}), .b ({signal_3039, signal_3038, signal_1257}), .clk ( clk ), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_3809, signal_3808, signal_1642}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1628 ( .a ({signal_8354, signal_8352, signal_8350}), .b ({signal_3051, signal_3050, signal_1263}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({signal_3811, signal_3810, signal_1643}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1629 ( .a ({signal_3025, signal_3024, signal_1250}), .b ({signal_3031, signal_3030, signal_1253}), .clk ( clk ), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_3813, signal_3812, signal_1644}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1630 ( .a ({signal_3059, signal_3058, signal_1267}), .b ({signal_3061, signal_3060, signal_1268}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({signal_3815, signal_3814, signal_1645}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1631 ( .a ({signal_8378, signal_8376, signal_8374}), .b ({signal_3005, signal_3004, signal_1240}), .clk ( clk ), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_3817, signal_3816, signal_1646}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1632 ( .a ({signal_3063, signal_3062, signal_1269}), .b ({signal_3065, signal_3064, signal_1270}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({signal_3819, signal_3818, signal_1647}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1633 ( .a ({signal_2995, signal_2994, signal_1235}), .b ({signal_3035, signal_3034, signal_1255}), .clk ( clk ), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_3821, signal_3820, signal_1648}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1634 ( .a ({signal_3071, signal_3070, signal_1273}), .b ({signal_3073, signal_3072, signal_1274}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({signal_3823, signal_3822, signal_1649}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1635 ( .a ({signal_2635, signal_2634, signal_1055}), .b ({signal_3033, signal_3032, signal_1254}), .clk ( clk ), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_3825, signal_3824, signal_1650}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1636 ( .a ({signal_8360, signal_8358, signal_8356}), .b ({signal_3007, signal_3006, signal_1241}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({signal_3827, signal_3826, signal_1651}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1637 ( .a ({signal_2997, signal_2996, signal_1236}), .b ({signal_2643, signal_2642, signal_1059}), .clk ( clk ), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_3829, signal_3828, signal_1652}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1638 ( .a ({signal_3085, signal_3084, signal_1280}), .b ({signal_3087, signal_3086, signal_1281}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({signal_3831, signal_3830, signal_1653}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1639 ( .a ({signal_3091, signal_3090, signal_1283}), .b ({signal_3093, signal_3092, signal_1284}), .clk ( clk ), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_3833, signal_3832, signal_1654}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1640 ( .a ({signal_2991, signal_2990, signal_1233}), .b ({signal_3097, signal_3096, signal_1286}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({signal_3835, signal_3834, signal_1655}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1641 ( .a ({signal_2999, signal_2998, signal_1237}), .b ({signal_3101, signal_3100, signal_1288}), .clk ( clk ), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_3837, signal_3836, signal_1656}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1642 ( .a ({signal_2643, signal_2642, signal_1059}), .b ({signal_3001, signal_3000, signal_1238}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({signal_3839, signal_3838, signal_1657}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1643 ( .a ({signal_3009, signal_3008, signal_1242}), .b ({signal_3011, signal_3010, signal_1243}), .clk ( clk ), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_3841, signal_3840, signal_1658}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1645 ( .a ({signal_3113, signal_3112, signal_1294}), .b ({signal_3115, signal_3114, signal_1295}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({signal_3845, signal_3844, signal_1660}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1646 ( .a ({signal_3001, signal_3000, signal_1238}), .b ({signal_3129, signal_3128, signal_1302}), .clk ( clk ), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_3847, signal_3846, signal_1661}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1647 ( .a ({signal_8384, signal_8382, signal_8380}), .b ({signal_3137, signal_3136, signal_1306}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({signal_3849, signal_3848, signal_1662}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1648 ( .a ({signal_3029, signal_3028, signal_1252}), .b ({signal_3145, signal_3144, signal_1310}), .clk ( clk ), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_3851, signal_3850, signal_1663}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1649 ( .a ({signal_8390, signal_8388, signal_8386}), .b ({signal_3291, signal_3290, signal_1383}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({signal_3853, signal_3852, signal_1664}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1650 ( .a ({signal_8066, signal_8062, signal_8058}), .b ({signal_3119, signal_3118, signal_1297}), .clk ( clk ), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_3855, signal_3854, signal_1665}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1651 ( .a ({signal_3013, signal_3012, signal_1244}), .b ({signal_3147, signal_3146, signal_1311}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({signal_3857, signal_3856, signal_1666}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1653 ( .a ({signal_3277, signal_3276, signal_1376}), .b ({signal_3159, signal_3158, signal_1317}), .clk ( clk ), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_3861, signal_3860, signal_1668}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1654 ( .a ({signal_2995, signal_2994, signal_1235}), .b ({signal_3163, signal_3162, signal_1319}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({signal_3863, signal_3862, signal_1669}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1655 ( .a ({signal_3305, signal_3304, signal_1390}), .b ({signal_2655, signal_2654, signal_1065}), .clk ( clk ), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_3865, signal_3864, signal_1670}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1656 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_3165, signal_3164, signal_1320}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({signal_3867, signal_3866, signal_1671}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1657 ( .a ({signal_3045, signal_3044, signal_1260}), .b ({signal_3125, signal_3124, signal_1300}), .clk ( clk ), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_3869, signal_3868, signal_1672}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1658 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_3167, signal_3166, signal_1321}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({signal_3871, signal_3870, signal_1673}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1659 ( .a ({signal_3157, signal_3156, signal_1316}), .b ({signal_3169, signal_3168, signal_1322}), .clk ( clk ), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_3873, signal_3872, signal_1674}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1660 ( .a ({signal_2651, signal_2650, signal_1063}), .b ({signal_3171, signal_3170, signal_1323}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({signal_3875, signal_3874, signal_1675}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1661 ( .a ({signal_3173, signal_3172, signal_1324}), .b ({signal_3175, signal_3174, signal_1325}), .clk ( clk ), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_3877, signal_3876, signal_1676}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1663 ( .a ({signal_3005, signal_3004, signal_1240}), .b ({signal_3119, signal_3118, signal_1297}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({signal_3881, signal_3880, signal_1678}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1664 ( .a ({signal_3053, signal_3052, signal_1264}), .b ({signal_3187, signal_3186, signal_1331}), .clk ( clk ), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_3883, signal_3882, signal_1679}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1665 ( .a ({signal_3009, signal_3008, signal_1242}), .b ({signal_3189, signal_3188, signal_1332}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({signal_3885, signal_3884, signal_1680}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1666 ( .a ({signal_3057, signal_3056, signal_1266}), .b ({signal_3193, signal_3192, signal_1334}), .clk ( clk ), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_3887, signal_3886, signal_1681}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1667 ( .a ({signal_3119, signal_3118, signal_1297}), .b ({signal_3199, signal_3198, signal_1337}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({signal_3889, signal_3888, signal_1682}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1668 ( .a ({signal_3067, signal_3066, signal_1271}), .b ({signal_3187, signal_3186, signal_1331}), .clk ( clk ), .r ({Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_3891, signal_3890, signal_1683}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1669 ( .a ({signal_8132, signal_8130, signal_8128}), .b ({signal_3165, signal_3164, signal_1320}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233]}), .c ({signal_3893, signal_3892, signal_1684}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1670 ( .a ({signal_3103, signal_3102, signal_1289}), .b ({signal_3205, signal_3204, signal_1340}), .clk ( clk ), .r ({Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({signal_3895, signal_3894, signal_1685}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1671 ( .a ({signal_8396, signal_8394, signal_8392}), .b ({signal_3207, signal_3206, signal_1341}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239]}), .c ({signal_3897, signal_3896, signal_1686}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1673 ( .a ({signal_3077, signal_3076, signal_1276}), .b ({signal_3185, signal_3184, signal_1330}), .clk ( clk ), .r ({Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({signal_3901, signal_3900, signal_1688}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1674 ( .a ({signal_3161, signal_3160, signal_1318}), .b ({signal_3361, signal_3360, signal_1418}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245]}), .c ({signal_3903, signal_3902, signal_1689}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1675 ( .a ({signal_3043, signal_3042, signal_1259}), .b ({signal_3173, signal_3172, signal_1324}), .clk ( clk ), .r ({Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({signal_3905, signal_3904, signal_1690}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1676 ( .a ({signal_3079, signal_3078, signal_1277}), .b ({signal_3217, signal_3216, signal_1346}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251]}), .c ({signal_3907, signal_3906, signal_1691}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1677 ( .a ({signal_3219, signal_3218, signal_1347}), .b ({signal_3221, signal_3220, signal_1348}), .clk ( clk ), .r ({Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({signal_3909, signal_3908, signal_1692}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1678 ( .a ({signal_3025, signal_3024, signal_1250}), .b ({signal_3223, signal_3222, signal_1349}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257]}), .c ({signal_3911, signal_3910, signal_1693}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1679 ( .a ({signal_3227, signal_3226, signal_1351}), .b ({signal_3229, signal_3228, signal_1352}), .clk ( clk ), .r ({Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_3913, signal_3912, signal_1694}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1680 ( .a ({signal_2995, signal_2994, signal_1235}), .b ({signal_3143, signal_3142, signal_1309}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263]}), .c ({signal_3915, signal_3914, signal_1695}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1681 ( .a ({signal_3235, signal_3234, signal_1355}), .b ({signal_3237, signal_3236, signal_1356}), .clk ( clk ), .r ({Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({signal_3917, signal_3916, signal_1696}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1682 ( .a ({signal_3155, signal_3154, signal_1315}), .b ({signal_3239, signal_3238, signal_1357}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269]}), .c ({signal_3919, signal_3918, signal_1697}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1684 ( .a ({signal_3103, signal_3102, signal_1289}), .b ({signal_3105, signal_3104, signal_1290}), .clk ( clk ), .r ({Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({signal_3923, signal_3922, signal_1699}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1687 ( .a ({signal_3011, signal_3010, signal_1243}), .b ({signal_3105, signal_3104, signal_1290}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275]}), .c ({signal_3929, signal_3928, signal_1702}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1693 ( .a ({signal_3105, signal_3104, signal_1290}), .b ({signal_3135, signal_3134, signal_1305}), .clk ( clk ), .r ({Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({signal_3941, signal_3940, signal_1708}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1698 ( .a ({signal_3111, signal_3110, signal_1293}), .b ({signal_3253, signal_3252, signal_1364}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281]}), .c ({signal_3951, signal_3950, signal_1713}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1700 ( .a ({signal_3801, signal_3800, signal_1638}), .b ({signal_3955, signal_3954, signal_1715}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1701 ( .a ({signal_3803, signal_3802, signal_1639}), .b ({signal_3957, signal_3956, signal_1716}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1702 ( .a ({signal_3807, signal_3806, signal_1641}), .b ({signal_3959, signal_3958, signal_1717}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1703 ( .a ({signal_3809, signal_3808, signal_1642}), .b ({signal_3961, signal_3960, signal_1718}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1704 ( .a ({signal_3811, signal_3810, signal_1643}), .b ({signal_3963, signal_3962, signal_1719}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1705 ( .a ({signal_3813, signal_3812, signal_1644}), .b ({signal_3965, signal_3964, signal_1720}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1706 ( .a ({signal_3817, signal_3816, signal_1646}), .b ({signal_3967, signal_3966, signal_1721}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1707 ( .a ({signal_3819, signal_3818, signal_1647}), .b ({signal_3969, signal_3968, signal_1722}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1708 ( .a ({signal_3821, signal_3820, signal_1648}), .b ({signal_3971, signal_3970, signal_1723}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1709 ( .a ({signal_3825, signal_3824, signal_1650}), .b ({signal_3973, signal_3972, signal_1724}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1710 ( .a ({signal_3827, signal_3826, signal_1651}), .b ({signal_3975, signal_3974, signal_1725}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1711 ( .a ({signal_3829, signal_3828, signal_1652}), .b ({signal_3977, signal_3976, signal_1726}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1712 ( .a ({signal_3837, signal_3836, signal_1656}), .b ({signal_3979, signal_3978, signal_1727}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1713 ( .a ({signal_3839, signal_3838, signal_1657}), .b ({signal_3981, signal_3980, signal_1728}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1714 ( .a ({signal_3841, signal_3840, signal_1658}), .b ({signal_3983, signal_3982, signal_1729}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1716 ( .a ({signal_3849, signal_3848, signal_1662}), .b ({signal_3987, signal_3986, signal_1731}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1717 ( .a ({signal_3851, signal_3850, signal_1663}), .b ({signal_3989, signal_3988, signal_1732}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1718 ( .a ({signal_3853, signal_3852, signal_1664}), .b ({signal_3991, signal_3990, signal_1733}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1719 ( .a ({signal_3855, signal_3854, signal_1665}), .b ({signal_3993, signal_3992, signal_1734}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1720 ( .a ({signal_3857, signal_3856, signal_1666}), .b ({signal_3995, signal_3994, signal_1735}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1722 ( .a ({signal_3863, signal_3862, signal_1669}), .b ({signal_3999, signal_3998, signal_1737}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1723 ( .a ({signal_3871, signal_3870, signal_1673}), .b ({signal_4001, signal_4000, signal_1738}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1724 ( .a ({signal_3877, signal_3876, signal_1676}), .b ({signal_4003, signal_4002, signal_1739}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1726 ( .a ({signal_3881, signal_3880, signal_1678}), .b ({signal_4007, signal_4006, signal_1741}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1727 ( .a ({signal_3883, signal_3882, signal_1679}), .b ({signal_4009, signal_4008, signal_1742}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1728 ( .a ({signal_3885, signal_3884, signal_1680}), .b ({signal_4011, signal_4010, signal_1743}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1729 ( .a ({signal_3887, signal_3886, signal_1681}), .b ({signal_4013, signal_4012, signal_1744}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1730 ( .a ({signal_3889, signal_3888, signal_1682}), .b ({signal_4015, signal_4014, signal_1745}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1731 ( .a ({signal_3897, signal_3896, signal_1686}), .b ({signal_4017, signal_4016, signal_1746}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1732 ( .a ({signal_3903, signal_3902, signal_1689}), .b ({signal_4019, signal_4018, signal_1747}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1733 ( .a ({signal_3911, signal_3910, signal_1693}), .b ({signal_4021, signal_4020, signal_1748}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1734 ( .a ({signal_3917, signal_3916, signal_1696}), .b ({signal_4023, signal_4022, signal_1749}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1735 ( .a ({signal_3919, signal_3918, signal_1697}), .b ({signal_4025, signal_4024, signal_1750}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1736 ( .a ({signal_3923, signal_3922, signal_1699}), .b ({signal_4027, signal_4026, signal_1751}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1739 ( .a ({signal_3929, signal_3928, signal_1702}), .b ({signal_4033, signal_4032, signal_1754}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1745 ( .a ({signal_3941, signal_3940, signal_1708}), .b ({signal_4045, signal_4044, signal_1760}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1749 ( .a ({signal_3951, signal_3950, signal_1713}), .b ({signal_4053, signal_4052, signal_1764}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1751 ( .a ({signal_2729, signal_2728, signal_1102}), .b ({signal_3539, signal_3538, signal_1507}), .clk ( clk ), .r ({Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({signal_4057, signal_4056, signal_1766}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1753 ( .a ({signal_8282, signal_8278, signal_8274}), .b ({signal_3541, signal_3540, signal_1508}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287]}), .c ({signal_4061, signal_4060, signal_1768}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1754 ( .a ({signal_8210, signal_8208, signal_8206}), .b ({signal_3543, signal_3542, signal_1509}), .clk ( clk ), .r ({Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_4063, signal_4062, signal_1769}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1755 ( .a ({signal_2691, signal_2690, signal_1083}), .b ({signal_3545, signal_3544, signal_1510}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293]}), .c ({signal_4065, signal_4064, signal_1770}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1756 ( .a ({signal_8270, signal_8268, signal_8266}), .b ({signal_3539, signal_3538, signal_1507}), .clk ( clk ), .r ({Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({signal_4067, signal_4066, signal_1771}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1757 ( .a ({signal_2789, signal_2788, signal_1132}), .b ({signal_3547, signal_3546, signal_1511}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299]}), .c ({signal_4069, signal_4068, signal_1772}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1758 ( .a ({signal_8348, signal_8346, signal_8344}), .b ({signal_3547, signal_3546, signal_1511}), .clk ( clk ), .r ({Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({signal_4071, signal_4070, signal_1773}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1760 ( .a ({signal_8402, signal_8400, signal_8398}), .b ({signal_3553, signal_3552, signal_1514}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305]}), .c ({signal_4075, signal_4074, signal_1775}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1761 ( .a ({signal_8408, signal_8406, signal_8404}), .b ({signal_3555, signal_3554, signal_1515}), .clk ( clk ), .r ({Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({signal_4077, signal_4076, signal_1776}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1762 ( .a ({signal_8090, signal_8088, signal_8086}), .b ({signal_3557, signal_3556, signal_1516}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311]}), .c ({signal_4079, signal_4078, signal_1777}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1764 ( .a ({signal_8240, signal_8238, signal_8236}), .b ({signal_3563, signal_3562, signal_1519}), .clk ( clk ), .r ({Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({signal_4083, signal_4082, signal_1779}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1765 ( .a ({signal_8384, signal_8382, signal_8380}), .b ({signal_3565, signal_3564, signal_1520}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317]}), .c ({signal_4085, signal_4084, signal_1780}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1766 ( .a ({signal_8108, signal_8106, signal_8104}), .b ({signal_3567, signal_3566, signal_1521}), .clk ( clk ), .r ({Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_4087, signal_4086, signal_1781}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1767 ( .a ({signal_8168, signal_8166, signal_8164}), .b ({signal_3569, signal_3568, signal_1522}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323]}), .c ({signal_4089, signal_4088, signal_1782}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1769 ( .a ({signal_2681, signal_2680, signal_1078}), .b ({signal_3569, signal_3568, signal_1522}), .clk ( clk ), .r ({Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({signal_4093, signal_4092, signal_1784}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1770 ( .a ({signal_2695, signal_2694, signal_1085}), .b ({signal_3581, signal_3580, signal_1528}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329]}), .c ({signal_4095, signal_4094, signal_1785}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1772 ( .a ({signal_8138, signal_8136, signal_8134}), .b ({signal_3567, signal_3566, signal_1521}), .clk ( clk ), .r ({Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({signal_4099, signal_4098, signal_1787}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1773 ( .a ({signal_2831, signal_2830, signal_1153}), .b ({signal_3595, signal_3594, signal_1535}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335]}), .c ({signal_4101, signal_4100, signal_1788}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1776 ( .a ({signal_8312, signal_8310, signal_8308}), .b ({signal_3565, signal_3564, signal_1520}), .clk ( clk ), .r ({Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({signal_4107, signal_4106, signal_1791}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1778 ( .a ({signal_8414, signal_8412, signal_8410}), .b ({signal_3619, signal_3618, signal_1547}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341]}), .c ({signal_4111, signal_4110, signal_1793}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1779 ( .a ({signal_2697, signal_2696, signal_1086}), .b ({signal_3621, signal_3620, signal_1548}), .clk ( clk ), .r ({Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({signal_4113, signal_4112, signal_1794}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1782 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_3631, signal_3630, signal_1553}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347]}), .c ({signal_4119, signal_4118, signal_1797}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1783 ( .a ({signal_8102, signal_8100, signal_8098}), .b ({signal_3633, signal_3632, signal_1554}), .clk ( clk ), .r ({Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_4121, signal_4120, signal_1798}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1784 ( .a ({signal_2689, signal_2688, signal_1082}), .b ({signal_3555, signal_3554, signal_1515}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353]}), .c ({signal_4123, signal_4122, signal_1799}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1785 ( .a ({signal_8300, signal_8298, signal_8296}), .b ({signal_3641, signal_3640, signal_1558}), .clk ( clk ), .r ({Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({signal_4125, signal_4124, signal_1800}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1786 ( .a ({signal_8228, signal_8226, signal_8224}), .b ({signal_3643, signal_3642, signal_1559}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359]}), .c ({signal_4127, signal_4126, signal_1801}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1835 ( .a ({signal_4057, signal_4056, signal_1766}), .b ({signal_4225, signal_4224, signal_1850}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1836 ( .a ({signal_4065, signal_4064, signal_1770}), .b ({signal_4227, signal_4226, signal_1851}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1837 ( .a ({signal_4069, signal_4068, signal_1772}), .b ({signal_4229, signal_4228, signal_1852}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1838 ( .a ({signal_4071, signal_4070, signal_1773}), .b ({signal_4231, signal_4230, signal_1853}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1839 ( .a ({signal_4075, signal_4074, signal_1775}), .b ({signal_4233, signal_4232, signal_1854}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1840 ( .a ({signal_4077, signal_4076, signal_1776}), .b ({signal_4235, signal_4234, signal_1855}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1841 ( .a ({signal_4079, signal_4078, signal_1777}), .b ({signal_4237, signal_4236, signal_1856}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1843 ( .a ({signal_4083, signal_4082, signal_1779}), .b ({signal_4241, signal_4240, signal_1858}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1844 ( .a ({signal_4085, signal_4084, signal_1780}), .b ({signal_4243, signal_4242, signal_1859}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1845 ( .a ({signal_4087, signal_4086, signal_1781}), .b ({signal_4245, signal_4244, signal_1860}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1846 ( .a ({signal_4093, signal_4092, signal_1784}), .b ({signal_4247, signal_4246, signal_1861}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1847 ( .a ({signal_4095, signal_4094, signal_1785}), .b ({signal_4249, signal_4248, signal_1862}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1848 ( .a ({signal_4099, signal_4098, signal_1787}), .b ({signal_4251, signal_4250, signal_1863}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1849 ( .a ({signal_4101, signal_4100, signal_1788}), .b ({signal_4253, signal_4252, signal_1864}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1850 ( .a ({signal_4107, signal_4106, signal_1791}), .b ({signal_4255, signal_4254, signal_1865}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1851 ( .a ({signal_4111, signal_4110, signal_1793}), .b ({signal_4257, signal_4256, signal_1866}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1852 ( .a ({signal_4113, signal_4112, signal_1794}), .b ({signal_4259, signal_4258, signal_1867}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1854 ( .a ({signal_4119, signal_4118, signal_1797}), .b ({signal_4263, signal_4262, signal_1869}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1855 ( .a ({signal_4121, signal_4120, signal_1798}), .b ({signal_4265, signal_4264, signal_1870}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1856 ( .a ({signal_4123, signal_4122, signal_1799}), .b ({signal_4267, signal_4266, signal_1871}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1857 ( .a ({signal_4125, signal_4124, signal_1800}), .b ({signal_4269, signal_4268, signal_1872}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1858 ( .a ({signal_4127, signal_4126, signal_1801}), .b ({signal_4271, signal_4270, signal_1873}) ) ;
    buf_clk cell_2824 ( .C ( clk ), .D ( signal_8415 ), .Q ( signal_8416 ) ) ;
    buf_clk cell_2826 ( .C ( clk ), .D ( signal_8417 ), .Q ( signal_8418 ) ) ;
    buf_clk cell_2828 ( .C ( clk ), .D ( signal_8419 ), .Q ( signal_8420 ) ) ;
    buf_clk cell_2830 ( .C ( clk ), .D ( signal_8421 ), .Q ( signal_8422 ) ) ;
    buf_clk cell_2832 ( .C ( clk ), .D ( signal_8423 ), .Q ( signal_8424 ) ) ;
    buf_clk cell_2834 ( .C ( clk ), .D ( signal_8425 ), .Q ( signal_8426 ) ) ;
    buf_clk cell_2836 ( .C ( clk ), .D ( signal_8427 ), .Q ( signal_8428 ) ) ;
    buf_clk cell_2838 ( .C ( clk ), .D ( signal_8429 ), .Q ( signal_8430 ) ) ;
    buf_clk cell_2840 ( .C ( clk ), .D ( signal_8431 ), .Q ( signal_8432 ) ) ;
    buf_clk cell_2842 ( .C ( clk ), .D ( signal_8433 ), .Q ( signal_8434 ) ) ;
    buf_clk cell_2844 ( .C ( clk ), .D ( signal_8435 ), .Q ( signal_8436 ) ) ;
    buf_clk cell_2846 ( .C ( clk ), .D ( signal_8437 ), .Q ( signal_8438 ) ) ;
    buf_clk cell_2848 ( .C ( clk ), .D ( signal_8439 ), .Q ( signal_8440 ) ) ;
    buf_clk cell_2850 ( .C ( clk ), .D ( signal_8441 ), .Q ( signal_8442 ) ) ;
    buf_clk cell_2852 ( .C ( clk ), .D ( signal_8443 ), .Q ( signal_8444 ) ) ;
    buf_clk cell_2854 ( .C ( clk ), .D ( signal_8445 ), .Q ( signal_8446 ) ) ;
    buf_clk cell_2856 ( .C ( clk ), .D ( signal_8447 ), .Q ( signal_8448 ) ) ;
    buf_clk cell_2858 ( .C ( clk ), .D ( signal_8449 ), .Q ( signal_8450 ) ) ;
    buf_clk cell_2860 ( .C ( clk ), .D ( signal_8451 ), .Q ( signal_8452 ) ) ;
    buf_clk cell_2862 ( .C ( clk ), .D ( signal_8453 ), .Q ( signal_8454 ) ) ;
    buf_clk cell_2864 ( .C ( clk ), .D ( signal_8455 ), .Q ( signal_8456 ) ) ;
    buf_clk cell_2866 ( .C ( clk ), .D ( signal_8457 ), .Q ( signal_8458 ) ) ;
    buf_clk cell_2868 ( .C ( clk ), .D ( signal_8459 ), .Q ( signal_8460 ) ) ;
    buf_clk cell_2870 ( .C ( clk ), .D ( signal_8461 ), .Q ( signal_8462 ) ) ;
    buf_clk cell_2872 ( .C ( clk ), .D ( signal_8463 ), .Q ( signal_8464 ) ) ;
    buf_clk cell_2874 ( .C ( clk ), .D ( signal_8465 ), .Q ( signal_8466 ) ) ;
    buf_clk cell_2876 ( .C ( clk ), .D ( signal_8467 ), .Q ( signal_8468 ) ) ;
    buf_clk cell_2878 ( .C ( clk ), .D ( signal_8469 ), .Q ( signal_8470 ) ) ;
    buf_clk cell_2880 ( .C ( clk ), .D ( signal_8471 ), .Q ( signal_8472 ) ) ;
    buf_clk cell_2882 ( .C ( clk ), .D ( signal_8473 ), .Q ( signal_8474 ) ) ;
    buf_clk cell_2884 ( .C ( clk ), .D ( signal_8475 ), .Q ( signal_8476 ) ) ;
    buf_clk cell_2886 ( .C ( clk ), .D ( signal_8477 ), .Q ( signal_8478 ) ) ;
    buf_clk cell_2888 ( .C ( clk ), .D ( signal_8479 ), .Q ( signal_8480 ) ) ;
    buf_clk cell_2894 ( .C ( clk ), .D ( signal_8485 ), .Q ( signal_8486 ) ) ;
    buf_clk cell_2900 ( .C ( clk ), .D ( signal_8491 ), .Q ( signal_8492 ) ) ;
    buf_clk cell_2906 ( .C ( clk ), .D ( signal_8497 ), .Q ( signal_8498 ) ) ;
    buf_clk cell_2908 ( .C ( clk ), .D ( signal_8499 ), .Q ( signal_8500 ) ) ;
    buf_clk cell_2910 ( .C ( clk ), .D ( signal_8501 ), .Q ( signal_8502 ) ) ;
    buf_clk cell_2912 ( .C ( clk ), .D ( signal_8503 ), .Q ( signal_8504 ) ) ;
    buf_clk cell_2914 ( .C ( clk ), .D ( signal_8505 ), .Q ( signal_8506 ) ) ;
    buf_clk cell_2916 ( .C ( clk ), .D ( signal_8507 ), .Q ( signal_8508 ) ) ;
    buf_clk cell_2918 ( .C ( clk ), .D ( signal_8509 ), .Q ( signal_8510 ) ) ;
    buf_clk cell_2920 ( .C ( clk ), .D ( signal_8511 ), .Q ( signal_8512 ) ) ;
    buf_clk cell_2922 ( .C ( clk ), .D ( signal_8513 ), .Q ( signal_8514 ) ) ;
    buf_clk cell_2924 ( .C ( clk ), .D ( signal_8515 ), .Q ( signal_8516 ) ) ;
    buf_clk cell_2926 ( .C ( clk ), .D ( signal_8517 ), .Q ( signal_8518 ) ) ;
    buf_clk cell_2928 ( .C ( clk ), .D ( signal_8519 ), .Q ( signal_8520 ) ) ;
    buf_clk cell_2930 ( .C ( clk ), .D ( signal_8521 ), .Q ( signal_8522 ) ) ;
    buf_clk cell_2932 ( .C ( clk ), .D ( signal_8523 ), .Q ( signal_8524 ) ) ;
    buf_clk cell_2934 ( .C ( clk ), .D ( signal_8525 ), .Q ( signal_8526 ) ) ;
    buf_clk cell_2936 ( .C ( clk ), .D ( signal_8527 ), .Q ( signal_8528 ) ) ;
    buf_clk cell_2938 ( .C ( clk ), .D ( signal_8529 ), .Q ( signal_8530 ) ) ;
    buf_clk cell_2940 ( .C ( clk ), .D ( signal_8531 ), .Q ( signal_8532 ) ) ;
    buf_clk cell_2942 ( .C ( clk ), .D ( signal_8533 ), .Q ( signal_8534 ) ) ;
    buf_clk cell_2944 ( .C ( clk ), .D ( signal_8535 ), .Q ( signal_8536 ) ) ;
    buf_clk cell_2946 ( .C ( clk ), .D ( signal_8537 ), .Q ( signal_8538 ) ) ;
    buf_clk cell_2948 ( .C ( clk ), .D ( signal_8539 ), .Q ( signal_8540 ) ) ;
    buf_clk cell_2950 ( .C ( clk ), .D ( signal_8541 ), .Q ( signal_8542 ) ) ;
    buf_clk cell_2952 ( .C ( clk ), .D ( signal_8543 ), .Q ( signal_8544 ) ) ;
    buf_clk cell_2954 ( .C ( clk ), .D ( signal_8545 ), .Q ( signal_8546 ) ) ;
    buf_clk cell_2956 ( .C ( clk ), .D ( signal_8547 ), .Q ( signal_8548 ) ) ;
    buf_clk cell_2958 ( .C ( clk ), .D ( signal_8549 ), .Q ( signal_8550 ) ) ;
    buf_clk cell_2960 ( .C ( clk ), .D ( signal_8551 ), .Q ( signal_8552 ) ) ;
    buf_clk cell_2962 ( .C ( clk ), .D ( signal_8553 ), .Q ( signal_8554 ) ) ;
    buf_clk cell_2964 ( .C ( clk ), .D ( signal_8555 ), .Q ( signal_8556 ) ) ;
    buf_clk cell_2966 ( .C ( clk ), .D ( signal_8557 ), .Q ( signal_8558 ) ) ;
    buf_clk cell_2968 ( .C ( clk ), .D ( signal_8559 ), .Q ( signal_8560 ) ) ;
    buf_clk cell_2970 ( .C ( clk ), .D ( signal_8561 ), .Q ( signal_8562 ) ) ;
    buf_clk cell_2972 ( .C ( clk ), .D ( signal_8563 ), .Q ( signal_8564 ) ) ;
    buf_clk cell_2974 ( .C ( clk ), .D ( signal_8565 ), .Q ( signal_8566 ) ) ;
    buf_clk cell_2976 ( .C ( clk ), .D ( signal_8567 ), .Q ( signal_8568 ) ) ;
    buf_clk cell_2978 ( .C ( clk ), .D ( signal_8569 ), .Q ( signal_8570 ) ) ;
    buf_clk cell_2980 ( .C ( clk ), .D ( signal_8571 ), .Q ( signal_8572 ) ) ;
    buf_clk cell_2982 ( .C ( clk ), .D ( signal_8573 ), .Q ( signal_8574 ) ) ;
    buf_clk cell_2984 ( .C ( clk ), .D ( signal_8575 ), .Q ( signal_8576 ) ) ;
    buf_clk cell_2986 ( .C ( clk ), .D ( signal_8577 ), .Q ( signal_8578 ) ) ;
    buf_clk cell_2988 ( .C ( clk ), .D ( signal_8579 ), .Q ( signal_8580 ) ) ;
    buf_clk cell_2990 ( .C ( clk ), .D ( signal_8581 ), .Q ( signal_8582 ) ) ;
    buf_clk cell_2992 ( .C ( clk ), .D ( signal_8583 ), .Q ( signal_8584 ) ) ;
    buf_clk cell_2994 ( .C ( clk ), .D ( signal_8585 ), .Q ( signal_8586 ) ) ;
    buf_clk cell_2996 ( .C ( clk ), .D ( signal_8587 ), .Q ( signal_8588 ) ) ;
    buf_clk cell_2998 ( .C ( clk ), .D ( signal_8589 ), .Q ( signal_8590 ) ) ;
    buf_clk cell_3000 ( .C ( clk ), .D ( signal_8591 ), .Q ( signal_8592 ) ) ;
    buf_clk cell_3002 ( .C ( clk ), .D ( signal_8593 ), .Q ( signal_8594 ) ) ;
    buf_clk cell_3004 ( .C ( clk ), .D ( signal_8595 ), .Q ( signal_8596 ) ) ;
    buf_clk cell_3006 ( .C ( clk ), .D ( signal_8597 ), .Q ( signal_8598 ) ) ;
    buf_clk cell_3008 ( .C ( clk ), .D ( signal_8599 ), .Q ( signal_8600 ) ) ;
    buf_clk cell_3010 ( .C ( clk ), .D ( signal_8601 ), .Q ( signal_8602 ) ) ;
    buf_clk cell_3012 ( .C ( clk ), .D ( signal_8603 ), .Q ( signal_8604 ) ) ;
    buf_clk cell_3014 ( .C ( clk ), .D ( signal_8605 ), .Q ( signal_8606 ) ) ;
    buf_clk cell_3016 ( .C ( clk ), .D ( signal_8607 ), .Q ( signal_8608 ) ) ;
    buf_clk cell_3018 ( .C ( clk ), .D ( signal_8609 ), .Q ( signal_8610 ) ) ;
    buf_clk cell_3020 ( .C ( clk ), .D ( signal_8611 ), .Q ( signal_8612 ) ) ;
    buf_clk cell_3022 ( .C ( clk ), .D ( signal_8613 ), .Q ( signal_8614 ) ) ;
    buf_clk cell_3024 ( .C ( clk ), .D ( signal_8615 ), .Q ( signal_8616 ) ) ;
    buf_clk cell_3026 ( .C ( clk ), .D ( signal_8617 ), .Q ( signal_8618 ) ) ;
    buf_clk cell_3030 ( .C ( clk ), .D ( signal_8621 ), .Q ( signal_8622 ) ) ;
    buf_clk cell_3034 ( .C ( clk ), .D ( signal_8625 ), .Q ( signal_8626 ) ) ;
    buf_clk cell_3038 ( .C ( clk ), .D ( signal_8629 ), .Q ( signal_8630 ) ) ;
    buf_clk cell_3040 ( .C ( clk ), .D ( signal_8631 ), .Q ( signal_8632 ) ) ;
    buf_clk cell_3042 ( .C ( clk ), .D ( signal_8633 ), .Q ( signal_8634 ) ) ;
    buf_clk cell_3044 ( .C ( clk ), .D ( signal_8635 ), .Q ( signal_8636 ) ) ;
    buf_clk cell_3046 ( .C ( clk ), .D ( signal_8637 ), .Q ( signal_8638 ) ) ;
    buf_clk cell_3048 ( .C ( clk ), .D ( signal_8639 ), .Q ( signal_8640 ) ) ;
    buf_clk cell_3050 ( .C ( clk ), .D ( signal_8641 ), .Q ( signal_8642 ) ) ;
    buf_clk cell_3054 ( .C ( clk ), .D ( signal_8645 ), .Q ( signal_8646 ) ) ;
    buf_clk cell_3058 ( .C ( clk ), .D ( signal_8649 ), .Q ( signal_8650 ) ) ;
    buf_clk cell_3062 ( .C ( clk ), .D ( signal_8653 ), .Q ( signal_8654 ) ) ;
    buf_clk cell_3064 ( .C ( clk ), .D ( signal_8655 ), .Q ( signal_8656 ) ) ;
    buf_clk cell_3066 ( .C ( clk ), .D ( signal_8657 ), .Q ( signal_8658 ) ) ;
    buf_clk cell_3068 ( .C ( clk ), .D ( signal_8659 ), .Q ( signal_8660 ) ) ;
    buf_clk cell_3070 ( .C ( clk ), .D ( signal_8661 ), .Q ( signal_8662 ) ) ;
    buf_clk cell_3072 ( .C ( clk ), .D ( signal_8663 ), .Q ( signal_8664 ) ) ;
    buf_clk cell_3074 ( .C ( clk ), .D ( signal_8665 ), .Q ( signal_8666 ) ) ;
    buf_clk cell_3076 ( .C ( clk ), .D ( signal_8667 ), .Q ( signal_8668 ) ) ;
    buf_clk cell_3078 ( .C ( clk ), .D ( signal_8669 ), .Q ( signal_8670 ) ) ;
    buf_clk cell_3080 ( .C ( clk ), .D ( signal_8671 ), .Q ( signal_8672 ) ) ;
    buf_clk cell_3082 ( .C ( clk ), .D ( signal_8673 ), .Q ( signal_8674 ) ) ;
    buf_clk cell_3084 ( .C ( clk ), .D ( signal_8675 ), .Q ( signal_8676 ) ) ;
    buf_clk cell_3086 ( .C ( clk ), .D ( signal_8677 ), .Q ( signal_8678 ) ) ;
    buf_clk cell_3088 ( .C ( clk ), .D ( signal_8679 ), .Q ( signal_8680 ) ) ;
    buf_clk cell_3090 ( .C ( clk ), .D ( signal_8681 ), .Q ( signal_8682 ) ) ;
    buf_clk cell_3092 ( .C ( clk ), .D ( signal_8683 ), .Q ( signal_8684 ) ) ;
    buf_clk cell_3094 ( .C ( clk ), .D ( signal_8685 ), .Q ( signal_8686 ) ) ;
    buf_clk cell_3096 ( .C ( clk ), .D ( signal_8687 ), .Q ( signal_8688 ) ) ;
    buf_clk cell_3098 ( .C ( clk ), .D ( signal_8689 ), .Q ( signal_8690 ) ) ;
    buf_clk cell_3100 ( .C ( clk ), .D ( signal_8691 ), .Q ( signal_8692 ) ) ;
    buf_clk cell_3102 ( .C ( clk ), .D ( signal_8693 ), .Q ( signal_8694 ) ) ;
    buf_clk cell_3104 ( .C ( clk ), .D ( signal_8695 ), .Q ( signal_8696 ) ) ;
    buf_clk cell_3106 ( .C ( clk ), .D ( signal_8697 ), .Q ( signal_8698 ) ) ;
    buf_clk cell_3108 ( .C ( clk ), .D ( signal_8699 ), .Q ( signal_8700 ) ) ;
    buf_clk cell_3110 ( .C ( clk ), .D ( signal_8701 ), .Q ( signal_8702 ) ) ;
    buf_clk cell_3112 ( .C ( clk ), .D ( signal_8703 ), .Q ( signal_8704 ) ) ;
    buf_clk cell_3114 ( .C ( clk ), .D ( signal_8705 ), .Q ( signal_8706 ) ) ;
    buf_clk cell_3116 ( .C ( clk ), .D ( signal_8707 ), .Q ( signal_8708 ) ) ;
    buf_clk cell_3118 ( .C ( clk ), .D ( signal_8709 ), .Q ( signal_8710 ) ) ;
    buf_clk cell_3120 ( .C ( clk ), .D ( signal_8711 ), .Q ( signal_8712 ) ) ;
    buf_clk cell_3122 ( .C ( clk ), .D ( signal_8713 ), .Q ( signal_8714 ) ) ;
    buf_clk cell_3124 ( .C ( clk ), .D ( signal_8715 ), .Q ( signal_8716 ) ) ;
    buf_clk cell_3126 ( .C ( clk ), .D ( signal_8717 ), .Q ( signal_8718 ) ) ;
    buf_clk cell_3128 ( .C ( clk ), .D ( signal_8719 ), .Q ( signal_8720 ) ) ;
    buf_clk cell_3132 ( .C ( clk ), .D ( signal_8723 ), .Q ( signal_8724 ) ) ;
    buf_clk cell_3136 ( .C ( clk ), .D ( signal_8727 ), .Q ( signal_8728 ) ) ;
    buf_clk cell_3140 ( .C ( clk ), .D ( signal_8731 ), .Q ( signal_8732 ) ) ;
    buf_clk cell_3142 ( .C ( clk ), .D ( signal_8733 ), .Q ( signal_8734 ) ) ;
    buf_clk cell_3144 ( .C ( clk ), .D ( signal_8735 ), .Q ( signal_8736 ) ) ;
    buf_clk cell_3146 ( .C ( clk ), .D ( signal_8737 ), .Q ( signal_8738 ) ) ;
    buf_clk cell_3150 ( .C ( clk ), .D ( signal_8741 ), .Q ( signal_8742 ) ) ;
    buf_clk cell_3154 ( .C ( clk ), .D ( signal_8745 ), .Q ( signal_8746 ) ) ;
    buf_clk cell_3158 ( .C ( clk ), .D ( signal_8749 ), .Q ( signal_8750 ) ) ;
    buf_clk cell_3160 ( .C ( clk ), .D ( signal_8751 ), .Q ( signal_8752 ) ) ;
    buf_clk cell_3162 ( .C ( clk ), .D ( signal_8753 ), .Q ( signal_8754 ) ) ;
    buf_clk cell_3164 ( .C ( clk ), .D ( signal_8755 ), .Q ( signal_8756 ) ) ;
    buf_clk cell_3166 ( .C ( clk ), .D ( signal_8757 ), .Q ( signal_8758 ) ) ;
    buf_clk cell_3168 ( .C ( clk ), .D ( signal_8759 ), .Q ( signal_8760 ) ) ;
    buf_clk cell_3170 ( .C ( clk ), .D ( signal_8761 ), .Q ( signal_8762 ) ) ;
    buf_clk cell_3172 ( .C ( clk ), .D ( signal_8763 ), .Q ( signal_8764 ) ) ;
    buf_clk cell_3174 ( .C ( clk ), .D ( signal_8765 ), .Q ( signal_8766 ) ) ;
    buf_clk cell_3176 ( .C ( clk ), .D ( signal_8767 ), .Q ( signal_8768 ) ) ;
    buf_clk cell_3182 ( .C ( clk ), .D ( signal_8773 ), .Q ( signal_8774 ) ) ;
    buf_clk cell_3188 ( .C ( clk ), .D ( signal_8779 ), .Q ( signal_8780 ) ) ;
    buf_clk cell_3194 ( .C ( clk ), .D ( signal_8785 ), .Q ( signal_8786 ) ) ;
    buf_clk cell_3196 ( .C ( clk ), .D ( signal_8787 ), .Q ( signal_8788 ) ) ;
    buf_clk cell_3198 ( .C ( clk ), .D ( signal_8789 ), .Q ( signal_8790 ) ) ;
    buf_clk cell_3200 ( .C ( clk ), .D ( signal_8791 ), .Q ( signal_8792 ) ) ;
    buf_clk cell_3202 ( .C ( clk ), .D ( signal_8793 ), .Q ( signal_8794 ) ) ;
    buf_clk cell_3204 ( .C ( clk ), .D ( signal_8795 ), .Q ( signal_8796 ) ) ;
    buf_clk cell_3206 ( .C ( clk ), .D ( signal_8797 ), .Q ( signal_8798 ) ) ;
    buf_clk cell_3208 ( .C ( clk ), .D ( signal_8799 ), .Q ( signal_8800 ) ) ;
    buf_clk cell_3210 ( .C ( clk ), .D ( signal_8801 ), .Q ( signal_8802 ) ) ;
    buf_clk cell_3212 ( .C ( clk ), .D ( signal_8803 ), .Q ( signal_8804 ) ) ;
    buf_clk cell_3214 ( .C ( clk ), .D ( signal_8805 ), .Q ( signal_8806 ) ) ;
    buf_clk cell_3216 ( .C ( clk ), .D ( signal_8807 ), .Q ( signal_8808 ) ) ;
    buf_clk cell_3218 ( .C ( clk ), .D ( signal_8809 ), .Q ( signal_8810 ) ) ;
    buf_clk cell_3222 ( .C ( clk ), .D ( signal_8813 ), .Q ( signal_8814 ) ) ;
    buf_clk cell_3226 ( .C ( clk ), .D ( signal_8817 ), .Q ( signal_8818 ) ) ;
    buf_clk cell_3230 ( .C ( clk ), .D ( signal_8821 ), .Q ( signal_8822 ) ) ;
    buf_clk cell_3232 ( .C ( clk ), .D ( signal_8823 ), .Q ( signal_8824 ) ) ;
    buf_clk cell_3234 ( .C ( clk ), .D ( signal_8825 ), .Q ( signal_8826 ) ) ;
    buf_clk cell_3236 ( .C ( clk ), .D ( signal_8827 ), .Q ( signal_8828 ) ) ;
    buf_clk cell_3238 ( .C ( clk ), .D ( signal_8829 ), .Q ( signal_8830 ) ) ;
    buf_clk cell_3240 ( .C ( clk ), .D ( signal_8831 ), .Q ( signal_8832 ) ) ;
    buf_clk cell_3242 ( .C ( clk ), .D ( signal_8833 ), .Q ( signal_8834 ) ) ;
    buf_clk cell_3244 ( .C ( clk ), .D ( signal_8835 ), .Q ( signal_8836 ) ) ;
    buf_clk cell_3246 ( .C ( clk ), .D ( signal_8837 ), .Q ( signal_8838 ) ) ;
    buf_clk cell_3248 ( .C ( clk ), .D ( signal_8839 ), .Q ( signal_8840 ) ) ;
    buf_clk cell_3250 ( .C ( clk ), .D ( signal_8841 ), .Q ( signal_8842 ) ) ;
    buf_clk cell_3252 ( .C ( clk ), .D ( signal_8843 ), .Q ( signal_8844 ) ) ;
    buf_clk cell_3254 ( .C ( clk ), .D ( signal_8845 ), .Q ( signal_8846 ) ) ;
    buf_clk cell_3256 ( .C ( clk ), .D ( signal_8847 ), .Q ( signal_8848 ) ) ;
    buf_clk cell_3258 ( .C ( clk ), .D ( signal_8849 ), .Q ( signal_8850 ) ) ;
    buf_clk cell_3260 ( .C ( clk ), .D ( signal_8851 ), .Q ( signal_8852 ) ) ;
    buf_clk cell_3262 ( .C ( clk ), .D ( signal_8853 ), .Q ( signal_8854 ) ) ;
    buf_clk cell_3264 ( .C ( clk ), .D ( signal_8855 ), .Q ( signal_8856 ) ) ;
    buf_clk cell_3266 ( .C ( clk ), .D ( signal_8857 ), .Q ( signal_8858 ) ) ;
    buf_clk cell_3268 ( .C ( clk ), .D ( signal_8859 ), .Q ( signal_8860 ) ) ;
    buf_clk cell_3270 ( .C ( clk ), .D ( signal_8861 ), .Q ( signal_8862 ) ) ;
    buf_clk cell_3272 ( .C ( clk ), .D ( signal_8863 ), .Q ( signal_8864 ) ) ;
    buf_clk cell_3274 ( .C ( clk ), .D ( signal_8865 ), .Q ( signal_8866 ) ) ;
    buf_clk cell_3276 ( .C ( clk ), .D ( signal_8867 ), .Q ( signal_8868 ) ) ;
    buf_clk cell_3278 ( .C ( clk ), .D ( signal_8869 ), .Q ( signal_8870 ) ) ;
    buf_clk cell_3280 ( .C ( clk ), .D ( signal_8871 ), .Q ( signal_8872 ) ) ;
    buf_clk cell_3282 ( .C ( clk ), .D ( signal_8873 ), .Q ( signal_8874 ) ) ;
    buf_clk cell_3284 ( .C ( clk ), .D ( signal_8875 ), .Q ( signal_8876 ) ) ;
    buf_clk cell_3288 ( .C ( clk ), .D ( signal_8879 ), .Q ( signal_8880 ) ) ;
    buf_clk cell_3292 ( .C ( clk ), .D ( signal_8883 ), .Q ( signal_8884 ) ) ;
    buf_clk cell_3296 ( .C ( clk ), .D ( signal_8887 ), .Q ( signal_8888 ) ) ;
    buf_clk cell_3298 ( .C ( clk ), .D ( signal_8889 ), .Q ( signal_8890 ) ) ;
    buf_clk cell_3300 ( .C ( clk ), .D ( signal_8891 ), .Q ( signal_8892 ) ) ;
    buf_clk cell_3302 ( .C ( clk ), .D ( signal_8893 ), .Q ( signal_8894 ) ) ;
    buf_clk cell_3304 ( .C ( clk ), .D ( signal_8895 ), .Q ( signal_8896 ) ) ;
    buf_clk cell_3306 ( .C ( clk ), .D ( signal_8897 ), .Q ( signal_8898 ) ) ;
    buf_clk cell_3308 ( .C ( clk ), .D ( signal_8899 ), .Q ( signal_8900 ) ) ;
    buf_clk cell_3310 ( .C ( clk ), .D ( signal_8901 ), .Q ( signal_8902 ) ) ;
    buf_clk cell_3312 ( .C ( clk ), .D ( signal_8903 ), .Q ( signal_8904 ) ) ;
    buf_clk cell_3314 ( .C ( clk ), .D ( signal_8905 ), .Q ( signal_8906 ) ) ;
    buf_clk cell_3316 ( .C ( clk ), .D ( signal_8907 ), .Q ( signal_8908 ) ) ;
    buf_clk cell_3318 ( .C ( clk ), .D ( signal_8909 ), .Q ( signal_8910 ) ) ;
    buf_clk cell_3320 ( .C ( clk ), .D ( signal_8911 ), .Q ( signal_8912 ) ) ;
    buf_clk cell_3322 ( .C ( clk ), .D ( signal_8913 ), .Q ( signal_8914 ) ) ;
    buf_clk cell_3324 ( .C ( clk ), .D ( signal_8915 ), .Q ( signal_8916 ) ) ;
    buf_clk cell_3326 ( .C ( clk ), .D ( signal_8917 ), .Q ( signal_8918 ) ) ;
    buf_clk cell_3328 ( .C ( clk ), .D ( signal_8919 ), .Q ( signal_8920 ) ) ;
    buf_clk cell_3330 ( .C ( clk ), .D ( signal_8921 ), .Q ( signal_8922 ) ) ;
    buf_clk cell_3332 ( .C ( clk ), .D ( signal_8923 ), .Q ( signal_8924 ) ) ;
    buf_clk cell_3346 ( .C ( clk ), .D ( signal_8937 ), .Q ( signal_8938 ) ) ;
    buf_clk cell_3350 ( .C ( clk ), .D ( signal_8941 ), .Q ( signal_8942 ) ) ;
    buf_clk cell_3354 ( .C ( clk ), .D ( signal_8945 ), .Q ( signal_8946 ) ) ;
    buf_clk cell_3364 ( .C ( clk ), .D ( signal_8955 ), .Q ( signal_8956 ) ) ;
    buf_clk cell_3368 ( .C ( clk ), .D ( signal_8959 ), .Q ( signal_8960 ) ) ;
    buf_clk cell_3372 ( .C ( clk ), .D ( signal_8963 ), .Q ( signal_8964 ) ) ;
    buf_clk cell_3376 ( .C ( clk ), .D ( signal_8967 ), .Q ( signal_8968 ) ) ;
    buf_clk cell_3380 ( .C ( clk ), .D ( signal_8971 ), .Q ( signal_8972 ) ) ;
    buf_clk cell_3384 ( .C ( clk ), .D ( signal_8975 ), .Q ( signal_8976 ) ) ;
    buf_clk cell_3388 ( .C ( clk ), .D ( signal_8979 ), .Q ( signal_8980 ) ) ;
    buf_clk cell_3392 ( .C ( clk ), .D ( signal_8983 ), .Q ( signal_8984 ) ) ;
    buf_clk cell_3396 ( .C ( clk ), .D ( signal_8987 ), .Q ( signal_8988 ) ) ;
    buf_clk cell_3404 ( .C ( clk ), .D ( signal_8995 ), .Q ( signal_8996 ) ) ;
    buf_clk cell_3412 ( .C ( clk ), .D ( signal_9003 ), .Q ( signal_9004 ) ) ;
    buf_clk cell_3420 ( .C ( clk ), .D ( signal_9011 ), .Q ( signal_9012 ) ) ;
    buf_clk cell_3436 ( .C ( clk ), .D ( signal_9027 ), .Q ( signal_9028 ) ) ;
    buf_clk cell_3440 ( .C ( clk ), .D ( signal_9031 ), .Q ( signal_9032 ) ) ;
    buf_clk cell_3444 ( .C ( clk ), .D ( signal_9035 ), .Q ( signal_9036 ) ) ;
    buf_clk cell_3460 ( .C ( clk ), .D ( signal_9051 ), .Q ( signal_9052 ) ) ;
    buf_clk cell_3464 ( .C ( clk ), .D ( signal_9055 ), .Q ( signal_9056 ) ) ;
    buf_clk cell_3468 ( .C ( clk ), .D ( signal_9059 ), .Q ( signal_9060 ) ) ;
    buf_clk cell_3502 ( .C ( clk ), .D ( signal_9093 ), .Q ( signal_9094 ) ) ;
    buf_clk cell_3506 ( .C ( clk ), .D ( signal_9097 ), .Q ( signal_9098 ) ) ;
    buf_clk cell_3510 ( .C ( clk ), .D ( signal_9101 ), .Q ( signal_9102 ) ) ;
    buf_clk cell_3538 ( .C ( clk ), .D ( signal_9129 ), .Q ( signal_9130 ) ) ;
    buf_clk cell_3542 ( .C ( clk ), .D ( signal_9133 ), .Q ( signal_9134 ) ) ;
    buf_clk cell_3546 ( .C ( clk ), .D ( signal_9137 ), .Q ( signal_9138 ) ) ;
    buf_clk cell_3562 ( .C ( clk ), .D ( signal_9153 ), .Q ( signal_9154 ) ) ;
    buf_clk cell_3566 ( .C ( clk ), .D ( signal_9157 ), .Q ( signal_9158 ) ) ;
    buf_clk cell_3570 ( .C ( clk ), .D ( signal_9161 ), .Q ( signal_9162 ) ) ;
    buf_clk cell_3574 ( .C ( clk ), .D ( signal_9165 ), .Q ( signal_9166 ) ) ;
    buf_clk cell_3578 ( .C ( clk ), .D ( signal_9169 ), .Q ( signal_9170 ) ) ;
    buf_clk cell_3582 ( .C ( clk ), .D ( signal_9173 ), .Q ( signal_9174 ) ) ;
    buf_clk cell_3586 ( .C ( clk ), .D ( signal_9177 ), .Q ( signal_9178 ) ) ;
    buf_clk cell_3590 ( .C ( clk ), .D ( signal_9181 ), .Q ( signal_9182 ) ) ;
    buf_clk cell_3594 ( .C ( clk ), .D ( signal_9185 ), .Q ( signal_9186 ) ) ;
    buf_clk cell_3598 ( .C ( clk ), .D ( signal_9189 ), .Q ( signal_9190 ) ) ;
    buf_clk cell_3602 ( .C ( clk ), .D ( signal_9193 ), .Q ( signal_9194 ) ) ;
    buf_clk cell_3606 ( .C ( clk ), .D ( signal_9197 ), .Q ( signal_9198 ) ) ;
    buf_clk cell_3640 ( .C ( clk ), .D ( signal_9231 ), .Q ( signal_9232 ) ) ;
    buf_clk cell_3644 ( .C ( clk ), .D ( signal_9235 ), .Q ( signal_9236 ) ) ;
    buf_clk cell_3648 ( .C ( clk ), .D ( signal_9239 ), .Q ( signal_9240 ) ) ;
    buf_clk cell_3652 ( .C ( clk ), .D ( signal_9243 ), .Q ( signal_9244 ) ) ;
    buf_clk cell_3656 ( .C ( clk ), .D ( signal_9247 ), .Q ( signal_9248 ) ) ;
    buf_clk cell_3660 ( .C ( clk ), .D ( signal_9251 ), .Q ( signal_9252 ) ) ;
    buf_clk cell_3664 ( .C ( clk ), .D ( signal_9255 ), .Q ( signal_9256 ) ) ;
    buf_clk cell_3668 ( .C ( clk ), .D ( signal_9259 ), .Q ( signal_9260 ) ) ;
    buf_clk cell_3672 ( .C ( clk ), .D ( signal_9263 ), .Q ( signal_9264 ) ) ;
    buf_clk cell_3682 ( .C ( clk ), .D ( signal_9273 ), .Q ( signal_9274 ) ) ;
    buf_clk cell_3686 ( .C ( clk ), .D ( signal_9277 ), .Q ( signal_9278 ) ) ;
    buf_clk cell_3690 ( .C ( clk ), .D ( signal_9281 ), .Q ( signal_9282 ) ) ;
    buf_clk cell_3724 ( .C ( clk ), .D ( signal_9315 ), .Q ( signal_9316 ) ) ;
    buf_clk cell_3728 ( .C ( clk ), .D ( signal_9319 ), .Q ( signal_9320 ) ) ;
    buf_clk cell_3732 ( .C ( clk ), .D ( signal_9323 ), .Q ( signal_9324 ) ) ;
    buf_clk cell_3736 ( .C ( clk ), .D ( signal_9327 ), .Q ( signal_9328 ) ) ;
    buf_clk cell_3740 ( .C ( clk ), .D ( signal_9331 ), .Q ( signal_9332 ) ) ;
    buf_clk cell_3744 ( .C ( clk ), .D ( signal_9335 ), .Q ( signal_9336 ) ) ;
    buf_clk cell_3754 ( .C ( clk ), .D ( signal_9345 ), .Q ( signal_9346 ) ) ;
    buf_clk cell_3758 ( .C ( clk ), .D ( signal_9349 ), .Q ( signal_9350 ) ) ;
    buf_clk cell_3762 ( .C ( clk ), .D ( signal_9353 ), .Q ( signal_9354 ) ) ;
    buf_clk cell_3778 ( .C ( clk ), .D ( signal_9369 ), .Q ( signal_9370 ) ) ;
    buf_clk cell_3782 ( .C ( clk ), .D ( signal_9373 ), .Q ( signal_9374 ) ) ;
    buf_clk cell_3786 ( .C ( clk ), .D ( signal_9377 ), .Q ( signal_9378 ) ) ;
    buf_clk cell_3790 ( .C ( clk ), .D ( signal_9381 ), .Q ( signal_9382 ) ) ;
    buf_clk cell_3794 ( .C ( clk ), .D ( signal_9385 ), .Q ( signal_9386 ) ) ;
    buf_clk cell_3798 ( .C ( clk ), .D ( signal_9389 ), .Q ( signal_9390 ) ) ;
    buf_clk cell_3802 ( .C ( clk ), .D ( signal_9393 ), .Q ( signal_9394 ) ) ;
    buf_clk cell_3806 ( .C ( clk ), .D ( signal_9397 ), .Q ( signal_9398 ) ) ;
    buf_clk cell_3810 ( .C ( clk ), .D ( signal_9401 ), .Q ( signal_9402 ) ) ;
    buf_clk cell_3820 ( .C ( clk ), .D ( signal_9411 ), .Q ( signal_9412 ) ) ;
    buf_clk cell_3824 ( .C ( clk ), .D ( signal_9415 ), .Q ( signal_9416 ) ) ;
    buf_clk cell_3828 ( .C ( clk ), .D ( signal_9419 ), .Q ( signal_9420 ) ) ;
    buf_clk cell_3832 ( .C ( clk ), .D ( signal_9423 ), .Q ( signal_9424 ) ) ;
    buf_clk cell_3836 ( .C ( clk ), .D ( signal_9427 ), .Q ( signal_9428 ) ) ;
    buf_clk cell_3840 ( .C ( clk ), .D ( signal_9431 ), .Q ( signal_9432 ) ) ;
    buf_clk cell_3850 ( .C ( clk ), .D ( signal_9441 ), .Q ( signal_9442 ) ) ;
    buf_clk cell_3854 ( .C ( clk ), .D ( signal_9445 ), .Q ( signal_9446 ) ) ;
    buf_clk cell_3858 ( .C ( clk ), .D ( signal_9449 ), .Q ( signal_9450 ) ) ;
    buf_clk cell_3880 ( .C ( clk ), .D ( signal_9471 ), .Q ( signal_9472 ) ) ;
    buf_clk cell_3884 ( .C ( clk ), .D ( signal_9475 ), .Q ( signal_9476 ) ) ;
    buf_clk cell_3888 ( .C ( clk ), .D ( signal_9479 ), .Q ( signal_9480 ) ) ;
    buf_clk cell_3898 ( .C ( clk ), .D ( signal_9489 ), .Q ( signal_9490 ) ) ;
    buf_clk cell_3904 ( .C ( clk ), .D ( signal_9495 ), .Q ( signal_9496 ) ) ;
    buf_clk cell_3910 ( .C ( clk ), .D ( signal_9501 ), .Q ( signal_9502 ) ) ;
    buf_clk cell_3916 ( .C ( clk ), .D ( signal_9507 ), .Q ( signal_9508 ) ) ;
    buf_clk cell_3922 ( .C ( clk ), .D ( signal_9513 ), .Q ( signal_9514 ) ) ;
    buf_clk cell_3928 ( .C ( clk ), .D ( signal_9519 ), .Q ( signal_9520 ) ) ;
    buf_clk cell_3934 ( .C ( clk ), .D ( signal_9525 ), .Q ( signal_9526 ) ) ;
    buf_clk cell_3940 ( .C ( clk ), .D ( signal_9531 ), .Q ( signal_9532 ) ) ;
    buf_clk cell_3946 ( .C ( clk ), .D ( signal_9537 ), .Q ( signal_9538 ) ) ;
    buf_clk cell_3964 ( .C ( clk ), .D ( signal_9555 ), .Q ( signal_9556 ) ) ;
    buf_clk cell_3970 ( .C ( clk ), .D ( signal_9561 ), .Q ( signal_9562 ) ) ;
    buf_clk cell_3976 ( .C ( clk ), .D ( signal_9567 ), .Q ( signal_9568 ) ) ;
    buf_clk cell_4042 ( .C ( clk ), .D ( signal_9633 ), .Q ( signal_9634 ) ) ;
    buf_clk cell_4048 ( .C ( clk ), .D ( signal_9639 ), .Q ( signal_9640 ) ) ;
    buf_clk cell_4054 ( .C ( clk ), .D ( signal_9645 ), .Q ( signal_9646 ) ) ;
    buf_clk cell_4132 ( .C ( clk ), .D ( signal_9723 ), .Q ( signal_9724 ) ) ;
    buf_clk cell_4138 ( .C ( clk ), .D ( signal_9729 ), .Q ( signal_9730 ) ) ;
    buf_clk cell_4144 ( .C ( clk ), .D ( signal_9735 ), .Q ( signal_9736 ) ) ;
    buf_clk cell_4180 ( .C ( clk ), .D ( signal_9771 ), .Q ( signal_9772 ) ) ;
    buf_clk cell_4186 ( .C ( clk ), .D ( signal_9777 ), .Q ( signal_9778 ) ) ;
    buf_clk cell_4192 ( .C ( clk ), .D ( signal_9783 ), .Q ( signal_9784 ) ) ;
    buf_clk cell_4264 ( .C ( clk ), .D ( signal_9855 ), .Q ( signal_9856 ) ) ;
    buf_clk cell_4270 ( .C ( clk ), .D ( signal_9861 ), .Q ( signal_9862 ) ) ;
    buf_clk cell_4276 ( .C ( clk ), .D ( signal_9867 ), .Q ( signal_9868 ) ) ;
    buf_clk cell_4294 ( .C ( clk ), .D ( signal_9885 ), .Q ( signal_9886 ) ) ;
    buf_clk cell_4300 ( .C ( clk ), .D ( signal_9891 ), .Q ( signal_9892 ) ) ;
    buf_clk cell_4306 ( .C ( clk ), .D ( signal_9897 ), .Q ( signal_9898 ) ) ;
    buf_clk cell_4378 ( .C ( clk ), .D ( signal_9969 ), .Q ( signal_9970 ) ) ;
    buf_clk cell_4384 ( .C ( clk ), .D ( signal_9975 ), .Q ( signal_9976 ) ) ;
    buf_clk cell_4390 ( .C ( clk ), .D ( signal_9981 ), .Q ( signal_9982 ) ) ;
    buf_clk cell_4420 ( .C ( clk ), .D ( signal_10011 ), .Q ( signal_10012 ) ) ;
    buf_clk cell_4426 ( .C ( clk ), .D ( signal_10017 ), .Q ( signal_10018 ) ) ;
    buf_clk cell_4432 ( .C ( clk ), .D ( signal_10023 ), .Q ( signal_10024 ) ) ;
    buf_clk cell_4438 ( .C ( clk ), .D ( signal_10029 ), .Q ( signal_10030 ) ) ;
    buf_clk cell_4444 ( .C ( clk ), .D ( signal_10035 ), .Q ( signal_10036 ) ) ;
    buf_clk cell_4450 ( .C ( clk ), .D ( signal_10041 ), .Q ( signal_10042 ) ) ;
    buf_clk cell_4456 ( .C ( clk ), .D ( signal_10047 ), .Q ( signal_10048 ) ) ;
    buf_clk cell_4462 ( .C ( clk ), .D ( signal_10053 ), .Q ( signal_10054 ) ) ;
    buf_clk cell_4468 ( .C ( clk ), .D ( signal_10059 ), .Q ( signal_10060 ) ) ;
    buf_clk cell_4498 ( .C ( clk ), .D ( signal_10089 ), .Q ( signal_10090 ) ) ;
    buf_clk cell_4506 ( .C ( clk ), .D ( signal_10097 ), .Q ( signal_10098 ) ) ;
    buf_clk cell_4514 ( .C ( clk ), .D ( signal_10105 ), .Q ( signal_10106 ) ) ;
    buf_clk cell_4756 ( .C ( clk ), .D ( signal_10347 ), .Q ( signal_10348 ) ) ;
    buf_clk cell_4764 ( .C ( clk ), .D ( signal_10355 ), .Q ( signal_10356 ) ) ;
    buf_clk cell_4772 ( .C ( clk ), .D ( signal_10363 ), .Q ( signal_10364 ) ) ;
    buf_clk cell_4852 ( .C ( clk ), .D ( signal_10443 ), .Q ( signal_10444 ) ) ;
    buf_clk cell_4860 ( .C ( clk ), .D ( signal_10451 ), .Q ( signal_10452 ) ) ;
    buf_clk cell_4868 ( .C ( clk ), .D ( signal_10459 ), .Q ( signal_10460 ) ) ;
    buf_clk cell_5002 ( .C ( clk ), .D ( signal_10593 ), .Q ( signal_10594 ) ) ;
    buf_clk cell_5012 ( .C ( clk ), .D ( signal_10603 ), .Q ( signal_10604 ) ) ;
    buf_clk cell_5022 ( .C ( clk ), .D ( signal_10613 ), .Q ( signal_10614 ) ) ;
    buf_clk cell_5146 ( .C ( clk ), .D ( signal_10737 ), .Q ( signal_10738 ) ) ;
    buf_clk cell_5156 ( .C ( clk ), .D ( signal_10747 ), .Q ( signal_10748 ) ) ;
    buf_clk cell_5166 ( .C ( clk ), .D ( signal_10757 ), .Q ( signal_10758 ) ) ;
    buf_clk cell_5314 ( .C ( clk ), .D ( signal_10905 ), .Q ( signal_10906 ) ) ;
    buf_clk cell_5324 ( .C ( clk ), .D ( signal_10915 ), .Q ( signal_10916 ) ) ;
    buf_clk cell_5334 ( .C ( clk ), .D ( signal_10925 ), .Q ( signal_10926 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_3333 ( .C ( clk ), .D ( signal_1550 ), .Q ( signal_8925 ) ) ;
    buf_clk cell_3335 ( .C ( clk ), .D ( signal_3624 ), .Q ( signal_8927 ) ) ;
    buf_clk cell_3337 ( .C ( clk ), .D ( signal_3625 ), .Q ( signal_8929 ) ) ;
    buf_clk cell_3339 ( .C ( clk ), .D ( signal_1566 ), .Q ( signal_8931 ) ) ;
    buf_clk cell_3341 ( .C ( clk ), .D ( signal_3656 ), .Q ( signal_8933 ) ) ;
    buf_clk cell_3343 ( .C ( clk ), .D ( signal_3657 ), .Q ( signal_8935 ) ) ;
    buf_clk cell_3347 ( .C ( clk ), .D ( signal_8938 ), .Q ( signal_8939 ) ) ;
    buf_clk cell_3351 ( .C ( clk ), .D ( signal_8942 ), .Q ( signal_8943 ) ) ;
    buf_clk cell_3355 ( .C ( clk ), .D ( signal_8946 ), .Q ( signal_8947 ) ) ;
    buf_clk cell_3357 ( .C ( clk ), .D ( signal_1604 ), .Q ( signal_8949 ) ) ;
    buf_clk cell_3359 ( .C ( clk ), .D ( signal_3732 ), .Q ( signal_8951 ) ) ;
    buf_clk cell_3361 ( .C ( clk ), .D ( signal_3733 ), .Q ( signal_8953 ) ) ;
    buf_clk cell_3365 ( .C ( clk ), .D ( signal_8956 ), .Q ( signal_8957 ) ) ;
    buf_clk cell_3369 ( .C ( clk ), .D ( signal_8960 ), .Q ( signal_8961 ) ) ;
    buf_clk cell_3373 ( .C ( clk ), .D ( signal_8964 ), .Q ( signal_8965 ) ) ;
    buf_clk cell_3377 ( .C ( clk ), .D ( signal_8968 ), .Q ( signal_8969 ) ) ;
    buf_clk cell_3381 ( .C ( clk ), .D ( signal_8972 ), .Q ( signal_8973 ) ) ;
    buf_clk cell_3385 ( .C ( clk ), .D ( signal_8976 ), .Q ( signal_8977 ) ) ;
    buf_clk cell_3389 ( .C ( clk ), .D ( signal_8980 ), .Q ( signal_8981 ) ) ;
    buf_clk cell_3393 ( .C ( clk ), .D ( signal_8984 ), .Q ( signal_8985 ) ) ;
    buf_clk cell_3397 ( .C ( clk ), .D ( signal_8988 ), .Q ( signal_8989 ) ) ;
    buf_clk cell_3405 ( .C ( clk ), .D ( signal_8996 ), .Q ( signal_8997 ) ) ;
    buf_clk cell_3413 ( .C ( clk ), .D ( signal_9004 ), .Q ( signal_9005 ) ) ;
    buf_clk cell_3421 ( .C ( clk ), .D ( signal_9012 ), .Q ( signal_9013 ) ) ;
    buf_clk cell_3423 ( .C ( clk ), .D ( signal_1576 ), .Q ( signal_9015 ) ) ;
    buf_clk cell_3425 ( .C ( clk ), .D ( signal_3676 ), .Q ( signal_9017 ) ) ;
    buf_clk cell_3427 ( .C ( clk ), .D ( signal_3677 ), .Q ( signal_9019 ) ) ;
    buf_clk cell_3429 ( .C ( clk ), .D ( signal_1582 ), .Q ( signal_9021 ) ) ;
    buf_clk cell_3431 ( .C ( clk ), .D ( signal_3688 ), .Q ( signal_9023 ) ) ;
    buf_clk cell_3433 ( .C ( clk ), .D ( signal_3689 ), .Q ( signal_9025 ) ) ;
    buf_clk cell_3437 ( .C ( clk ), .D ( signal_9028 ), .Q ( signal_9029 ) ) ;
    buf_clk cell_3441 ( .C ( clk ), .D ( signal_9032 ), .Q ( signal_9033 ) ) ;
    buf_clk cell_3445 ( .C ( clk ), .D ( signal_9036 ), .Q ( signal_9037 ) ) ;
    buf_clk cell_3447 ( .C ( clk ), .D ( signal_1632 ), .Q ( signal_9039 ) ) ;
    buf_clk cell_3449 ( .C ( clk ), .D ( signal_3788 ), .Q ( signal_9041 ) ) ;
    buf_clk cell_3451 ( .C ( clk ), .D ( signal_3789 ), .Q ( signal_9043 ) ) ;
    buf_clk cell_3453 ( .C ( clk ), .D ( signal_1597 ), .Q ( signal_9045 ) ) ;
    buf_clk cell_3455 ( .C ( clk ), .D ( signal_3718 ), .Q ( signal_9047 ) ) ;
    buf_clk cell_3457 ( .C ( clk ), .D ( signal_3719 ), .Q ( signal_9049 ) ) ;
    buf_clk cell_3461 ( .C ( clk ), .D ( signal_9052 ), .Q ( signal_9053 ) ) ;
    buf_clk cell_3465 ( .C ( clk ), .D ( signal_9056 ), .Q ( signal_9057 ) ) ;
    buf_clk cell_3469 ( .C ( clk ), .D ( signal_9060 ), .Q ( signal_9061 ) ) ;
    buf_clk cell_3471 ( .C ( clk ), .D ( signal_1595 ), .Q ( signal_9063 ) ) ;
    buf_clk cell_3473 ( .C ( clk ), .D ( signal_3714 ), .Q ( signal_9065 ) ) ;
    buf_clk cell_3475 ( .C ( clk ), .D ( signal_3715 ), .Q ( signal_9067 ) ) ;
    buf_clk cell_3477 ( .C ( clk ), .D ( signal_1551 ), .Q ( signal_9069 ) ) ;
    buf_clk cell_3479 ( .C ( clk ), .D ( signal_3626 ), .Q ( signal_9071 ) ) ;
    buf_clk cell_3481 ( .C ( clk ), .D ( signal_3627 ), .Q ( signal_9073 ) ) ;
    buf_clk cell_3483 ( .C ( clk ), .D ( signal_1613 ), .Q ( signal_9075 ) ) ;
    buf_clk cell_3485 ( .C ( clk ), .D ( signal_3750 ), .Q ( signal_9077 ) ) ;
    buf_clk cell_3487 ( .C ( clk ), .D ( signal_3751 ), .Q ( signal_9079 ) ) ;
    buf_clk cell_3489 ( .C ( clk ), .D ( signal_1690 ), .Q ( signal_9081 ) ) ;
    buf_clk cell_3491 ( .C ( clk ), .D ( signal_3904 ), .Q ( signal_9083 ) ) ;
    buf_clk cell_3493 ( .C ( clk ), .D ( signal_3905 ), .Q ( signal_9085 ) ) ;
    buf_clk cell_3495 ( .C ( clk ), .D ( signal_1555 ), .Q ( signal_9087 ) ) ;
    buf_clk cell_3497 ( .C ( clk ), .D ( signal_3634 ), .Q ( signal_9089 ) ) ;
    buf_clk cell_3499 ( .C ( clk ), .D ( signal_3635 ), .Q ( signal_9091 ) ) ;
    buf_clk cell_3503 ( .C ( clk ), .D ( signal_9094 ), .Q ( signal_9095 ) ) ;
    buf_clk cell_3507 ( .C ( clk ), .D ( signal_9098 ), .Q ( signal_9099 ) ) ;
    buf_clk cell_3511 ( .C ( clk ), .D ( signal_9102 ), .Q ( signal_9103 ) ) ;
    buf_clk cell_3513 ( .C ( clk ), .D ( signal_1562 ), .Q ( signal_9105 ) ) ;
    buf_clk cell_3515 ( .C ( clk ), .D ( signal_3648 ), .Q ( signal_9107 ) ) ;
    buf_clk cell_3517 ( .C ( clk ), .D ( signal_3649 ), .Q ( signal_9109 ) ) ;
    buf_clk cell_3519 ( .C ( clk ), .D ( signal_1694 ), .Q ( signal_9111 ) ) ;
    buf_clk cell_3521 ( .C ( clk ), .D ( signal_3912 ), .Q ( signal_9113 ) ) ;
    buf_clk cell_3523 ( .C ( clk ), .D ( signal_3913 ), .Q ( signal_9115 ) ) ;
    buf_clk cell_3525 ( .C ( clk ), .D ( signal_1636 ), .Q ( signal_9117 ) ) ;
    buf_clk cell_3527 ( .C ( clk ), .D ( signal_3796 ), .Q ( signal_9119 ) ) ;
    buf_clk cell_3529 ( .C ( clk ), .D ( signal_3797 ), .Q ( signal_9121 ) ) ;
    buf_clk cell_3531 ( .C ( clk ), .D ( signal_1568 ), .Q ( signal_9123 ) ) ;
    buf_clk cell_3533 ( .C ( clk ), .D ( signal_3660 ), .Q ( signal_9125 ) ) ;
    buf_clk cell_3535 ( .C ( clk ), .D ( signal_3661 ), .Q ( signal_9127 ) ) ;
    buf_clk cell_3539 ( .C ( clk ), .D ( signal_9130 ), .Q ( signal_9131 ) ) ;
    buf_clk cell_3543 ( .C ( clk ), .D ( signal_9134 ), .Q ( signal_9135 ) ) ;
    buf_clk cell_3547 ( .C ( clk ), .D ( signal_9138 ), .Q ( signal_9139 ) ) ;
    buf_clk cell_3549 ( .C ( clk ), .D ( signal_1853 ), .Q ( signal_9141 ) ) ;
    buf_clk cell_3551 ( .C ( clk ), .D ( signal_4230 ), .Q ( signal_9143 ) ) ;
    buf_clk cell_3553 ( .C ( clk ), .D ( signal_4231 ), .Q ( signal_9145 ) ) ;
    buf_clk cell_3555 ( .C ( clk ), .D ( signal_8860 ), .Q ( signal_9147 ) ) ;
    buf_clk cell_3557 ( .C ( clk ), .D ( signal_8862 ), .Q ( signal_9149 ) ) ;
    buf_clk cell_3559 ( .C ( clk ), .D ( signal_8864 ), .Q ( signal_9151 ) ) ;
    buf_clk cell_3563 ( .C ( clk ), .D ( signal_9154 ), .Q ( signal_9155 ) ) ;
    buf_clk cell_3567 ( .C ( clk ), .D ( signal_9158 ), .Q ( signal_9159 ) ) ;
    buf_clk cell_3571 ( .C ( clk ), .D ( signal_9162 ), .Q ( signal_9163 ) ) ;
    buf_clk cell_3575 ( .C ( clk ), .D ( signal_9166 ), .Q ( signal_9167 ) ) ;
    buf_clk cell_3579 ( .C ( clk ), .D ( signal_9170 ), .Q ( signal_9171 ) ) ;
    buf_clk cell_3583 ( .C ( clk ), .D ( signal_9174 ), .Q ( signal_9175 ) ) ;
    buf_clk cell_3587 ( .C ( clk ), .D ( signal_9178 ), .Q ( signal_9179 ) ) ;
    buf_clk cell_3591 ( .C ( clk ), .D ( signal_9182 ), .Q ( signal_9183 ) ) ;
    buf_clk cell_3595 ( .C ( clk ), .D ( signal_9186 ), .Q ( signal_9187 ) ) ;
    buf_clk cell_3599 ( .C ( clk ), .D ( signal_9190 ), .Q ( signal_9191 ) ) ;
    buf_clk cell_3603 ( .C ( clk ), .D ( signal_9194 ), .Q ( signal_9195 ) ) ;
    buf_clk cell_3607 ( .C ( clk ), .D ( signal_9198 ), .Q ( signal_9199 ) ) ;
    buf_clk cell_3609 ( .C ( clk ), .D ( signal_8788 ), .Q ( signal_9201 ) ) ;
    buf_clk cell_3611 ( .C ( clk ), .D ( signal_8790 ), .Q ( signal_9203 ) ) ;
    buf_clk cell_3613 ( .C ( clk ), .D ( signal_8792 ), .Q ( signal_9205 ) ) ;
    buf_clk cell_3615 ( .C ( clk ), .D ( signal_8662 ), .Q ( signal_9207 ) ) ;
    buf_clk cell_3617 ( .C ( clk ), .D ( signal_8664 ), .Q ( signal_9209 ) ) ;
    buf_clk cell_3619 ( .C ( clk ), .D ( signal_8666 ), .Q ( signal_9211 ) ) ;
    buf_clk cell_3621 ( .C ( clk ), .D ( signal_1854 ), .Q ( signal_9213 ) ) ;
    buf_clk cell_3623 ( .C ( clk ), .D ( signal_4232 ), .Q ( signal_9215 ) ) ;
    buf_clk cell_3625 ( .C ( clk ), .D ( signal_4233 ), .Q ( signal_9217 ) ) ;
    buf_clk cell_3627 ( .C ( clk ), .D ( signal_8452 ), .Q ( signal_9219 ) ) ;
    buf_clk cell_3629 ( .C ( clk ), .D ( signal_8454 ), .Q ( signal_9221 ) ) ;
    buf_clk cell_3631 ( .C ( clk ), .D ( signal_8456 ), .Q ( signal_9223 ) ) ;
    buf_clk cell_3633 ( .C ( clk ), .D ( signal_8896 ), .Q ( signal_9225 ) ) ;
    buf_clk cell_3635 ( .C ( clk ), .D ( signal_8898 ), .Q ( signal_9227 ) ) ;
    buf_clk cell_3637 ( .C ( clk ), .D ( signal_8900 ), .Q ( signal_9229 ) ) ;
    buf_clk cell_3641 ( .C ( clk ), .D ( signal_9232 ), .Q ( signal_9233 ) ) ;
    buf_clk cell_3645 ( .C ( clk ), .D ( signal_9236 ), .Q ( signal_9237 ) ) ;
    buf_clk cell_3649 ( .C ( clk ), .D ( signal_9240 ), .Q ( signal_9241 ) ) ;
    buf_clk cell_3653 ( .C ( clk ), .D ( signal_9244 ), .Q ( signal_9245 ) ) ;
    buf_clk cell_3657 ( .C ( clk ), .D ( signal_9248 ), .Q ( signal_9249 ) ) ;
    buf_clk cell_3661 ( .C ( clk ), .D ( signal_9252 ), .Q ( signal_9253 ) ) ;
    buf_clk cell_3665 ( .C ( clk ), .D ( signal_9256 ), .Q ( signal_9257 ) ) ;
    buf_clk cell_3669 ( .C ( clk ), .D ( signal_9260 ), .Q ( signal_9261 ) ) ;
    buf_clk cell_3673 ( .C ( clk ), .D ( signal_9264 ), .Q ( signal_9265 ) ) ;
    buf_clk cell_3675 ( .C ( clk ), .D ( signal_1862 ), .Q ( signal_9267 ) ) ;
    buf_clk cell_3677 ( .C ( clk ), .D ( signal_4248 ), .Q ( signal_9269 ) ) ;
    buf_clk cell_3679 ( .C ( clk ), .D ( signal_4249 ), .Q ( signal_9271 ) ) ;
    buf_clk cell_3683 ( .C ( clk ), .D ( signal_9274 ), .Q ( signal_9275 ) ) ;
    buf_clk cell_3687 ( .C ( clk ), .D ( signal_9278 ), .Q ( signal_9279 ) ) ;
    buf_clk cell_3691 ( .C ( clk ), .D ( signal_9282 ), .Q ( signal_9283 ) ) ;
    buf_clk cell_3693 ( .C ( clk ), .D ( signal_8500 ), .Q ( signal_9285 ) ) ;
    buf_clk cell_3695 ( .C ( clk ), .D ( signal_8502 ), .Q ( signal_9287 ) ) ;
    buf_clk cell_3697 ( .C ( clk ), .D ( signal_8504 ), .Q ( signal_9289 ) ) ;
    buf_clk cell_3699 ( .C ( clk ), .D ( signal_1866 ), .Q ( signal_9291 ) ) ;
    buf_clk cell_3701 ( .C ( clk ), .D ( signal_4256 ), .Q ( signal_9293 ) ) ;
    buf_clk cell_3703 ( .C ( clk ), .D ( signal_4257 ), .Q ( signal_9295 ) ) ;
    buf_clk cell_3705 ( .C ( clk ), .D ( signal_8422 ), .Q ( signal_9297 ) ) ;
    buf_clk cell_3707 ( .C ( clk ), .D ( signal_8424 ), .Q ( signal_9299 ) ) ;
    buf_clk cell_3709 ( .C ( clk ), .D ( signal_8426 ), .Q ( signal_9301 ) ) ;
    buf_clk cell_3711 ( .C ( clk ), .D ( signal_1873 ), .Q ( signal_9303 ) ) ;
    buf_clk cell_3713 ( .C ( clk ), .D ( signal_4270 ), .Q ( signal_9305 ) ) ;
    buf_clk cell_3715 ( .C ( clk ), .D ( signal_4271 ), .Q ( signal_9307 ) ) ;
    buf_clk cell_3717 ( .C ( clk ), .D ( signal_1851 ), .Q ( signal_9309 ) ) ;
    buf_clk cell_3719 ( .C ( clk ), .D ( signal_4226 ), .Q ( signal_9311 ) ) ;
    buf_clk cell_3721 ( .C ( clk ), .D ( signal_4227 ), .Q ( signal_9313 ) ) ;
    buf_clk cell_3725 ( .C ( clk ), .D ( signal_9316 ), .Q ( signal_9317 ) ) ;
    buf_clk cell_3729 ( .C ( clk ), .D ( signal_9320 ), .Q ( signal_9321 ) ) ;
    buf_clk cell_3733 ( .C ( clk ), .D ( signal_9324 ), .Q ( signal_9325 ) ) ;
    buf_clk cell_3737 ( .C ( clk ), .D ( signal_9328 ), .Q ( signal_9329 ) ) ;
    buf_clk cell_3741 ( .C ( clk ), .D ( signal_9332 ), .Q ( signal_9333 ) ) ;
    buf_clk cell_3745 ( .C ( clk ), .D ( signal_9336 ), .Q ( signal_9337 ) ) ;
    buf_clk cell_3747 ( .C ( clk ), .D ( signal_1571 ), .Q ( signal_9339 ) ) ;
    buf_clk cell_3749 ( .C ( clk ), .D ( signal_3666 ), .Q ( signal_9341 ) ) ;
    buf_clk cell_3751 ( .C ( clk ), .D ( signal_3667 ), .Q ( signal_9343 ) ) ;
    buf_clk cell_3755 ( .C ( clk ), .D ( signal_9346 ), .Q ( signal_9347 ) ) ;
    buf_clk cell_3759 ( .C ( clk ), .D ( signal_9350 ), .Q ( signal_9351 ) ) ;
    buf_clk cell_3763 ( .C ( clk ), .D ( signal_9354 ), .Q ( signal_9355 ) ) ;
    buf_clk cell_3765 ( .C ( clk ), .D ( signal_1540 ), .Q ( signal_9357 ) ) ;
    buf_clk cell_3767 ( .C ( clk ), .D ( signal_3604 ), .Q ( signal_9359 ) ) ;
    buf_clk cell_3769 ( .C ( clk ), .D ( signal_3605 ), .Q ( signal_9361 ) ) ;
    buf_clk cell_3771 ( .C ( clk ), .D ( signal_1872 ), .Q ( signal_9363 ) ) ;
    buf_clk cell_3773 ( .C ( clk ), .D ( signal_4268 ), .Q ( signal_9365 ) ) ;
    buf_clk cell_3775 ( .C ( clk ), .D ( signal_4269 ), .Q ( signal_9367 ) ) ;
    buf_clk cell_3779 ( .C ( clk ), .D ( signal_9370 ), .Q ( signal_9371 ) ) ;
    buf_clk cell_3783 ( .C ( clk ), .D ( signal_9374 ), .Q ( signal_9375 ) ) ;
    buf_clk cell_3787 ( .C ( clk ), .D ( signal_9378 ), .Q ( signal_9379 ) ) ;
    buf_clk cell_3791 ( .C ( clk ), .D ( signal_9382 ), .Q ( signal_9383 ) ) ;
    buf_clk cell_3795 ( .C ( clk ), .D ( signal_9386 ), .Q ( signal_9387 ) ) ;
    buf_clk cell_3799 ( .C ( clk ), .D ( signal_9390 ), .Q ( signal_9391 ) ) ;
    buf_clk cell_3803 ( .C ( clk ), .D ( signal_9394 ), .Q ( signal_9395 ) ) ;
    buf_clk cell_3807 ( .C ( clk ), .D ( signal_9398 ), .Q ( signal_9399 ) ) ;
    buf_clk cell_3811 ( .C ( clk ), .D ( signal_9402 ), .Q ( signal_9403 ) ) ;
    buf_clk cell_3813 ( .C ( clk ), .D ( signal_1583 ), .Q ( signal_9405 ) ) ;
    buf_clk cell_3815 ( .C ( clk ), .D ( signal_3690 ), .Q ( signal_9407 ) ) ;
    buf_clk cell_3817 ( .C ( clk ), .D ( signal_3691 ), .Q ( signal_9409 ) ) ;
    buf_clk cell_3821 ( .C ( clk ), .D ( signal_9412 ), .Q ( signal_9413 ) ) ;
    buf_clk cell_3825 ( .C ( clk ), .D ( signal_9416 ), .Q ( signal_9417 ) ) ;
    buf_clk cell_3829 ( .C ( clk ), .D ( signal_9420 ), .Q ( signal_9421 ) ) ;
    buf_clk cell_3833 ( .C ( clk ), .D ( signal_9424 ), .Q ( signal_9425 ) ) ;
    buf_clk cell_3837 ( .C ( clk ), .D ( signal_9428 ), .Q ( signal_9429 ) ) ;
    buf_clk cell_3841 ( .C ( clk ), .D ( signal_9432 ), .Q ( signal_9433 ) ) ;
    buf_clk cell_3843 ( .C ( clk ), .D ( signal_1600 ), .Q ( signal_9435 ) ) ;
    buf_clk cell_3845 ( .C ( clk ), .D ( signal_3724 ), .Q ( signal_9437 ) ) ;
    buf_clk cell_3847 ( .C ( clk ), .D ( signal_3725 ), .Q ( signal_9439 ) ) ;
    buf_clk cell_3851 ( .C ( clk ), .D ( signal_9442 ), .Q ( signal_9443 ) ) ;
    buf_clk cell_3855 ( .C ( clk ), .D ( signal_9446 ), .Q ( signal_9447 ) ) ;
    buf_clk cell_3859 ( .C ( clk ), .D ( signal_9450 ), .Q ( signal_9451 ) ) ;
    buf_clk cell_3861 ( .C ( clk ), .D ( signal_1870 ), .Q ( signal_9453 ) ) ;
    buf_clk cell_3863 ( .C ( clk ), .D ( signal_4264 ), .Q ( signal_9455 ) ) ;
    buf_clk cell_3865 ( .C ( clk ), .D ( signal_4265 ), .Q ( signal_9457 ) ) ;
    buf_clk cell_3867 ( .C ( clk ), .D ( signal_1312 ), .Q ( signal_9459 ) ) ;
    buf_clk cell_3869 ( .C ( clk ), .D ( signal_3148 ), .Q ( signal_9461 ) ) ;
    buf_clk cell_3871 ( .C ( clk ), .D ( signal_3149 ), .Q ( signal_9463 ) ) ;
    buf_clk cell_3873 ( .C ( clk ), .D ( signal_8476 ), .Q ( signal_9465 ) ) ;
    buf_clk cell_3875 ( .C ( clk ), .D ( signal_8478 ), .Q ( signal_9467 ) ) ;
    buf_clk cell_3877 ( .C ( clk ), .D ( signal_8480 ), .Q ( signal_9469 ) ) ;
    buf_clk cell_3881 ( .C ( clk ), .D ( signal_9472 ), .Q ( signal_9473 ) ) ;
    buf_clk cell_3885 ( .C ( clk ), .D ( signal_9476 ), .Q ( signal_9477 ) ) ;
    buf_clk cell_3889 ( .C ( clk ), .D ( signal_9480 ), .Q ( signal_9481 ) ) ;
    buf_clk cell_3899 ( .C ( clk ), .D ( signal_9490 ), .Q ( signal_9491 ) ) ;
    buf_clk cell_3905 ( .C ( clk ), .D ( signal_9496 ), .Q ( signal_9497 ) ) ;
    buf_clk cell_3911 ( .C ( clk ), .D ( signal_9502 ), .Q ( signal_9503 ) ) ;
    buf_clk cell_3917 ( .C ( clk ), .D ( signal_9508 ), .Q ( signal_9509 ) ) ;
    buf_clk cell_3923 ( .C ( clk ), .D ( signal_9514 ), .Q ( signal_9515 ) ) ;
    buf_clk cell_3929 ( .C ( clk ), .D ( signal_9520 ), .Q ( signal_9521 ) ) ;
    buf_clk cell_3935 ( .C ( clk ), .D ( signal_9526 ), .Q ( signal_9527 ) ) ;
    buf_clk cell_3941 ( .C ( clk ), .D ( signal_9532 ), .Q ( signal_9533 ) ) ;
    buf_clk cell_3947 ( .C ( clk ), .D ( signal_9538 ), .Q ( signal_9539 ) ) ;
    buf_clk cell_3951 ( .C ( clk ), .D ( signal_1537 ), .Q ( signal_9543 ) ) ;
    buf_clk cell_3955 ( .C ( clk ), .D ( signal_3598 ), .Q ( signal_9547 ) ) ;
    buf_clk cell_3959 ( .C ( clk ), .D ( signal_3599 ), .Q ( signal_9551 ) ) ;
    buf_clk cell_3965 ( .C ( clk ), .D ( signal_9556 ), .Q ( signal_9557 ) ) ;
    buf_clk cell_3971 ( .C ( clk ), .D ( signal_9562 ), .Q ( signal_9563 ) ) ;
    buf_clk cell_3977 ( .C ( clk ), .D ( signal_9568 ), .Q ( signal_9569 ) ) ;
    buf_clk cell_3981 ( .C ( clk ), .D ( signal_1552 ), .Q ( signal_9573 ) ) ;
    buf_clk cell_3985 ( .C ( clk ), .D ( signal_3628 ), .Q ( signal_9577 ) ) ;
    buf_clk cell_3989 ( .C ( clk ), .D ( signal_3629 ), .Q ( signal_9581 ) ) ;
    buf_clk cell_3993 ( .C ( clk ), .D ( signal_1618 ), .Q ( signal_9585 ) ) ;
    buf_clk cell_3997 ( .C ( clk ), .D ( signal_3760 ), .Q ( signal_9589 ) ) ;
    buf_clk cell_4001 ( .C ( clk ), .D ( signal_3761 ), .Q ( signal_9593 ) ) ;
    buf_clk cell_4005 ( .C ( clk ), .D ( signal_1560 ), .Q ( signal_9597 ) ) ;
    buf_clk cell_4009 ( .C ( clk ), .D ( signal_3644 ), .Q ( signal_9601 ) ) ;
    buf_clk cell_4013 ( .C ( clk ), .D ( signal_3645 ), .Q ( signal_9605 ) ) ;
    buf_clk cell_4017 ( .C ( clk ), .D ( signal_1622 ), .Q ( signal_9609 ) ) ;
    buf_clk cell_4021 ( .C ( clk ), .D ( signal_3768 ), .Q ( signal_9613 ) ) ;
    buf_clk cell_4025 ( .C ( clk ), .D ( signal_3769 ), .Q ( signal_9617 ) ) ;
    buf_clk cell_4029 ( .C ( clk ), .D ( signal_1533 ), .Q ( signal_9621 ) ) ;
    buf_clk cell_4033 ( .C ( clk ), .D ( signal_3590 ), .Q ( signal_9625 ) ) ;
    buf_clk cell_4037 ( .C ( clk ), .D ( signal_3591 ), .Q ( signal_9629 ) ) ;
    buf_clk cell_4043 ( .C ( clk ), .D ( signal_9634 ), .Q ( signal_9635 ) ) ;
    buf_clk cell_4049 ( .C ( clk ), .D ( signal_9640 ), .Q ( signal_9641 ) ) ;
    buf_clk cell_4055 ( .C ( clk ), .D ( signal_9646 ), .Q ( signal_9647 ) ) ;
    buf_clk cell_4059 ( .C ( clk ), .D ( signal_8518 ), .Q ( signal_9651 ) ) ;
    buf_clk cell_4063 ( .C ( clk ), .D ( signal_8520 ), .Q ( signal_9655 ) ) ;
    buf_clk cell_4067 ( .C ( clk ), .D ( signal_8522 ), .Q ( signal_9659 ) ) ;
    buf_clk cell_4101 ( .C ( clk ), .D ( signal_1591 ), .Q ( signal_9693 ) ) ;
    buf_clk cell_4105 ( .C ( clk ), .D ( signal_3706 ), .Q ( signal_9697 ) ) ;
    buf_clk cell_4109 ( .C ( clk ), .D ( signal_3707 ), .Q ( signal_9701 ) ) ;
    buf_clk cell_4133 ( .C ( clk ), .D ( signal_9724 ), .Q ( signal_9725 ) ) ;
    buf_clk cell_4139 ( .C ( clk ), .D ( signal_9730 ), .Q ( signal_9731 ) ) ;
    buf_clk cell_4145 ( .C ( clk ), .D ( signal_9736 ), .Q ( signal_9737 ) ) ;
    buf_clk cell_4155 ( .C ( clk ), .D ( signal_1621 ), .Q ( signal_9747 ) ) ;
    buf_clk cell_4159 ( .C ( clk ), .D ( signal_3766 ), .Q ( signal_9751 ) ) ;
    buf_clk cell_4163 ( .C ( clk ), .D ( signal_3767 ), .Q ( signal_9755 ) ) ;
    buf_clk cell_4181 ( .C ( clk ), .D ( signal_9772 ), .Q ( signal_9773 ) ) ;
    buf_clk cell_4187 ( .C ( clk ), .D ( signal_9778 ), .Q ( signal_9779 ) ) ;
    buf_clk cell_4193 ( .C ( clk ), .D ( signal_9784 ), .Q ( signal_9785 ) ) ;
    buf_clk cell_4197 ( .C ( clk ), .D ( signal_8902 ), .Q ( signal_9789 ) ) ;
    buf_clk cell_4201 ( .C ( clk ), .D ( signal_8904 ), .Q ( signal_9793 ) ) ;
    buf_clk cell_4205 ( .C ( clk ), .D ( signal_8906 ), .Q ( signal_9797 ) ) ;
    buf_clk cell_4221 ( .C ( clk ), .D ( signal_1606 ), .Q ( signal_9813 ) ) ;
    buf_clk cell_4225 ( .C ( clk ), .D ( signal_3736 ), .Q ( signal_9817 ) ) ;
    buf_clk cell_4229 ( .C ( clk ), .D ( signal_3737 ), .Q ( signal_9821 ) ) ;
    buf_clk cell_4233 ( .C ( clk ), .D ( signal_1691 ), .Q ( signal_9825 ) ) ;
    buf_clk cell_4237 ( .C ( clk ), .D ( signal_3906 ), .Q ( signal_9829 ) ) ;
    buf_clk cell_4241 ( .C ( clk ), .D ( signal_3907 ), .Q ( signal_9833 ) ) ;
    buf_clk cell_4245 ( .C ( clk ), .D ( signal_1570 ), .Q ( signal_9837 ) ) ;
    buf_clk cell_4249 ( .C ( clk ), .D ( signal_3664 ), .Q ( signal_9841 ) ) ;
    buf_clk cell_4253 ( .C ( clk ), .D ( signal_3665 ), .Q ( signal_9845 ) ) ;
    buf_clk cell_4265 ( .C ( clk ), .D ( signal_9856 ), .Q ( signal_9857 ) ) ;
    buf_clk cell_4271 ( .C ( clk ), .D ( signal_9862 ), .Q ( signal_9863 ) ) ;
    buf_clk cell_4277 ( .C ( clk ), .D ( signal_9868 ), .Q ( signal_9869 ) ) ;
    buf_clk cell_4281 ( .C ( clk ), .D ( signal_1584 ), .Q ( signal_9873 ) ) ;
    buf_clk cell_4285 ( .C ( clk ), .D ( signal_3692 ), .Q ( signal_9877 ) ) ;
    buf_clk cell_4289 ( .C ( clk ), .D ( signal_3693 ), .Q ( signal_9881 ) ) ;
    buf_clk cell_4295 ( .C ( clk ), .D ( signal_9886 ), .Q ( signal_9887 ) ) ;
    buf_clk cell_4301 ( .C ( clk ), .D ( signal_9892 ), .Q ( signal_9893 ) ) ;
    buf_clk cell_4307 ( .C ( clk ), .D ( signal_9898 ), .Q ( signal_9899 ) ) ;
    buf_clk cell_4311 ( .C ( clk ), .D ( signal_1590 ), .Q ( signal_9903 ) ) ;
    buf_clk cell_4315 ( .C ( clk ), .D ( signal_3704 ), .Q ( signal_9907 ) ) ;
    buf_clk cell_4319 ( .C ( clk ), .D ( signal_3705 ), .Q ( signal_9911 ) ) ;
    buf_clk cell_4323 ( .C ( clk ), .D ( signal_1675 ), .Q ( signal_9915 ) ) ;
    buf_clk cell_4327 ( .C ( clk ), .D ( signal_3874 ), .Q ( signal_9919 ) ) ;
    buf_clk cell_4331 ( .C ( clk ), .D ( signal_3875 ), .Q ( signal_9923 ) ) ;
    buf_clk cell_4335 ( .C ( clk ), .D ( signal_1598 ), .Q ( signal_9927 ) ) ;
    buf_clk cell_4339 ( .C ( clk ), .D ( signal_3720 ), .Q ( signal_9931 ) ) ;
    buf_clk cell_4343 ( .C ( clk ), .D ( signal_3721 ), .Q ( signal_9935 ) ) ;
    buf_clk cell_4353 ( .C ( clk ), .D ( signal_1601 ), .Q ( signal_9945 ) ) ;
    buf_clk cell_4357 ( .C ( clk ), .D ( signal_3726 ), .Q ( signal_9949 ) ) ;
    buf_clk cell_4361 ( .C ( clk ), .D ( signal_3727 ), .Q ( signal_9953 ) ) ;
    buf_clk cell_4365 ( .C ( clk ), .D ( signal_1543 ), .Q ( signal_9957 ) ) ;
    buf_clk cell_4369 ( .C ( clk ), .D ( signal_3610 ), .Q ( signal_9961 ) ) ;
    buf_clk cell_4373 ( .C ( clk ), .D ( signal_3611 ), .Q ( signal_9965 ) ) ;
    buf_clk cell_4379 ( .C ( clk ), .D ( signal_9970 ), .Q ( signal_9971 ) ) ;
    buf_clk cell_4385 ( .C ( clk ), .D ( signal_9976 ), .Q ( signal_9977 ) ) ;
    buf_clk cell_4391 ( .C ( clk ), .D ( signal_9982 ), .Q ( signal_9983 ) ) ;
    buf_clk cell_4407 ( .C ( clk ), .D ( signal_1625 ), .Q ( signal_9999 ) ) ;
    buf_clk cell_4411 ( .C ( clk ), .D ( signal_3774 ), .Q ( signal_10003 ) ) ;
    buf_clk cell_4415 ( .C ( clk ), .D ( signal_3775 ), .Q ( signal_10007 ) ) ;
    buf_clk cell_4421 ( .C ( clk ), .D ( signal_10012 ), .Q ( signal_10013 ) ) ;
    buf_clk cell_4427 ( .C ( clk ), .D ( signal_10018 ), .Q ( signal_10019 ) ) ;
    buf_clk cell_4433 ( .C ( clk ), .D ( signal_10024 ), .Q ( signal_10025 ) ) ;
    buf_clk cell_4439 ( .C ( clk ), .D ( signal_10030 ), .Q ( signal_10031 ) ) ;
    buf_clk cell_4445 ( .C ( clk ), .D ( signal_10036 ), .Q ( signal_10037 ) ) ;
    buf_clk cell_4451 ( .C ( clk ), .D ( signal_10042 ), .Q ( signal_10043 ) ) ;
    buf_clk cell_4457 ( .C ( clk ), .D ( signal_10048 ), .Q ( signal_10049 ) ) ;
    buf_clk cell_4463 ( .C ( clk ), .D ( signal_10054 ), .Q ( signal_10055 ) ) ;
    buf_clk cell_4469 ( .C ( clk ), .D ( signal_10060 ), .Q ( signal_10061 ) ) ;
    buf_clk cell_4473 ( .C ( clk ), .D ( signal_8774 ), .Q ( signal_10065 ) ) ;
    buf_clk cell_4477 ( .C ( clk ), .D ( signal_8780 ), .Q ( signal_10069 ) ) ;
    buf_clk cell_4481 ( .C ( clk ), .D ( signal_8786 ), .Q ( signal_10073 ) ) ;
    buf_clk cell_4499 ( .C ( clk ), .D ( signal_10090 ), .Q ( signal_10091 ) ) ;
    buf_clk cell_4507 ( .C ( clk ), .D ( signal_10098 ), .Q ( signal_10099 ) ) ;
    buf_clk cell_4515 ( .C ( clk ), .D ( signal_10106 ), .Q ( signal_10107 ) ) ;
    buf_clk cell_4533 ( .C ( clk ), .D ( signal_1645 ), .Q ( signal_10125 ) ) ;
    buf_clk cell_4539 ( .C ( clk ), .D ( signal_3814 ), .Q ( signal_10131 ) ) ;
    buf_clk cell_4545 ( .C ( clk ), .D ( signal_3815 ), .Q ( signal_10137 ) ) ;
    buf_clk cell_4551 ( .C ( clk ), .D ( signal_1616 ), .Q ( signal_10143 ) ) ;
    buf_clk cell_4557 ( .C ( clk ), .D ( signal_3756 ), .Q ( signal_10149 ) ) ;
    buf_clk cell_4563 ( .C ( clk ), .D ( signal_3757 ), .Q ( signal_10155 ) ) ;
    buf_clk cell_4581 ( .C ( clk ), .D ( signal_1534 ), .Q ( signal_10173 ) ) ;
    buf_clk cell_4587 ( .C ( clk ), .D ( signal_3592 ), .Q ( signal_10179 ) ) ;
    buf_clk cell_4593 ( .C ( clk ), .D ( signal_3593 ), .Q ( signal_10185 ) ) ;
    buf_clk cell_4635 ( .C ( clk ), .D ( signal_1850 ), .Q ( signal_10227 ) ) ;
    buf_clk cell_4641 ( .C ( clk ), .D ( signal_4224 ), .Q ( signal_10233 ) ) ;
    buf_clk cell_4647 ( .C ( clk ), .D ( signal_4225 ), .Q ( signal_10239 ) ) ;
    buf_clk cell_4653 ( .C ( clk ), .D ( signal_1631 ), .Q ( signal_10245 ) ) ;
    buf_clk cell_4659 ( .C ( clk ), .D ( signal_3786 ), .Q ( signal_10251 ) ) ;
    buf_clk cell_4665 ( .C ( clk ), .D ( signal_3787 ), .Q ( signal_10257 ) ) ;
    buf_clk cell_4671 ( .C ( clk ), .D ( signal_1683 ), .Q ( signal_10263 ) ) ;
    buf_clk cell_4677 ( .C ( clk ), .D ( signal_3890 ), .Q ( signal_10269 ) ) ;
    buf_clk cell_4683 ( .C ( clk ), .D ( signal_3891 ), .Q ( signal_10275 ) ) ;
    buf_clk cell_4707 ( .C ( clk ), .D ( signal_1299 ), .Q ( signal_10299 ) ) ;
    buf_clk cell_4713 ( .C ( clk ), .D ( signal_3122 ), .Q ( signal_10305 ) ) ;
    buf_clk cell_4719 ( .C ( clk ), .D ( signal_3123 ), .Q ( signal_10311 ) ) ;
    buf_clk cell_4731 ( .C ( clk ), .D ( signal_1557 ), .Q ( signal_10323 ) ) ;
    buf_clk cell_4737 ( .C ( clk ), .D ( signal_3638 ), .Q ( signal_10329 ) ) ;
    buf_clk cell_4743 ( .C ( clk ), .D ( signal_3639 ), .Q ( signal_10335 ) ) ;
    buf_clk cell_4757 ( .C ( clk ), .D ( signal_10348 ), .Q ( signal_10349 ) ) ;
    buf_clk cell_4765 ( .C ( clk ), .D ( signal_10356 ), .Q ( signal_10357 ) ) ;
    buf_clk cell_4773 ( .C ( clk ), .D ( signal_10364 ), .Q ( signal_10365 ) ) ;
    buf_clk cell_4803 ( .C ( clk ), .D ( signal_1506 ), .Q ( signal_10395 ) ) ;
    buf_clk cell_4809 ( .C ( clk ), .D ( signal_3536 ), .Q ( signal_10401 ) ) ;
    buf_clk cell_4815 ( .C ( clk ), .D ( signal_3537 ), .Q ( signal_10407 ) ) ;
    buf_clk cell_4821 ( .C ( clk ), .D ( signal_1593 ), .Q ( signal_10413 ) ) ;
    buf_clk cell_4827 ( .C ( clk ), .D ( signal_3710 ), .Q ( signal_10419 ) ) ;
    buf_clk cell_4833 ( .C ( clk ), .D ( signal_3711 ), .Q ( signal_10425 ) ) ;
    buf_clk cell_4853 ( .C ( clk ), .D ( signal_10444 ), .Q ( signal_10445 ) ) ;
    buf_clk cell_4861 ( .C ( clk ), .D ( signal_10452 ), .Q ( signal_10453 ) ) ;
    buf_clk cell_4869 ( .C ( clk ), .D ( signal_10460 ), .Q ( signal_10461 ) ) ;
    buf_clk cell_4875 ( .C ( clk ), .D ( signal_1338 ), .Q ( signal_10467 ) ) ;
    buf_clk cell_4881 ( .C ( clk ), .D ( signal_3200 ), .Q ( signal_10473 ) ) ;
    buf_clk cell_4887 ( .C ( clk ), .D ( signal_3201 ), .Q ( signal_10479 ) ) ;
    buf_clk cell_4893 ( .C ( clk ), .D ( signal_8464 ), .Q ( signal_10485 ) ) ;
    buf_clk cell_4899 ( .C ( clk ), .D ( signal_8466 ), .Q ( signal_10491 ) ) ;
    buf_clk cell_4905 ( .C ( clk ), .D ( signal_8468 ), .Q ( signal_10497 ) ) ;
    buf_clk cell_4923 ( .C ( clk ), .D ( signal_8734 ), .Q ( signal_10515 ) ) ;
    buf_clk cell_4929 ( .C ( clk ), .D ( signal_8736 ), .Q ( signal_10521 ) ) ;
    buf_clk cell_4935 ( .C ( clk ), .D ( signal_8738 ), .Q ( signal_10527 ) ) ;
    buf_clk cell_4953 ( .C ( clk ), .D ( signal_1637 ), .Q ( signal_10545 ) ) ;
    buf_clk cell_4959 ( .C ( clk ), .D ( signal_3798 ), .Q ( signal_10551 ) ) ;
    buf_clk cell_4965 ( .C ( clk ), .D ( signal_3799 ), .Q ( signal_10557 ) ) ;
    buf_clk cell_4971 ( .C ( clk ), .D ( signal_1518 ), .Q ( signal_10563 ) ) ;
    buf_clk cell_4977 ( .C ( clk ), .D ( signal_3560 ), .Q ( signal_10569 ) ) ;
    buf_clk cell_4983 ( .C ( clk ), .D ( signal_3561 ), .Q ( signal_10575 ) ) ;
    buf_clk cell_5003 ( .C ( clk ), .D ( signal_10594 ), .Q ( signal_10595 ) ) ;
    buf_clk cell_5013 ( .C ( clk ), .D ( signal_10604 ), .Q ( signal_10605 ) ) ;
    buf_clk cell_5023 ( .C ( clk ), .D ( signal_10614 ), .Q ( signal_10615 ) ) ;
    buf_clk cell_5049 ( .C ( clk ), .D ( signal_1619 ), .Q ( signal_10641 ) ) ;
    buf_clk cell_5057 ( .C ( clk ), .D ( signal_3762 ), .Q ( signal_10649 ) ) ;
    buf_clk cell_5065 ( .C ( clk ), .D ( signal_3763 ), .Q ( signal_10657 ) ) ;
    buf_clk cell_5073 ( .C ( clk ), .D ( signal_1350 ), .Q ( signal_10665 ) ) ;
    buf_clk cell_5081 ( .C ( clk ), .D ( signal_3224 ), .Q ( signal_10673 ) ) ;
    buf_clk cell_5089 ( .C ( clk ), .D ( signal_3225 ), .Q ( signal_10681 ) ) ;
    buf_clk cell_5147 ( .C ( clk ), .D ( signal_10738 ), .Q ( signal_10739 ) ) ;
    buf_clk cell_5157 ( .C ( clk ), .D ( signal_10748 ), .Q ( signal_10749 ) ) ;
    buf_clk cell_5167 ( .C ( clk ), .D ( signal_10758 ), .Q ( signal_10759 ) ) ;
    buf_clk cell_5199 ( .C ( clk ), .D ( signal_1575 ), .Q ( signal_10791 ) ) ;
    buf_clk cell_5207 ( .C ( clk ), .D ( signal_3674 ), .Q ( signal_10799 ) ) ;
    buf_clk cell_5215 ( .C ( clk ), .D ( signal_3675 ), .Q ( signal_10807 ) ) ;
    buf_clk cell_5241 ( .C ( clk ), .D ( signal_1587 ), .Q ( signal_10833 ) ) ;
    buf_clk cell_5249 ( .C ( clk ), .D ( signal_3698 ), .Q ( signal_10841 ) ) ;
    buf_clk cell_5257 ( .C ( clk ), .D ( signal_3699 ), .Q ( signal_10849 ) ) ;
    buf_clk cell_5265 ( .C ( clk ), .D ( signal_1861 ), .Q ( signal_10857 ) ) ;
    buf_clk cell_5273 ( .C ( clk ), .D ( signal_4246 ), .Q ( signal_10865 ) ) ;
    buf_clk cell_5281 ( .C ( clk ), .D ( signal_4247 ), .Q ( signal_10873 ) ) ;
    buf_clk cell_5289 ( .C ( clk ), .D ( signal_1258 ), .Q ( signal_10881 ) ) ;
    buf_clk cell_5297 ( .C ( clk ), .D ( signal_3040 ), .Q ( signal_10889 ) ) ;
    buf_clk cell_5305 ( .C ( clk ), .D ( signal_3041 ), .Q ( signal_10897 ) ) ;
    buf_clk cell_5315 ( .C ( clk ), .D ( signal_10906 ), .Q ( signal_10907 ) ) ;
    buf_clk cell_5325 ( .C ( clk ), .D ( signal_10916 ), .Q ( signal_10917 ) ) ;
    buf_clk cell_5335 ( .C ( clk ), .D ( signal_10926 ), .Q ( signal_10927 ) ) ;
    buf_clk cell_5343 ( .C ( clk ), .D ( signal_8512 ), .Q ( signal_10935 ) ) ;
    buf_clk cell_5351 ( .C ( clk ), .D ( signal_8514 ), .Q ( signal_10943 ) ) ;
    buf_clk cell_5359 ( .C ( clk ), .D ( signal_8516 ), .Q ( signal_10951 ) ) ;
    buf_clk cell_5367 ( .C ( clk ), .D ( signal_1614 ), .Q ( signal_10959 ) ) ;
    buf_clk cell_5375 ( .C ( clk ), .D ( signal_3752 ), .Q ( signal_10967 ) ) ;
    buf_clk cell_5383 ( .C ( clk ), .D ( signal_3753 ), .Q ( signal_10975 ) ) ;
    buf_clk cell_5397 ( .C ( clk ), .D ( signal_1549 ), .Q ( signal_10989 ) ) ;
    buf_clk cell_5405 ( .C ( clk ), .D ( signal_3622 ), .Q ( signal_10997 ) ) ;
    buf_clk cell_5413 ( .C ( clk ), .D ( signal_3623 ), .Q ( signal_11005 ) ) ;
    buf_clk cell_5421 ( .C ( clk ), .D ( signal_1578 ), .Q ( signal_11013 ) ) ;
    buf_clk cell_5429 ( .C ( clk ), .D ( signal_3680 ), .Q ( signal_11021 ) ) ;
    buf_clk cell_5437 ( .C ( clk ), .D ( signal_3681 ), .Q ( signal_11029 ) ) ;
    buf_clk cell_5445 ( .C ( clk ), .D ( signal_1581 ), .Q ( signal_11037 ) ) ;
    buf_clk cell_5453 ( .C ( clk ), .D ( signal_3686 ), .Q ( signal_11045 ) ) ;
    buf_clk cell_5461 ( .C ( clk ), .D ( signal_3687 ), .Q ( signal_11053 ) ) ;
    buf_clk cell_5571 ( .C ( clk ), .D ( signal_1505 ), .Q ( signal_11163 ) ) ;
    buf_clk cell_5581 ( .C ( clk ), .D ( signal_3534 ), .Q ( signal_11173 ) ) ;
    buf_clk cell_5591 ( .C ( clk ), .D ( signal_3535 ), .Q ( signal_11183 ) ) ;
    buf_clk cell_5649 ( .C ( clk ), .D ( signal_1589 ), .Q ( signal_11241 ) ) ;
    buf_clk cell_5659 ( .C ( clk ), .D ( signal_3702 ), .Q ( signal_11251 ) ) ;
    buf_clk cell_5669 ( .C ( clk ), .D ( signal_3703 ), .Q ( signal_11261 ) ) ;
    buf_clk cell_6255 ( .C ( clk ), .D ( signal_1527 ), .Q ( signal_11847 ) ) ;
    buf_clk cell_6269 ( .C ( clk ), .D ( signal_3578 ), .Q ( signal_11861 ) ) ;
    buf_clk cell_6283 ( .C ( clk ), .D ( signal_3579 ), .Q ( signal_11875 ) ) ;
    buf_clk cell_6321 ( .C ( clk ), .D ( signal_1633 ), .Q ( signal_11913 ) ) ;
    buf_clk cell_6335 ( .C ( clk ), .D ( signal_3790 ), .Q ( signal_11927 ) ) ;
    buf_clk cell_6349 ( .C ( clk ), .D ( signal_3791 ), .Q ( signal_11941 ) ) ;
    buf_clk cell_6441 ( .C ( clk ), .D ( signal_1588 ), .Q ( signal_12033 ) ) ;
    buf_clk cell_6457 ( .C ( clk ), .D ( signal_3700 ), .Q ( signal_12049 ) ) ;
    buf_clk cell_6473 ( .C ( clk ), .D ( signal_3701 ), .Q ( signal_12065 ) ) ;
    buf_clk cell_6501 ( .C ( clk ), .D ( signal_1602 ), .Q ( signal_12093 ) ) ;
    buf_clk cell_6517 ( .C ( clk ), .D ( signal_3728 ), .Q ( signal_12109 ) ) ;
    buf_clk cell_6533 ( .C ( clk ), .D ( signal_3729 ), .Q ( signal_12125 ) ) ;
    buf_clk cell_6735 ( .C ( clk ), .D ( signal_1539 ), .Q ( signal_12327 ) ) ;
    buf_clk cell_6753 ( .C ( clk ), .D ( signal_3602 ), .Q ( signal_12345 ) ) ;
    buf_clk cell_6771 ( .C ( clk ), .D ( signal_3603 ), .Q ( signal_12363 ) ) ;
    buf_clk cell_6885 ( .C ( clk ), .D ( signal_1603 ), .Q ( signal_12477 ) ) ;
    buf_clk cell_6905 ( .C ( clk ), .D ( signal_3730 ), .Q ( signal_12497 ) ) ;
    buf_clk cell_6925 ( .C ( clk ), .D ( signal_3731 ), .Q ( signal_12517 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1644 ( .a ({signal_3109, signal_3108, signal_1292}), .b ({signal_8420, signal_8418, signal_8416}), .clk ( clk ), .r ({Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({signal_3843, signal_3842, signal_1659}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1652 ( .a ({signal_8426, signal_8424, signal_8422}), .b ({signal_3295, signal_3294, signal_1385}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365]}), .c ({signal_3859, signal_3858, signal_1667}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1662 ( .a ({signal_8432, signal_8430, signal_8428}), .b ({signal_3183, signal_3182, signal_1329}), .clk ( clk ), .r ({Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({signal_3879, signal_3878, signal_1677}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1672 ( .a ({signal_8438, signal_8436, signal_8434}), .b ({signal_3211, signal_3210, signal_1343}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371]}), .c ({signal_3899, signal_3898, signal_1687}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1683 ( .a ({signal_8444, signal_8442, signal_8440}), .b ({signal_3241, signal_3240, signal_1358}), .clk ( clk ), .r ({Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({signal_3921, signal_3920, signal_1698}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1685 ( .a ({signal_8450, signal_8448, signal_8446}), .b ({signal_3245, signal_3244, signal_1360}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377]}), .c ({signal_3925, signal_3924, signal_1700}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1686 ( .a ({signal_8456, signal_8454, signal_8452}), .b ({signal_3417, signal_3416, signal_1446}), .clk ( clk ), .r ({Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_3927, signal_3926, signal_1701}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1688 ( .a ({signal_8462, signal_8460, signal_8458}), .b ({signal_3417, signal_3416, signal_1446}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383]}), .c ({signal_3931, signal_3930, signal_1703}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1689 ( .a ({signal_8462, signal_8460, signal_8458}), .b ({signal_3445, signal_3444, signal_1460}), .clk ( clk ), .r ({Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({signal_3933, signal_3932, signal_1704}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1690 ( .a ({signal_8468, signal_8466, signal_8464}), .b ({signal_3447, signal_3446, signal_1461}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389]}), .c ({signal_3935, signal_3934, signal_1705}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1691 ( .a ({signal_8474, signal_8472, signal_8470}), .b ({signal_3449, signal_3448, signal_1462}), .clk ( clk ), .r ({Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({signal_3937, signal_3936, signal_1706}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1692 ( .a ({signal_8480, signal_8478, signal_8476}), .b ({signal_3425, signal_3424, signal_1450}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395]}), .c ({signal_3939, signal_3938, signal_1707}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1694 ( .a ({signal_8498, signal_8492, signal_8486}), .b ({signal_3481, signal_3480, signal_1478}), .clk ( clk ), .r ({Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({signal_3943, signal_3942, signal_1709}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1695 ( .a ({signal_8504, signal_8502, signal_8500}), .b ({signal_3251, signal_3250, signal_1363}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401]}), .c ({signal_3945, signal_3944, signal_1710}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1696 ( .a ({signal_8510, signal_8508, signal_8506}), .b ({signal_3395, signal_3394, signal_1435}), .clk ( clk ), .r ({Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({signal_3947, signal_3946, signal_1711}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1697 ( .a ({signal_8516, signal_8514, signal_8512}), .b ({signal_3473, signal_3472, signal_1474}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407]}), .c ({signal_3949, signal_3948, signal_1712}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1699 ( .a ({signal_8522, signal_8520, signal_8518}), .b ({signal_3519, signal_3518, signal_1497}), .clk ( clk ), .r ({Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_3953, signal_3952, signal_1714}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1715 ( .a ({signal_3843, signal_3842, signal_1659}), .b ({signal_3985, signal_3984, signal_1730}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1721 ( .a ({signal_3859, signal_3858, signal_1667}), .b ({signal_3997, signal_3996, signal_1736}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1725 ( .a ({signal_3879, signal_3878, signal_1677}), .b ({signal_4005, signal_4004, signal_1740}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1737 ( .a ({signal_3925, signal_3924, signal_1700}), .b ({signal_4029, signal_4028, signal_1752}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1738 ( .a ({signal_3927, signal_3926, signal_1701}), .b ({signal_4031, signal_4030, signal_1753}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1740 ( .a ({signal_3931, signal_3930, signal_1703}), .b ({signal_4035, signal_4034, signal_1755}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1741 ( .a ({signal_3933, signal_3932, signal_1704}), .b ({signal_4037, signal_4036, signal_1756}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1742 ( .a ({signal_3935, signal_3934, signal_1705}), .b ({signal_4039, signal_4038, signal_1757}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1743 ( .a ({signal_3937, signal_3936, signal_1706}), .b ({signal_4041, signal_4040, signal_1758}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1744 ( .a ({signal_3939, signal_3938, signal_1707}), .b ({signal_4043, signal_4042, signal_1759}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1746 ( .a ({signal_3943, signal_3942, signal_1709}), .b ({signal_4047, signal_4046, signal_1761}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1747 ( .a ({signal_3947, signal_3946, signal_1711}), .b ({signal_4049, signal_4048, signal_1762}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1748 ( .a ({signal_3949, signal_3948, signal_1712}), .b ({signal_4051, signal_4050, signal_1763}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1750 ( .a ({signal_3953, signal_3952, signal_1714}), .b ({signal_4055, signal_4054, signal_1765}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1752 ( .a ({signal_3587, signal_3586, signal_1531}), .b ({signal_3589, signal_3588, signal_1532}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413]}), .c ({signal_4059, signal_4058, signal_1767}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1759 ( .a ({signal_8528, signal_8526, signal_8524}), .b ({signal_3549, signal_3548, signal_1512}), .clk ( clk ), .r ({Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({signal_4073, signal_4072, signal_1774}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1763 ( .a ({signal_8534, signal_8532, signal_8530}), .b ({signal_3559, signal_3558, signal_1517}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419]}), .c ({signal_4081, signal_4080, signal_1778}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1768 ( .a ({signal_3575, signal_3574, signal_1525}), .b ({signal_3577, signal_3576, signal_1526}), .clk ( clk ), .r ({Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({signal_4091, signal_4090, signal_1783}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1771 ( .a ({signal_3571, signal_3570, signal_1523}), .b ({signal_3585, signal_3584, signal_1530}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425]}), .c ({signal_4097, signal_4096, signal_1786}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1774 ( .a ({signal_8540, signal_8538, signal_8536}), .b ({signal_3597, signal_3596, signal_1536}), .clk ( clk ), .r ({Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({signal_4103, signal_4102, signal_1789}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1775 ( .a ({signal_3607, signal_3606, signal_1541}), .b ({signal_3609, signal_3608, signal_1542}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431]}), .c ({signal_4105, signal_4104, signal_1790}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1777 ( .a ({signal_8546, signal_8544, signal_8542}), .b ({signal_3617, signal_3616, signal_1546}), .clk ( clk ), .r ({Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({signal_4109, signal_4108, signal_1792}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1780 ( .a ({signal_8552, signal_8550, signal_8548}), .b ({signal_3823, signal_3822, signal_1649}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437]}), .c ({signal_4115, signal_4114, signal_1795}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1781 ( .a ({signal_3713, signal_3712, signal_1594}), .b ({signal_3747, signal_3746, signal_1611}), .clk ( clk ), .r ({Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_4117, signal_4116, signal_1796}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1787 ( .a ({signal_8558, signal_8556, signal_8554}), .b ({signal_3647, signal_3646, signal_1561}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443]}), .c ({signal_4129, signal_4128, signal_1802}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1788 ( .a ({signal_3651, signal_3650, signal_1563}), .b ({signal_8564, signal_8562, signal_8560}), .clk ( clk ), .r ({Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({signal_4131, signal_4130, signal_1803}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1789 ( .a ({signal_8570, signal_8568, signal_8566}), .b ({signal_3831, signal_3830, signal_1653}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449]}), .c ({signal_4133, signal_4132, signal_1804}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1790 ( .a ({signal_8576, signal_8574, signal_8572}), .b ({signal_3833, signal_3832, signal_1654}), .clk ( clk ), .r ({Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({signal_4135, signal_4134, signal_1805}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1791 ( .a ({signal_8582, signal_8580, signal_8578}), .b ({signal_3835, signal_3834, signal_1655}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455]}), .c ({signal_4137, signal_4136, signal_1806}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1792 ( .a ({signal_3657, signal_3656, signal_1566}), .b ({signal_3659, signal_3658, signal_1567}), .clk ( clk ), .r ({Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({signal_4139, signal_4138, signal_1807}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1793 ( .a ({signal_3099, signal_3098, signal_1287}), .b ({signal_3661, signal_3660, signal_1568}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461]}), .c ({signal_4141, signal_4140, signal_1808}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1794 ( .a ({signal_3805, signal_3804, signal_1640}), .b ({signal_3663, signal_3662, signal_1569}), .clk ( clk ), .r ({Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({signal_4143, signal_4142, signal_1809}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1795 ( .a ({signal_8468, signal_8466, signal_8464}), .b ({signal_3667, signal_3666, signal_1571}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467]}), .c ({signal_4145, signal_4144, signal_1810}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1796 ( .a ({signal_3551, signal_3550, signal_1513}), .b ({signal_3669, signal_3668, signal_1572}), .clk ( clk ), .r ({Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_4147, signal_4146, signal_1811}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1797 ( .a ({signal_8588, signal_8586, signal_8584}), .b ({signal_3671, signal_3670, signal_1573}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473]}), .c ({signal_4149, signal_4148, signal_1812}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1798 ( .a ({signal_8594, signal_8592, signal_8590}), .b ({signal_3845, signal_3844, signal_1660}), .clk ( clk ), .r ({Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({signal_4151, signal_4150, signal_1813}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1799 ( .a ({signal_8600, signal_8598, signal_8596}), .b ({signal_3673, signal_3672, signal_1574}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479]}), .c ({signal_4153, signal_4152, signal_1814}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1800 ( .a ({signal_8606, signal_8604, signal_8602}), .b ({signal_3679, signal_3678, signal_1577}), .clk ( clk ), .r ({Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({signal_4155, signal_4154, signal_1815}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1801 ( .a ({signal_8612, signal_8610, signal_8608}), .b ({signal_3847, signal_3846, signal_1661}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485]}), .c ({signal_4157, signal_4156, signal_1816}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1802 ( .a ({signal_8618, signal_8616, signal_8614}), .b ({signal_3657, signal_3656, signal_1566}), .clk ( clk ), .r ({Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({signal_4159, signal_4158, signal_1817}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1803 ( .a ({signal_3683, signal_3682, signal_1579}), .b ({signal_3685, signal_3684, signal_1580}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491]}), .c ({signal_4161, signal_4160, signal_1818}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1804 ( .a ({signal_3573, signal_3572, signal_1524}), .b ({signal_3695, signal_3694, signal_1585}), .clk ( clk ), .r ({Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({signal_4163, signal_4162, signal_1819}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1805 ( .a ({signal_3673, signal_3672, signal_1574}), .b ({signal_3697, signal_3696, signal_1586}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497]}), .c ({signal_4165, signal_4164, signal_1820}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1806 ( .a ({signal_8630, signal_8626, signal_8622}), .b ({signal_3861, signal_3860, signal_1668}), .clk ( clk ), .r ({Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_4167, signal_4166, signal_1821}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1807 ( .a ({signal_8636, signal_8634, signal_8632}), .b ({signal_3857, signal_3856, signal_1666}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503]}), .c ({signal_4169, signal_4168, signal_1822}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1808 ( .a ({signal_8642, signal_8640, signal_8638}), .b ({signal_3865, signal_3864, signal_1670}), .clk ( clk ), .r ({Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({signal_4171, signal_4170, signal_1823}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1809 ( .a ({signal_8654, signal_8650, signal_8646}), .b ({signal_3867, signal_3866, signal_1671}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509]}), .c ({signal_4173, signal_4172, signal_1824}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1810 ( .a ({signal_3783, signal_3782, signal_1629}), .b ({signal_3785, signal_3784, signal_1630}), .clk ( clk ), .r ({Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({signal_4175, signal_4174, signal_1825}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1811 ( .a ({signal_3583, signal_3582, signal_1529}), .b ({signal_3869, signal_3868, signal_1672}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515]}), .c ({signal_4177, signal_4176, signal_1826}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1812 ( .a ({signal_3601, signal_3600, signal_1538}), .b ({signal_3723, signal_3722, signal_1599}), .clk ( clk ), .r ({Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({signal_4179, signal_4178, signal_1827}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1813 ( .a ({signal_3613, signal_3612, signal_1544}), .b ({signal_3735, signal_3734, signal_1605}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521]}), .c ({signal_4181, signal_4180, signal_1828}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1814 ( .a ({signal_3615, signal_3614, signal_1545}), .b ({signal_3739, signal_3738, signal_1607}), .clk ( clk ), .r ({Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({signal_4183, signal_4182, signal_1829}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1815 ( .a ({signal_8660, signal_8658, signal_8656}), .b ({signal_3741, signal_3740, signal_1608}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527]}), .c ({signal_4185, signal_4184, signal_1830}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1816 ( .a ({signal_8666, signal_8664, signal_8662}), .b ({signal_3893, signal_3892, signal_1684}), .clk ( clk ), .r ({Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_4187, signal_4186, signal_1831}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1817 ( .a ({signal_8672, signal_8670, signal_8668}), .b ({signal_3895, signal_3894, signal_1685}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533]}), .c ({signal_4189, signal_4188, signal_1832}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1818 ( .a ({signal_3667, signal_3666, signal_1571}), .b ({signal_3717, signal_3716, signal_1596}), .clk ( clk ), .r ({Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({signal_4191, signal_4190, signal_1833}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1820 ( .a ({signal_3213, signal_3212, signal_1344}), .b ({signal_3745, signal_3744, signal_1610}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539]}), .c ({signal_4195, signal_4194, signal_1835}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1821 ( .a ({signal_8678, signal_8676, signal_8674}), .b ({signal_3749, signal_3748, signal_1612}), .clk ( clk ), .r ({Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({signal_4197, signal_4196, signal_1836}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1822 ( .a ({signal_8684, signal_8682, signal_8680}), .b ({signal_3755, signal_3754, signal_1615}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545]}), .c ({signal_4199, signal_4198, signal_1837}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1823 ( .a ({signal_3637, signal_3636, signal_1556}), .b ({signal_3759, signal_3758, signal_1617}), .clk ( clk ), .r ({Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({signal_4201, signal_4200, signal_1838}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1824 ( .a ({signal_8690, signal_8688, signal_8686}), .b ({signal_3909, signal_3908, signal_1692}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551]}), .c ({signal_4203, signal_4202, signal_1839}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1825 ( .a ({signal_8696, signal_8694, signal_8692}), .b ({signal_3765, signal_3764, signal_1620}), .clk ( clk ), .r ({Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({signal_4205, signal_4204, signal_1840}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1826 ( .a ({signal_8702, signal_8700, signal_8698}), .b ({signal_3755, signal_3754, signal_1615}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557]}), .c ({signal_4207, signal_4206, signal_1841}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1827 ( .a ({signal_8708, signal_8706, signal_8704}), .b ({signal_3915, signal_3914, signal_1695}), .clk ( clk ), .r ({Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_4209, signal_4208, signal_1842}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1828 ( .a ({signal_3653, signal_3652, signal_1564}), .b ({signal_3771, signal_3770, signal_1623}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563]}), .c ({signal_4211, signal_4210, signal_1843}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1829 ( .a ({signal_8714, signal_8712, signal_8710}), .b ({signal_3773, signal_3772, signal_1624}), .clk ( clk ), .r ({Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({signal_4213, signal_4212, signal_1844}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1830 ( .a ({signal_3777, signal_3776, signal_1626}), .b ({signal_3779, signal_3778, signal_1627}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569]}), .c ({signal_4215, signal_4214, signal_1845}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1831 ( .a ({signal_3709, signal_3708, signal_1592}), .b ({signal_3781, signal_3780, signal_1628}), .clk ( clk ), .r ({Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({signal_4217, signal_4216, signal_1846}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1832 ( .a ({signal_3571, signal_3570, signal_1523}), .b ({signal_3793, signal_3792, signal_1634}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575]}), .c ({signal_4219, signal_4218, signal_1847}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1833 ( .a ({signal_3249, signal_3248, signal_1362}), .b ({signal_3795, signal_3794, signal_1635}), .clk ( clk ), .r ({Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({signal_4221, signal_4220, signal_1848}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1842 ( .a ({signal_4081, signal_4080, signal_1778}), .b ({signal_4239, signal_4238, signal_1857}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1853 ( .a ({signal_4115, signal_4114, signal_1795}), .b ({signal_4261, signal_4260, signal_1868}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1859 ( .a ({signal_4135, signal_4134, signal_1805}), .b ({signal_4273, signal_4272, signal_1874}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1860 ( .a ({signal_4139, signal_4138, signal_1807}), .b ({signal_4275, signal_4274, signal_1875}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1861 ( .a ({signal_4149, signal_4148, signal_1812}), .b ({signal_4277, signal_4276, signal_1876}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1862 ( .a ({signal_4157, signal_4156, signal_1816}), .b ({signal_4279, signal_4278, signal_1877}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1863 ( .a ({signal_4159, signal_4158, signal_1817}), .b ({signal_4281, signal_4280, signal_1878}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1864 ( .a ({signal_4167, signal_4166, signal_1821}), .b ({signal_4283, signal_4282, signal_1879}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1865 ( .a ({signal_4169, signal_4168, signal_1822}), .b ({signal_4285, signal_4284, signal_1880}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1866 ( .a ({signal_4171, signal_4170, signal_1823}), .b ({signal_4287, signal_4286, signal_1881}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1867 ( .a ({signal_4173, signal_4172, signal_1824}), .b ({signal_4289, signal_4288, signal_1882}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1868 ( .a ({signal_4181, signal_4180, signal_1828}), .b ({signal_4291, signal_4290, signal_1883}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1869 ( .a ({signal_4183, signal_4182, signal_1829}), .b ({signal_4293, signal_4292, signal_1884}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1870 ( .a ({signal_4187, signal_4186, signal_1831}), .b ({signal_4295, signal_4294, signal_1885}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1871 ( .a ({signal_4189, signal_4188, signal_1832}), .b ({signal_4297, signal_4296, signal_1886}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1873 ( .a ({signal_4209, signal_4208, signal_1842}), .b ({signal_4301, signal_4300, signal_1888}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1874 ( .a ({signal_4213, signal_4212, signal_1844}), .b ({signal_4303, signal_4302, signal_1889}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1876 ( .a ({signal_3955, signal_3954, signal_1715}), .b ({signal_8720, signal_8718, signal_8716}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581]}), .c ({signal_4307, signal_4306, signal_1891}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1877 ( .a ({signal_8732, signal_8728, signal_8724}), .b ({signal_3957, signal_3956, signal_1716}), .clk ( clk ), .r ({Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({signal_4309, signal_4308, signal_1892}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1878 ( .a ({signal_8738, signal_8736, signal_8734}), .b ({signal_3959, signal_3958, signal_1717}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587]}), .c ({signal_4311, signal_4310, signal_1893}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1879 ( .a ({signal_8462, signal_8460, signal_8458}), .b ({signal_3961, signal_3960, signal_1718}), .clk ( clk ), .r ({Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_4313, signal_4312, signal_1894}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1880 ( .a ({signal_8522, signal_8520, signal_8518}), .b ({signal_4061, signal_4060, signal_1768}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593]}), .c ({signal_4315, signal_4314, signal_1895}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1881 ( .a ({signal_8750, signal_8746, signal_8742}), .b ({signal_3963, signal_3962, signal_1719}), .clk ( clk ), .r ({Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({signal_4317, signal_4316, signal_1896}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1882 ( .a ({signal_3965, signal_3964, signal_1720}), .b ({signal_8756, signal_8754, signal_8752}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599]}), .c ({signal_4319, signal_4318, signal_1897}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1883 ( .a ({signal_8762, signal_8760, signal_8758}), .b ({signal_3967, signal_3966, signal_1721}), .clk ( clk ), .r ({Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({signal_4321, signal_4320, signal_1898}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1884 ( .a ({signal_8768, signal_8766, signal_8764}), .b ({signal_3969, signal_3968, signal_1722}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605]}), .c ({signal_4323, signal_4322, signal_1899}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1885 ( .a ({signal_8786, signal_8780, signal_8774}), .b ({signal_3971, signal_3970, signal_1723}), .clk ( clk ), .r ({Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({signal_4325, signal_4324, signal_1900}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1886 ( .a ({signal_8480, signal_8478, signal_8476}), .b ({signal_4063, signal_4062, signal_1769}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611]}), .c ({signal_4327, signal_4326, signal_1901}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1887 ( .a ({signal_8792, signal_8790, signal_8788}), .b ({signal_3973, signal_3972, signal_1724}), .clk ( clk ), .r ({Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({signal_4329, signal_4328, signal_1902}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1888 ( .a ({signal_8798, signal_8796, signal_8794}), .b ({signal_3977, signal_3976, signal_1726}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617]}), .c ({signal_4331, signal_4330, signal_1903}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1889 ( .a ({signal_8804, signal_8802, signal_8800}), .b ({signal_4067, signal_4066, signal_1771}), .clk ( clk ), .r ({Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_4333, signal_4332, signal_1904}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1890 ( .a ({signal_8462, signal_8460, signal_8458}), .b ({signal_3979, signal_3978, signal_1727}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623]}), .c ({signal_4335, signal_4334, signal_1905}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1891 ( .a ({signal_8522, signal_8520, signal_8518}), .b ({signal_3981, signal_3980, signal_1728}), .clk ( clk ), .r ({Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({signal_4337, signal_4336, signal_1906}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1892 ( .a ({signal_8810, signal_8808, signal_8806}), .b ({signal_3983, signal_3982, signal_1729}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629]}), .c ({signal_4339, signal_4338, signal_1907}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1894 ( .a ({signal_8534, signal_8532, signal_8530}), .b ({signal_3987, signal_3986, signal_1731}), .clk ( clk ), .r ({Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({signal_4343, signal_4342, signal_1909}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1895 ( .a ({signal_8822, signal_8818, signal_8814}), .b ({signal_3989, signal_3988, signal_1732}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635]}), .c ({signal_4345, signal_4344, signal_1910}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1896 ( .a ({signal_8828, signal_8826, signal_8824}), .b ({signal_3991, signal_3990, signal_1733}), .clk ( clk ), .r ({Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({signal_4347, signal_4346, signal_1911}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1897 ( .a ({signal_8834, signal_8832, signal_8830}), .b ({signal_3993, signal_3992, signal_1734}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641]}), .c ({signal_4349, signal_4348, signal_1912}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1898 ( .a ({signal_8840, signal_8838, signal_8836}), .b ({signal_4089, signal_4088, signal_1782}), .clk ( clk ), .r ({Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({signal_4351, signal_4350, signal_1913}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1899 ( .a ({signal_8846, signal_8844, signal_8842}), .b ({signal_3995, signal_3994, signal_1735}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647]}), .c ({signal_4353, signal_4352, signal_1914}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1900 ( .a ({signal_8798, signal_8796, signal_8794}), .b ({signal_3999, signal_3998, signal_1737}), .clk ( clk ), .r ({Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_4355, signal_4354, signal_1915}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1901 ( .a ({signal_4001, signal_4000, signal_1738}), .b ({signal_3873, signal_3872, signal_1674}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653]}), .c ({signal_4357, signal_4356, signal_1916}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1903 ( .a ({signal_8468, signal_8466, signal_8464}), .b ({signal_4003, signal_4002, signal_1739}), .clk ( clk ), .r ({Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({signal_4361, signal_4360, signal_1918}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1905 ( .a ({signal_8828, signal_8826, signal_8824}), .b ({signal_4007, signal_4006, signal_1741}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659]}), .c ({signal_4365, signal_4364, signal_1920}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1906 ( .a ({signal_8516, signal_8514, signal_8512}), .b ({signal_4009, signal_4008, signal_1742}), .clk ( clk ), .r ({Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({signal_4367, signal_4366, signal_1921}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1907 ( .a ({signal_8666, signal_8664, signal_8662}), .b ({signal_4011, signal_4010, signal_1743}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665]}), .c ({signal_4369, signal_4368, signal_1922}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1908 ( .a ({signal_8750, signal_8746, signal_8742}), .b ({signal_4013, signal_4012, signal_1744}), .clk ( clk ), .r ({Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({signal_4371, signal_4370, signal_1923}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1909 ( .a ({signal_8852, signal_8850, signal_8848}), .b ({signal_4089, signal_4088, signal_1782}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671]}), .c ({signal_4373, signal_4372, signal_1924}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1910 ( .a ({signal_8858, signal_8856, signal_8854}), .b ({signal_4015, signal_4014, signal_1745}), .clk ( clk ), .r ({Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({signal_4375, signal_4374, signal_1925}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1913 ( .a ({signal_8864, signal_8862, signal_8860}), .b ({signal_4017, signal_4016, signal_1746}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677]}), .c ({signal_4381, signal_4380, signal_1928}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1914 ( .a ({signal_8516, signal_8514, signal_8512}), .b ({signal_4019, signal_4018, signal_1747}), .clk ( clk ), .r ({Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_4383, signal_4382, signal_1929}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1915 ( .a ({signal_8462, signal_8460, signal_8458}), .b ({signal_4021, signal_4020, signal_1748}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683]}), .c ({signal_4385, signal_4384, signal_1930}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1916 ( .a ({signal_8870, signal_8868, signal_8866}), .b ({signal_3975, signal_3974, signal_1725}), .clk ( clk ), .r ({Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({signal_4387, signal_4386, signal_1931}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1917 ( .a ({signal_8876, signal_8874, signal_8872}), .b ({signal_3983, signal_3982, signal_1729}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689]}), .c ({signal_4389, signal_4388, signal_1932}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1919 ( .a ({signal_8888, signal_8884, signal_8880}), .b ({signal_4023, signal_4022, signal_1749}), .clk ( clk ), .r ({Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({signal_4393, signal_4392, signal_1934}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1920 ( .a ({signal_8666, signal_8664, signal_8662}), .b ({signal_4025, signal_4024, signal_1750}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695]}), .c ({signal_4395, signal_4394, signal_1935}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1923 ( .a ({signal_8894, signal_8892, signal_8890}), .b ({signal_4027, signal_4026, signal_1751}), .clk ( clk ), .r ({Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({signal_4401, signal_4400, signal_1938}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1927 ( .a ({signal_8900, signal_8898, signal_8896}), .b ({signal_4033, signal_4032, signal_1754}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701]}), .c ({signal_4409, signal_4408, signal_1942}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1932 ( .a ({signal_8456, signal_8454, signal_8452}), .b ({signal_4045, signal_4044, signal_1760}), .clk ( clk ), .r ({Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({signal_4419, signal_4418, signal_1947}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1944 ( .a ({signal_8906, signal_8904, signal_8902}), .b ({signal_4053, signal_4052, signal_1764}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707]}), .c ({signal_4443, signal_4442, signal_1959}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1948 ( .a ({signal_4309, signal_4308, signal_1892}), .b ({signal_4451, signal_4450, signal_1963}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1949 ( .a ({signal_4311, signal_4310, signal_1893}), .b ({signal_4453, signal_4452, signal_1964}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1950 ( .a ({signal_4315, signal_4314, signal_1895}), .b ({signal_4455, signal_4454, signal_1965}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1951 ( .a ({signal_4319, signal_4318, signal_1897}), .b ({signal_4457, signal_4456, signal_1966}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1952 ( .a ({signal_4321, signal_4320, signal_1898}), .b ({signal_4459, signal_4458, signal_1967}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1953 ( .a ({signal_4325, signal_4324, signal_1900}), .b ({signal_4461, signal_4460, signal_1968}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1954 ( .a ({signal_4327, signal_4326, signal_1901}), .b ({signal_4463, signal_4462, signal_1969}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1955 ( .a ({signal_4329, signal_4328, signal_1902}), .b ({signal_4465, signal_4464, signal_1970}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1956 ( .a ({signal_4331, signal_4330, signal_1903}), .b ({signal_4467, signal_4466, signal_1971}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1957 ( .a ({signal_4333, signal_4332, signal_1904}), .b ({signal_4469, signal_4468, signal_1972}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1958 ( .a ({signal_4335, signal_4334, signal_1905}), .b ({signal_4471, signal_4470, signal_1973}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1959 ( .a ({signal_4337, signal_4336, signal_1906}), .b ({signal_4473, signal_4472, signal_1974}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1960 ( .a ({signal_4339, signal_4338, signal_1907}), .b ({signal_4475, signal_4474, signal_1975}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1962 ( .a ({signal_4343, signal_4342, signal_1909}), .b ({signal_4479, signal_4478, signal_1977}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1963 ( .a ({signal_4345, signal_4344, signal_1910}), .b ({signal_4481, signal_4480, signal_1978}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1964 ( .a ({signal_4347, signal_4346, signal_1911}), .b ({signal_4483, signal_4482, signal_1979}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1965 ( .a ({signal_4349, signal_4348, signal_1912}), .b ({signal_4485, signal_4484, signal_1980}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1966 ( .a ({signal_4351, signal_4350, signal_1913}), .b ({signal_4487, signal_4486, signal_1981}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1967 ( .a ({signal_4353, signal_4352, signal_1914}), .b ({signal_4489, signal_4488, signal_1982}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1968 ( .a ({signal_4355, signal_4354, signal_1915}), .b ({signal_4491, signal_4490, signal_1983}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1970 ( .a ({signal_4361, signal_4360, signal_1918}), .b ({signal_4495, signal_4494, signal_1985}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1972 ( .a ({signal_4365, signal_4364, signal_1920}), .b ({signal_4499, signal_4498, signal_1987}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1973 ( .a ({signal_4367, signal_4366, signal_1921}), .b ({signal_4501, signal_4500, signal_1988}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1974 ( .a ({signal_4369, signal_4368, signal_1922}), .b ({signal_4503, signal_4502, signal_1989}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1975 ( .a ({signal_4371, signal_4370, signal_1923}), .b ({signal_4505, signal_4504, signal_1990}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1976 ( .a ({signal_4373, signal_4372, signal_1924}), .b ({signal_4507, signal_4506, signal_1991}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1977 ( .a ({signal_4375, signal_4374, signal_1925}), .b ({signal_4509, signal_4508, signal_1992}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1979 ( .a ({signal_4381, signal_4380, signal_1928}), .b ({signal_4513, signal_4512, signal_1994}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1980 ( .a ({signal_4383, signal_4382, signal_1929}), .b ({signal_4515, signal_4514, signal_1995}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1981 ( .a ({signal_4385, signal_4384, signal_1930}), .b ({signal_4517, signal_4516, signal_1996}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1982 ( .a ({signal_4387, signal_4386, signal_1931}), .b ({signal_4519, signal_4518, signal_1997}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1983 ( .a ({signal_4389, signal_4388, signal_1932}), .b ({signal_4521, signal_4520, signal_1998}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1984 ( .a ({signal_4393, signal_4392, signal_1934}), .b ({signal_4523, signal_4522, signal_1999}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1985 ( .a ({signal_4395, signal_4394, signal_1935}), .b ({signal_4525, signal_4524, signal_2000}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1988 ( .a ({signal_4401, signal_4400, signal_1938}), .b ({signal_4531, signal_4530, signal_2003}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1990 ( .a ({signal_4409, signal_4408, signal_1942}), .b ({signal_4535, signal_4534, signal_2005}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1991 ( .a ({signal_4419, signal_4418, signal_1947}), .b ({signal_4537, signal_4536, signal_2006}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1996 ( .a ({signal_4443, signal_4442, signal_1959}), .b ({signal_4547, signal_4546, signal_2011}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2000 ( .a ({signal_4251, signal_4250, signal_1863}), .b ({signal_3713, signal_3712, signal_1594}), .clk ( clk ), .r ({Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_4555, signal_4554, signal_2015}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2001 ( .a ({signal_4229, signal_4228, signal_1852}), .b ({signal_3655, signal_3654, signal_1565}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713]}), .c ({signal_4557, signal_4556, signal_2016}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2003 ( .a ({signal_4235, signal_4234, signal_1855}), .b ({signal_4237, signal_4236, signal_1856}), .clk ( clk ), .r ({Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({signal_4561, signal_4560, signal_2018}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2004 ( .a ({signal_8912, signal_8910, signal_8908}), .b ({signal_4241, signal_4240, signal_1858}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719]}), .c ({signal_4563, signal_4562, signal_2019}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2005 ( .a ({signal_8678, signal_8676, signal_8674}), .b ({signal_4243, signal_4242, signal_1859}), .clk ( clk ), .r ({Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({signal_4565, signal_4564, signal_2020}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2006 ( .a ({signal_8918, signal_8916, signal_8914}), .b ({signal_4245, signal_4244, signal_1860}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725]}), .c ({signal_4567, signal_4566, signal_2021}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2008 ( .a ({signal_8924, signal_8922, signal_8920}), .b ({signal_4253, signal_4252, signal_1864}), .clk ( clk ), .r ({Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({signal_4571, signal_4570, signal_2023}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2011 ( .a ({signal_8678, signal_8676, signal_8674}), .b ({signal_4255, signal_4254, signal_1865}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731]}), .c ({signal_4577, signal_4576, signal_2026}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2012 ( .a ({signal_3743, signal_3742, signal_1609}), .b ({signal_4259, signal_4258, signal_1867}), .clk ( clk ), .r ({Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({signal_4579, signal_4578, signal_2027}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2014 ( .a ({signal_4263, signal_4262, signal_1869}), .b ({signal_3901, signal_3900, signal_1688}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737]}), .c ({signal_4583, signal_4582, signal_2029}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2015 ( .a ({signal_3739, signal_3738, signal_1607}), .b ({signal_4267, signal_4266, signal_1871}), .clk ( clk ), .r ({Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_4585, signal_4584, signal_2030}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2048 ( .a ({signal_4563, signal_4562, signal_2019}), .b ({signal_4651, signal_4650, signal_2063}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2052 ( .a ({signal_4577, signal_4576, signal_2026}), .b ({signal_4659, signal_4658, signal_2067}) ) ;
    buf_clk cell_3334 ( .C ( clk ), .D ( signal_8925 ), .Q ( signal_8926 ) ) ;
    buf_clk cell_3336 ( .C ( clk ), .D ( signal_8927 ), .Q ( signal_8928 ) ) ;
    buf_clk cell_3338 ( .C ( clk ), .D ( signal_8929 ), .Q ( signal_8930 ) ) ;
    buf_clk cell_3340 ( .C ( clk ), .D ( signal_8931 ), .Q ( signal_8932 ) ) ;
    buf_clk cell_3342 ( .C ( clk ), .D ( signal_8933 ), .Q ( signal_8934 ) ) ;
    buf_clk cell_3344 ( .C ( clk ), .D ( signal_8935 ), .Q ( signal_8936 ) ) ;
    buf_clk cell_3348 ( .C ( clk ), .D ( signal_8939 ), .Q ( signal_8940 ) ) ;
    buf_clk cell_3352 ( .C ( clk ), .D ( signal_8943 ), .Q ( signal_8944 ) ) ;
    buf_clk cell_3356 ( .C ( clk ), .D ( signal_8947 ), .Q ( signal_8948 ) ) ;
    buf_clk cell_3358 ( .C ( clk ), .D ( signal_8949 ), .Q ( signal_8950 ) ) ;
    buf_clk cell_3360 ( .C ( clk ), .D ( signal_8951 ), .Q ( signal_8952 ) ) ;
    buf_clk cell_3362 ( .C ( clk ), .D ( signal_8953 ), .Q ( signal_8954 ) ) ;
    buf_clk cell_3366 ( .C ( clk ), .D ( signal_8957 ), .Q ( signal_8958 ) ) ;
    buf_clk cell_3370 ( .C ( clk ), .D ( signal_8961 ), .Q ( signal_8962 ) ) ;
    buf_clk cell_3374 ( .C ( clk ), .D ( signal_8965 ), .Q ( signal_8966 ) ) ;
    buf_clk cell_3378 ( .C ( clk ), .D ( signal_8969 ), .Q ( signal_8970 ) ) ;
    buf_clk cell_3382 ( .C ( clk ), .D ( signal_8973 ), .Q ( signal_8974 ) ) ;
    buf_clk cell_3386 ( .C ( clk ), .D ( signal_8977 ), .Q ( signal_8978 ) ) ;
    buf_clk cell_3390 ( .C ( clk ), .D ( signal_8981 ), .Q ( signal_8982 ) ) ;
    buf_clk cell_3394 ( .C ( clk ), .D ( signal_8985 ), .Q ( signal_8986 ) ) ;
    buf_clk cell_3398 ( .C ( clk ), .D ( signal_8989 ), .Q ( signal_8990 ) ) ;
    buf_clk cell_3406 ( .C ( clk ), .D ( signal_8997 ), .Q ( signal_8998 ) ) ;
    buf_clk cell_3414 ( .C ( clk ), .D ( signal_9005 ), .Q ( signal_9006 ) ) ;
    buf_clk cell_3422 ( .C ( clk ), .D ( signal_9013 ), .Q ( signal_9014 ) ) ;
    buf_clk cell_3424 ( .C ( clk ), .D ( signal_9015 ), .Q ( signal_9016 ) ) ;
    buf_clk cell_3426 ( .C ( clk ), .D ( signal_9017 ), .Q ( signal_9018 ) ) ;
    buf_clk cell_3428 ( .C ( clk ), .D ( signal_9019 ), .Q ( signal_9020 ) ) ;
    buf_clk cell_3430 ( .C ( clk ), .D ( signal_9021 ), .Q ( signal_9022 ) ) ;
    buf_clk cell_3432 ( .C ( clk ), .D ( signal_9023 ), .Q ( signal_9024 ) ) ;
    buf_clk cell_3434 ( .C ( clk ), .D ( signal_9025 ), .Q ( signal_9026 ) ) ;
    buf_clk cell_3438 ( .C ( clk ), .D ( signal_9029 ), .Q ( signal_9030 ) ) ;
    buf_clk cell_3442 ( .C ( clk ), .D ( signal_9033 ), .Q ( signal_9034 ) ) ;
    buf_clk cell_3446 ( .C ( clk ), .D ( signal_9037 ), .Q ( signal_9038 ) ) ;
    buf_clk cell_3448 ( .C ( clk ), .D ( signal_9039 ), .Q ( signal_9040 ) ) ;
    buf_clk cell_3450 ( .C ( clk ), .D ( signal_9041 ), .Q ( signal_9042 ) ) ;
    buf_clk cell_3452 ( .C ( clk ), .D ( signal_9043 ), .Q ( signal_9044 ) ) ;
    buf_clk cell_3454 ( .C ( clk ), .D ( signal_9045 ), .Q ( signal_9046 ) ) ;
    buf_clk cell_3456 ( .C ( clk ), .D ( signal_9047 ), .Q ( signal_9048 ) ) ;
    buf_clk cell_3458 ( .C ( clk ), .D ( signal_9049 ), .Q ( signal_9050 ) ) ;
    buf_clk cell_3462 ( .C ( clk ), .D ( signal_9053 ), .Q ( signal_9054 ) ) ;
    buf_clk cell_3466 ( .C ( clk ), .D ( signal_9057 ), .Q ( signal_9058 ) ) ;
    buf_clk cell_3470 ( .C ( clk ), .D ( signal_9061 ), .Q ( signal_9062 ) ) ;
    buf_clk cell_3472 ( .C ( clk ), .D ( signal_9063 ), .Q ( signal_9064 ) ) ;
    buf_clk cell_3474 ( .C ( clk ), .D ( signal_9065 ), .Q ( signal_9066 ) ) ;
    buf_clk cell_3476 ( .C ( clk ), .D ( signal_9067 ), .Q ( signal_9068 ) ) ;
    buf_clk cell_3478 ( .C ( clk ), .D ( signal_9069 ), .Q ( signal_9070 ) ) ;
    buf_clk cell_3480 ( .C ( clk ), .D ( signal_9071 ), .Q ( signal_9072 ) ) ;
    buf_clk cell_3482 ( .C ( clk ), .D ( signal_9073 ), .Q ( signal_9074 ) ) ;
    buf_clk cell_3484 ( .C ( clk ), .D ( signal_9075 ), .Q ( signal_9076 ) ) ;
    buf_clk cell_3486 ( .C ( clk ), .D ( signal_9077 ), .Q ( signal_9078 ) ) ;
    buf_clk cell_3488 ( .C ( clk ), .D ( signal_9079 ), .Q ( signal_9080 ) ) ;
    buf_clk cell_3490 ( .C ( clk ), .D ( signal_9081 ), .Q ( signal_9082 ) ) ;
    buf_clk cell_3492 ( .C ( clk ), .D ( signal_9083 ), .Q ( signal_9084 ) ) ;
    buf_clk cell_3494 ( .C ( clk ), .D ( signal_9085 ), .Q ( signal_9086 ) ) ;
    buf_clk cell_3496 ( .C ( clk ), .D ( signal_9087 ), .Q ( signal_9088 ) ) ;
    buf_clk cell_3498 ( .C ( clk ), .D ( signal_9089 ), .Q ( signal_9090 ) ) ;
    buf_clk cell_3500 ( .C ( clk ), .D ( signal_9091 ), .Q ( signal_9092 ) ) ;
    buf_clk cell_3504 ( .C ( clk ), .D ( signal_9095 ), .Q ( signal_9096 ) ) ;
    buf_clk cell_3508 ( .C ( clk ), .D ( signal_9099 ), .Q ( signal_9100 ) ) ;
    buf_clk cell_3512 ( .C ( clk ), .D ( signal_9103 ), .Q ( signal_9104 ) ) ;
    buf_clk cell_3514 ( .C ( clk ), .D ( signal_9105 ), .Q ( signal_9106 ) ) ;
    buf_clk cell_3516 ( .C ( clk ), .D ( signal_9107 ), .Q ( signal_9108 ) ) ;
    buf_clk cell_3518 ( .C ( clk ), .D ( signal_9109 ), .Q ( signal_9110 ) ) ;
    buf_clk cell_3520 ( .C ( clk ), .D ( signal_9111 ), .Q ( signal_9112 ) ) ;
    buf_clk cell_3522 ( .C ( clk ), .D ( signal_9113 ), .Q ( signal_9114 ) ) ;
    buf_clk cell_3524 ( .C ( clk ), .D ( signal_9115 ), .Q ( signal_9116 ) ) ;
    buf_clk cell_3526 ( .C ( clk ), .D ( signal_9117 ), .Q ( signal_9118 ) ) ;
    buf_clk cell_3528 ( .C ( clk ), .D ( signal_9119 ), .Q ( signal_9120 ) ) ;
    buf_clk cell_3530 ( .C ( clk ), .D ( signal_9121 ), .Q ( signal_9122 ) ) ;
    buf_clk cell_3532 ( .C ( clk ), .D ( signal_9123 ), .Q ( signal_9124 ) ) ;
    buf_clk cell_3534 ( .C ( clk ), .D ( signal_9125 ), .Q ( signal_9126 ) ) ;
    buf_clk cell_3536 ( .C ( clk ), .D ( signal_9127 ), .Q ( signal_9128 ) ) ;
    buf_clk cell_3540 ( .C ( clk ), .D ( signal_9131 ), .Q ( signal_9132 ) ) ;
    buf_clk cell_3544 ( .C ( clk ), .D ( signal_9135 ), .Q ( signal_9136 ) ) ;
    buf_clk cell_3548 ( .C ( clk ), .D ( signal_9139 ), .Q ( signal_9140 ) ) ;
    buf_clk cell_3550 ( .C ( clk ), .D ( signal_9141 ), .Q ( signal_9142 ) ) ;
    buf_clk cell_3552 ( .C ( clk ), .D ( signal_9143 ), .Q ( signal_9144 ) ) ;
    buf_clk cell_3554 ( .C ( clk ), .D ( signal_9145 ), .Q ( signal_9146 ) ) ;
    buf_clk cell_3556 ( .C ( clk ), .D ( signal_9147 ), .Q ( signal_9148 ) ) ;
    buf_clk cell_3558 ( .C ( clk ), .D ( signal_9149 ), .Q ( signal_9150 ) ) ;
    buf_clk cell_3560 ( .C ( clk ), .D ( signal_9151 ), .Q ( signal_9152 ) ) ;
    buf_clk cell_3564 ( .C ( clk ), .D ( signal_9155 ), .Q ( signal_9156 ) ) ;
    buf_clk cell_3568 ( .C ( clk ), .D ( signal_9159 ), .Q ( signal_9160 ) ) ;
    buf_clk cell_3572 ( .C ( clk ), .D ( signal_9163 ), .Q ( signal_9164 ) ) ;
    buf_clk cell_3576 ( .C ( clk ), .D ( signal_9167 ), .Q ( signal_9168 ) ) ;
    buf_clk cell_3580 ( .C ( clk ), .D ( signal_9171 ), .Q ( signal_9172 ) ) ;
    buf_clk cell_3584 ( .C ( clk ), .D ( signal_9175 ), .Q ( signal_9176 ) ) ;
    buf_clk cell_3588 ( .C ( clk ), .D ( signal_9179 ), .Q ( signal_9180 ) ) ;
    buf_clk cell_3592 ( .C ( clk ), .D ( signal_9183 ), .Q ( signal_9184 ) ) ;
    buf_clk cell_3596 ( .C ( clk ), .D ( signal_9187 ), .Q ( signal_9188 ) ) ;
    buf_clk cell_3600 ( .C ( clk ), .D ( signal_9191 ), .Q ( signal_9192 ) ) ;
    buf_clk cell_3604 ( .C ( clk ), .D ( signal_9195 ), .Q ( signal_9196 ) ) ;
    buf_clk cell_3608 ( .C ( clk ), .D ( signal_9199 ), .Q ( signal_9200 ) ) ;
    buf_clk cell_3610 ( .C ( clk ), .D ( signal_9201 ), .Q ( signal_9202 ) ) ;
    buf_clk cell_3612 ( .C ( clk ), .D ( signal_9203 ), .Q ( signal_9204 ) ) ;
    buf_clk cell_3614 ( .C ( clk ), .D ( signal_9205 ), .Q ( signal_9206 ) ) ;
    buf_clk cell_3616 ( .C ( clk ), .D ( signal_9207 ), .Q ( signal_9208 ) ) ;
    buf_clk cell_3618 ( .C ( clk ), .D ( signal_9209 ), .Q ( signal_9210 ) ) ;
    buf_clk cell_3620 ( .C ( clk ), .D ( signal_9211 ), .Q ( signal_9212 ) ) ;
    buf_clk cell_3622 ( .C ( clk ), .D ( signal_9213 ), .Q ( signal_9214 ) ) ;
    buf_clk cell_3624 ( .C ( clk ), .D ( signal_9215 ), .Q ( signal_9216 ) ) ;
    buf_clk cell_3626 ( .C ( clk ), .D ( signal_9217 ), .Q ( signal_9218 ) ) ;
    buf_clk cell_3628 ( .C ( clk ), .D ( signal_9219 ), .Q ( signal_9220 ) ) ;
    buf_clk cell_3630 ( .C ( clk ), .D ( signal_9221 ), .Q ( signal_9222 ) ) ;
    buf_clk cell_3632 ( .C ( clk ), .D ( signal_9223 ), .Q ( signal_9224 ) ) ;
    buf_clk cell_3634 ( .C ( clk ), .D ( signal_9225 ), .Q ( signal_9226 ) ) ;
    buf_clk cell_3636 ( .C ( clk ), .D ( signal_9227 ), .Q ( signal_9228 ) ) ;
    buf_clk cell_3638 ( .C ( clk ), .D ( signal_9229 ), .Q ( signal_9230 ) ) ;
    buf_clk cell_3642 ( .C ( clk ), .D ( signal_9233 ), .Q ( signal_9234 ) ) ;
    buf_clk cell_3646 ( .C ( clk ), .D ( signal_9237 ), .Q ( signal_9238 ) ) ;
    buf_clk cell_3650 ( .C ( clk ), .D ( signal_9241 ), .Q ( signal_9242 ) ) ;
    buf_clk cell_3654 ( .C ( clk ), .D ( signal_9245 ), .Q ( signal_9246 ) ) ;
    buf_clk cell_3658 ( .C ( clk ), .D ( signal_9249 ), .Q ( signal_9250 ) ) ;
    buf_clk cell_3662 ( .C ( clk ), .D ( signal_9253 ), .Q ( signal_9254 ) ) ;
    buf_clk cell_3666 ( .C ( clk ), .D ( signal_9257 ), .Q ( signal_9258 ) ) ;
    buf_clk cell_3670 ( .C ( clk ), .D ( signal_9261 ), .Q ( signal_9262 ) ) ;
    buf_clk cell_3674 ( .C ( clk ), .D ( signal_9265 ), .Q ( signal_9266 ) ) ;
    buf_clk cell_3676 ( .C ( clk ), .D ( signal_9267 ), .Q ( signal_9268 ) ) ;
    buf_clk cell_3678 ( .C ( clk ), .D ( signal_9269 ), .Q ( signal_9270 ) ) ;
    buf_clk cell_3680 ( .C ( clk ), .D ( signal_9271 ), .Q ( signal_9272 ) ) ;
    buf_clk cell_3684 ( .C ( clk ), .D ( signal_9275 ), .Q ( signal_9276 ) ) ;
    buf_clk cell_3688 ( .C ( clk ), .D ( signal_9279 ), .Q ( signal_9280 ) ) ;
    buf_clk cell_3692 ( .C ( clk ), .D ( signal_9283 ), .Q ( signal_9284 ) ) ;
    buf_clk cell_3694 ( .C ( clk ), .D ( signal_9285 ), .Q ( signal_9286 ) ) ;
    buf_clk cell_3696 ( .C ( clk ), .D ( signal_9287 ), .Q ( signal_9288 ) ) ;
    buf_clk cell_3698 ( .C ( clk ), .D ( signal_9289 ), .Q ( signal_9290 ) ) ;
    buf_clk cell_3700 ( .C ( clk ), .D ( signal_9291 ), .Q ( signal_9292 ) ) ;
    buf_clk cell_3702 ( .C ( clk ), .D ( signal_9293 ), .Q ( signal_9294 ) ) ;
    buf_clk cell_3704 ( .C ( clk ), .D ( signal_9295 ), .Q ( signal_9296 ) ) ;
    buf_clk cell_3706 ( .C ( clk ), .D ( signal_9297 ), .Q ( signal_9298 ) ) ;
    buf_clk cell_3708 ( .C ( clk ), .D ( signal_9299 ), .Q ( signal_9300 ) ) ;
    buf_clk cell_3710 ( .C ( clk ), .D ( signal_9301 ), .Q ( signal_9302 ) ) ;
    buf_clk cell_3712 ( .C ( clk ), .D ( signal_9303 ), .Q ( signal_9304 ) ) ;
    buf_clk cell_3714 ( .C ( clk ), .D ( signal_9305 ), .Q ( signal_9306 ) ) ;
    buf_clk cell_3716 ( .C ( clk ), .D ( signal_9307 ), .Q ( signal_9308 ) ) ;
    buf_clk cell_3718 ( .C ( clk ), .D ( signal_9309 ), .Q ( signal_9310 ) ) ;
    buf_clk cell_3720 ( .C ( clk ), .D ( signal_9311 ), .Q ( signal_9312 ) ) ;
    buf_clk cell_3722 ( .C ( clk ), .D ( signal_9313 ), .Q ( signal_9314 ) ) ;
    buf_clk cell_3726 ( .C ( clk ), .D ( signal_9317 ), .Q ( signal_9318 ) ) ;
    buf_clk cell_3730 ( .C ( clk ), .D ( signal_9321 ), .Q ( signal_9322 ) ) ;
    buf_clk cell_3734 ( .C ( clk ), .D ( signal_9325 ), .Q ( signal_9326 ) ) ;
    buf_clk cell_3738 ( .C ( clk ), .D ( signal_9329 ), .Q ( signal_9330 ) ) ;
    buf_clk cell_3742 ( .C ( clk ), .D ( signal_9333 ), .Q ( signal_9334 ) ) ;
    buf_clk cell_3746 ( .C ( clk ), .D ( signal_9337 ), .Q ( signal_9338 ) ) ;
    buf_clk cell_3748 ( .C ( clk ), .D ( signal_9339 ), .Q ( signal_9340 ) ) ;
    buf_clk cell_3750 ( .C ( clk ), .D ( signal_9341 ), .Q ( signal_9342 ) ) ;
    buf_clk cell_3752 ( .C ( clk ), .D ( signal_9343 ), .Q ( signal_9344 ) ) ;
    buf_clk cell_3756 ( .C ( clk ), .D ( signal_9347 ), .Q ( signal_9348 ) ) ;
    buf_clk cell_3760 ( .C ( clk ), .D ( signal_9351 ), .Q ( signal_9352 ) ) ;
    buf_clk cell_3764 ( .C ( clk ), .D ( signal_9355 ), .Q ( signal_9356 ) ) ;
    buf_clk cell_3766 ( .C ( clk ), .D ( signal_9357 ), .Q ( signal_9358 ) ) ;
    buf_clk cell_3768 ( .C ( clk ), .D ( signal_9359 ), .Q ( signal_9360 ) ) ;
    buf_clk cell_3770 ( .C ( clk ), .D ( signal_9361 ), .Q ( signal_9362 ) ) ;
    buf_clk cell_3772 ( .C ( clk ), .D ( signal_9363 ), .Q ( signal_9364 ) ) ;
    buf_clk cell_3774 ( .C ( clk ), .D ( signal_9365 ), .Q ( signal_9366 ) ) ;
    buf_clk cell_3776 ( .C ( clk ), .D ( signal_9367 ), .Q ( signal_9368 ) ) ;
    buf_clk cell_3780 ( .C ( clk ), .D ( signal_9371 ), .Q ( signal_9372 ) ) ;
    buf_clk cell_3784 ( .C ( clk ), .D ( signal_9375 ), .Q ( signal_9376 ) ) ;
    buf_clk cell_3788 ( .C ( clk ), .D ( signal_9379 ), .Q ( signal_9380 ) ) ;
    buf_clk cell_3792 ( .C ( clk ), .D ( signal_9383 ), .Q ( signal_9384 ) ) ;
    buf_clk cell_3796 ( .C ( clk ), .D ( signal_9387 ), .Q ( signal_9388 ) ) ;
    buf_clk cell_3800 ( .C ( clk ), .D ( signal_9391 ), .Q ( signal_9392 ) ) ;
    buf_clk cell_3804 ( .C ( clk ), .D ( signal_9395 ), .Q ( signal_9396 ) ) ;
    buf_clk cell_3808 ( .C ( clk ), .D ( signal_9399 ), .Q ( signal_9400 ) ) ;
    buf_clk cell_3812 ( .C ( clk ), .D ( signal_9403 ), .Q ( signal_9404 ) ) ;
    buf_clk cell_3814 ( .C ( clk ), .D ( signal_9405 ), .Q ( signal_9406 ) ) ;
    buf_clk cell_3816 ( .C ( clk ), .D ( signal_9407 ), .Q ( signal_9408 ) ) ;
    buf_clk cell_3818 ( .C ( clk ), .D ( signal_9409 ), .Q ( signal_9410 ) ) ;
    buf_clk cell_3822 ( .C ( clk ), .D ( signal_9413 ), .Q ( signal_9414 ) ) ;
    buf_clk cell_3826 ( .C ( clk ), .D ( signal_9417 ), .Q ( signal_9418 ) ) ;
    buf_clk cell_3830 ( .C ( clk ), .D ( signal_9421 ), .Q ( signal_9422 ) ) ;
    buf_clk cell_3834 ( .C ( clk ), .D ( signal_9425 ), .Q ( signal_9426 ) ) ;
    buf_clk cell_3838 ( .C ( clk ), .D ( signal_9429 ), .Q ( signal_9430 ) ) ;
    buf_clk cell_3842 ( .C ( clk ), .D ( signal_9433 ), .Q ( signal_9434 ) ) ;
    buf_clk cell_3844 ( .C ( clk ), .D ( signal_9435 ), .Q ( signal_9436 ) ) ;
    buf_clk cell_3846 ( .C ( clk ), .D ( signal_9437 ), .Q ( signal_9438 ) ) ;
    buf_clk cell_3848 ( .C ( clk ), .D ( signal_9439 ), .Q ( signal_9440 ) ) ;
    buf_clk cell_3852 ( .C ( clk ), .D ( signal_9443 ), .Q ( signal_9444 ) ) ;
    buf_clk cell_3856 ( .C ( clk ), .D ( signal_9447 ), .Q ( signal_9448 ) ) ;
    buf_clk cell_3860 ( .C ( clk ), .D ( signal_9451 ), .Q ( signal_9452 ) ) ;
    buf_clk cell_3862 ( .C ( clk ), .D ( signal_9453 ), .Q ( signal_9454 ) ) ;
    buf_clk cell_3864 ( .C ( clk ), .D ( signal_9455 ), .Q ( signal_9456 ) ) ;
    buf_clk cell_3866 ( .C ( clk ), .D ( signal_9457 ), .Q ( signal_9458 ) ) ;
    buf_clk cell_3868 ( .C ( clk ), .D ( signal_9459 ), .Q ( signal_9460 ) ) ;
    buf_clk cell_3870 ( .C ( clk ), .D ( signal_9461 ), .Q ( signal_9462 ) ) ;
    buf_clk cell_3872 ( .C ( clk ), .D ( signal_9463 ), .Q ( signal_9464 ) ) ;
    buf_clk cell_3874 ( .C ( clk ), .D ( signal_9465 ), .Q ( signal_9466 ) ) ;
    buf_clk cell_3876 ( .C ( clk ), .D ( signal_9467 ), .Q ( signal_9468 ) ) ;
    buf_clk cell_3878 ( .C ( clk ), .D ( signal_9469 ), .Q ( signal_9470 ) ) ;
    buf_clk cell_3882 ( .C ( clk ), .D ( signal_9473 ), .Q ( signal_9474 ) ) ;
    buf_clk cell_3886 ( .C ( clk ), .D ( signal_9477 ), .Q ( signal_9478 ) ) ;
    buf_clk cell_3890 ( .C ( clk ), .D ( signal_9481 ), .Q ( signal_9482 ) ) ;
    buf_clk cell_3900 ( .C ( clk ), .D ( signal_9491 ), .Q ( signal_9492 ) ) ;
    buf_clk cell_3906 ( .C ( clk ), .D ( signal_9497 ), .Q ( signal_9498 ) ) ;
    buf_clk cell_3912 ( .C ( clk ), .D ( signal_9503 ), .Q ( signal_9504 ) ) ;
    buf_clk cell_3918 ( .C ( clk ), .D ( signal_9509 ), .Q ( signal_9510 ) ) ;
    buf_clk cell_3924 ( .C ( clk ), .D ( signal_9515 ), .Q ( signal_9516 ) ) ;
    buf_clk cell_3930 ( .C ( clk ), .D ( signal_9521 ), .Q ( signal_9522 ) ) ;
    buf_clk cell_3936 ( .C ( clk ), .D ( signal_9527 ), .Q ( signal_9528 ) ) ;
    buf_clk cell_3942 ( .C ( clk ), .D ( signal_9533 ), .Q ( signal_9534 ) ) ;
    buf_clk cell_3948 ( .C ( clk ), .D ( signal_9539 ), .Q ( signal_9540 ) ) ;
    buf_clk cell_3952 ( .C ( clk ), .D ( signal_9543 ), .Q ( signal_9544 ) ) ;
    buf_clk cell_3956 ( .C ( clk ), .D ( signal_9547 ), .Q ( signal_9548 ) ) ;
    buf_clk cell_3960 ( .C ( clk ), .D ( signal_9551 ), .Q ( signal_9552 ) ) ;
    buf_clk cell_3966 ( .C ( clk ), .D ( signal_9557 ), .Q ( signal_9558 ) ) ;
    buf_clk cell_3972 ( .C ( clk ), .D ( signal_9563 ), .Q ( signal_9564 ) ) ;
    buf_clk cell_3978 ( .C ( clk ), .D ( signal_9569 ), .Q ( signal_9570 ) ) ;
    buf_clk cell_3982 ( .C ( clk ), .D ( signal_9573 ), .Q ( signal_9574 ) ) ;
    buf_clk cell_3986 ( .C ( clk ), .D ( signal_9577 ), .Q ( signal_9578 ) ) ;
    buf_clk cell_3990 ( .C ( clk ), .D ( signal_9581 ), .Q ( signal_9582 ) ) ;
    buf_clk cell_3994 ( .C ( clk ), .D ( signal_9585 ), .Q ( signal_9586 ) ) ;
    buf_clk cell_3998 ( .C ( clk ), .D ( signal_9589 ), .Q ( signal_9590 ) ) ;
    buf_clk cell_4002 ( .C ( clk ), .D ( signal_9593 ), .Q ( signal_9594 ) ) ;
    buf_clk cell_4006 ( .C ( clk ), .D ( signal_9597 ), .Q ( signal_9598 ) ) ;
    buf_clk cell_4010 ( .C ( clk ), .D ( signal_9601 ), .Q ( signal_9602 ) ) ;
    buf_clk cell_4014 ( .C ( clk ), .D ( signal_9605 ), .Q ( signal_9606 ) ) ;
    buf_clk cell_4018 ( .C ( clk ), .D ( signal_9609 ), .Q ( signal_9610 ) ) ;
    buf_clk cell_4022 ( .C ( clk ), .D ( signal_9613 ), .Q ( signal_9614 ) ) ;
    buf_clk cell_4026 ( .C ( clk ), .D ( signal_9617 ), .Q ( signal_9618 ) ) ;
    buf_clk cell_4030 ( .C ( clk ), .D ( signal_9621 ), .Q ( signal_9622 ) ) ;
    buf_clk cell_4034 ( .C ( clk ), .D ( signal_9625 ), .Q ( signal_9626 ) ) ;
    buf_clk cell_4038 ( .C ( clk ), .D ( signal_9629 ), .Q ( signal_9630 ) ) ;
    buf_clk cell_4044 ( .C ( clk ), .D ( signal_9635 ), .Q ( signal_9636 ) ) ;
    buf_clk cell_4050 ( .C ( clk ), .D ( signal_9641 ), .Q ( signal_9642 ) ) ;
    buf_clk cell_4056 ( .C ( clk ), .D ( signal_9647 ), .Q ( signal_9648 ) ) ;
    buf_clk cell_4060 ( .C ( clk ), .D ( signal_9651 ), .Q ( signal_9652 ) ) ;
    buf_clk cell_4064 ( .C ( clk ), .D ( signal_9655 ), .Q ( signal_9656 ) ) ;
    buf_clk cell_4068 ( .C ( clk ), .D ( signal_9659 ), .Q ( signal_9660 ) ) ;
    buf_clk cell_4102 ( .C ( clk ), .D ( signal_9693 ), .Q ( signal_9694 ) ) ;
    buf_clk cell_4106 ( .C ( clk ), .D ( signal_9697 ), .Q ( signal_9698 ) ) ;
    buf_clk cell_4110 ( .C ( clk ), .D ( signal_9701 ), .Q ( signal_9702 ) ) ;
    buf_clk cell_4134 ( .C ( clk ), .D ( signal_9725 ), .Q ( signal_9726 ) ) ;
    buf_clk cell_4140 ( .C ( clk ), .D ( signal_9731 ), .Q ( signal_9732 ) ) ;
    buf_clk cell_4146 ( .C ( clk ), .D ( signal_9737 ), .Q ( signal_9738 ) ) ;
    buf_clk cell_4156 ( .C ( clk ), .D ( signal_9747 ), .Q ( signal_9748 ) ) ;
    buf_clk cell_4160 ( .C ( clk ), .D ( signal_9751 ), .Q ( signal_9752 ) ) ;
    buf_clk cell_4164 ( .C ( clk ), .D ( signal_9755 ), .Q ( signal_9756 ) ) ;
    buf_clk cell_4182 ( .C ( clk ), .D ( signal_9773 ), .Q ( signal_9774 ) ) ;
    buf_clk cell_4188 ( .C ( clk ), .D ( signal_9779 ), .Q ( signal_9780 ) ) ;
    buf_clk cell_4194 ( .C ( clk ), .D ( signal_9785 ), .Q ( signal_9786 ) ) ;
    buf_clk cell_4198 ( .C ( clk ), .D ( signal_9789 ), .Q ( signal_9790 ) ) ;
    buf_clk cell_4202 ( .C ( clk ), .D ( signal_9793 ), .Q ( signal_9794 ) ) ;
    buf_clk cell_4206 ( .C ( clk ), .D ( signal_9797 ), .Q ( signal_9798 ) ) ;
    buf_clk cell_4222 ( .C ( clk ), .D ( signal_9813 ), .Q ( signal_9814 ) ) ;
    buf_clk cell_4226 ( .C ( clk ), .D ( signal_9817 ), .Q ( signal_9818 ) ) ;
    buf_clk cell_4230 ( .C ( clk ), .D ( signal_9821 ), .Q ( signal_9822 ) ) ;
    buf_clk cell_4234 ( .C ( clk ), .D ( signal_9825 ), .Q ( signal_9826 ) ) ;
    buf_clk cell_4238 ( .C ( clk ), .D ( signal_9829 ), .Q ( signal_9830 ) ) ;
    buf_clk cell_4242 ( .C ( clk ), .D ( signal_9833 ), .Q ( signal_9834 ) ) ;
    buf_clk cell_4246 ( .C ( clk ), .D ( signal_9837 ), .Q ( signal_9838 ) ) ;
    buf_clk cell_4250 ( .C ( clk ), .D ( signal_9841 ), .Q ( signal_9842 ) ) ;
    buf_clk cell_4254 ( .C ( clk ), .D ( signal_9845 ), .Q ( signal_9846 ) ) ;
    buf_clk cell_4266 ( .C ( clk ), .D ( signal_9857 ), .Q ( signal_9858 ) ) ;
    buf_clk cell_4272 ( .C ( clk ), .D ( signal_9863 ), .Q ( signal_9864 ) ) ;
    buf_clk cell_4278 ( .C ( clk ), .D ( signal_9869 ), .Q ( signal_9870 ) ) ;
    buf_clk cell_4282 ( .C ( clk ), .D ( signal_9873 ), .Q ( signal_9874 ) ) ;
    buf_clk cell_4286 ( .C ( clk ), .D ( signal_9877 ), .Q ( signal_9878 ) ) ;
    buf_clk cell_4290 ( .C ( clk ), .D ( signal_9881 ), .Q ( signal_9882 ) ) ;
    buf_clk cell_4296 ( .C ( clk ), .D ( signal_9887 ), .Q ( signal_9888 ) ) ;
    buf_clk cell_4302 ( .C ( clk ), .D ( signal_9893 ), .Q ( signal_9894 ) ) ;
    buf_clk cell_4308 ( .C ( clk ), .D ( signal_9899 ), .Q ( signal_9900 ) ) ;
    buf_clk cell_4312 ( .C ( clk ), .D ( signal_9903 ), .Q ( signal_9904 ) ) ;
    buf_clk cell_4316 ( .C ( clk ), .D ( signal_9907 ), .Q ( signal_9908 ) ) ;
    buf_clk cell_4320 ( .C ( clk ), .D ( signal_9911 ), .Q ( signal_9912 ) ) ;
    buf_clk cell_4324 ( .C ( clk ), .D ( signal_9915 ), .Q ( signal_9916 ) ) ;
    buf_clk cell_4328 ( .C ( clk ), .D ( signal_9919 ), .Q ( signal_9920 ) ) ;
    buf_clk cell_4332 ( .C ( clk ), .D ( signal_9923 ), .Q ( signal_9924 ) ) ;
    buf_clk cell_4336 ( .C ( clk ), .D ( signal_9927 ), .Q ( signal_9928 ) ) ;
    buf_clk cell_4340 ( .C ( clk ), .D ( signal_9931 ), .Q ( signal_9932 ) ) ;
    buf_clk cell_4344 ( .C ( clk ), .D ( signal_9935 ), .Q ( signal_9936 ) ) ;
    buf_clk cell_4354 ( .C ( clk ), .D ( signal_9945 ), .Q ( signal_9946 ) ) ;
    buf_clk cell_4358 ( .C ( clk ), .D ( signal_9949 ), .Q ( signal_9950 ) ) ;
    buf_clk cell_4362 ( .C ( clk ), .D ( signal_9953 ), .Q ( signal_9954 ) ) ;
    buf_clk cell_4366 ( .C ( clk ), .D ( signal_9957 ), .Q ( signal_9958 ) ) ;
    buf_clk cell_4370 ( .C ( clk ), .D ( signal_9961 ), .Q ( signal_9962 ) ) ;
    buf_clk cell_4374 ( .C ( clk ), .D ( signal_9965 ), .Q ( signal_9966 ) ) ;
    buf_clk cell_4380 ( .C ( clk ), .D ( signal_9971 ), .Q ( signal_9972 ) ) ;
    buf_clk cell_4386 ( .C ( clk ), .D ( signal_9977 ), .Q ( signal_9978 ) ) ;
    buf_clk cell_4392 ( .C ( clk ), .D ( signal_9983 ), .Q ( signal_9984 ) ) ;
    buf_clk cell_4408 ( .C ( clk ), .D ( signal_9999 ), .Q ( signal_10000 ) ) ;
    buf_clk cell_4412 ( .C ( clk ), .D ( signal_10003 ), .Q ( signal_10004 ) ) ;
    buf_clk cell_4416 ( .C ( clk ), .D ( signal_10007 ), .Q ( signal_10008 ) ) ;
    buf_clk cell_4422 ( .C ( clk ), .D ( signal_10013 ), .Q ( signal_10014 ) ) ;
    buf_clk cell_4428 ( .C ( clk ), .D ( signal_10019 ), .Q ( signal_10020 ) ) ;
    buf_clk cell_4434 ( .C ( clk ), .D ( signal_10025 ), .Q ( signal_10026 ) ) ;
    buf_clk cell_4440 ( .C ( clk ), .D ( signal_10031 ), .Q ( signal_10032 ) ) ;
    buf_clk cell_4446 ( .C ( clk ), .D ( signal_10037 ), .Q ( signal_10038 ) ) ;
    buf_clk cell_4452 ( .C ( clk ), .D ( signal_10043 ), .Q ( signal_10044 ) ) ;
    buf_clk cell_4458 ( .C ( clk ), .D ( signal_10049 ), .Q ( signal_10050 ) ) ;
    buf_clk cell_4464 ( .C ( clk ), .D ( signal_10055 ), .Q ( signal_10056 ) ) ;
    buf_clk cell_4470 ( .C ( clk ), .D ( signal_10061 ), .Q ( signal_10062 ) ) ;
    buf_clk cell_4474 ( .C ( clk ), .D ( signal_10065 ), .Q ( signal_10066 ) ) ;
    buf_clk cell_4478 ( .C ( clk ), .D ( signal_10069 ), .Q ( signal_10070 ) ) ;
    buf_clk cell_4482 ( .C ( clk ), .D ( signal_10073 ), .Q ( signal_10074 ) ) ;
    buf_clk cell_4500 ( .C ( clk ), .D ( signal_10091 ), .Q ( signal_10092 ) ) ;
    buf_clk cell_4508 ( .C ( clk ), .D ( signal_10099 ), .Q ( signal_10100 ) ) ;
    buf_clk cell_4516 ( .C ( clk ), .D ( signal_10107 ), .Q ( signal_10108 ) ) ;
    buf_clk cell_4534 ( .C ( clk ), .D ( signal_10125 ), .Q ( signal_10126 ) ) ;
    buf_clk cell_4540 ( .C ( clk ), .D ( signal_10131 ), .Q ( signal_10132 ) ) ;
    buf_clk cell_4546 ( .C ( clk ), .D ( signal_10137 ), .Q ( signal_10138 ) ) ;
    buf_clk cell_4552 ( .C ( clk ), .D ( signal_10143 ), .Q ( signal_10144 ) ) ;
    buf_clk cell_4558 ( .C ( clk ), .D ( signal_10149 ), .Q ( signal_10150 ) ) ;
    buf_clk cell_4564 ( .C ( clk ), .D ( signal_10155 ), .Q ( signal_10156 ) ) ;
    buf_clk cell_4582 ( .C ( clk ), .D ( signal_10173 ), .Q ( signal_10174 ) ) ;
    buf_clk cell_4588 ( .C ( clk ), .D ( signal_10179 ), .Q ( signal_10180 ) ) ;
    buf_clk cell_4594 ( .C ( clk ), .D ( signal_10185 ), .Q ( signal_10186 ) ) ;
    buf_clk cell_4636 ( .C ( clk ), .D ( signal_10227 ), .Q ( signal_10228 ) ) ;
    buf_clk cell_4642 ( .C ( clk ), .D ( signal_10233 ), .Q ( signal_10234 ) ) ;
    buf_clk cell_4648 ( .C ( clk ), .D ( signal_10239 ), .Q ( signal_10240 ) ) ;
    buf_clk cell_4654 ( .C ( clk ), .D ( signal_10245 ), .Q ( signal_10246 ) ) ;
    buf_clk cell_4660 ( .C ( clk ), .D ( signal_10251 ), .Q ( signal_10252 ) ) ;
    buf_clk cell_4666 ( .C ( clk ), .D ( signal_10257 ), .Q ( signal_10258 ) ) ;
    buf_clk cell_4672 ( .C ( clk ), .D ( signal_10263 ), .Q ( signal_10264 ) ) ;
    buf_clk cell_4678 ( .C ( clk ), .D ( signal_10269 ), .Q ( signal_10270 ) ) ;
    buf_clk cell_4684 ( .C ( clk ), .D ( signal_10275 ), .Q ( signal_10276 ) ) ;
    buf_clk cell_4708 ( .C ( clk ), .D ( signal_10299 ), .Q ( signal_10300 ) ) ;
    buf_clk cell_4714 ( .C ( clk ), .D ( signal_10305 ), .Q ( signal_10306 ) ) ;
    buf_clk cell_4720 ( .C ( clk ), .D ( signal_10311 ), .Q ( signal_10312 ) ) ;
    buf_clk cell_4732 ( .C ( clk ), .D ( signal_10323 ), .Q ( signal_10324 ) ) ;
    buf_clk cell_4738 ( .C ( clk ), .D ( signal_10329 ), .Q ( signal_10330 ) ) ;
    buf_clk cell_4744 ( .C ( clk ), .D ( signal_10335 ), .Q ( signal_10336 ) ) ;
    buf_clk cell_4758 ( .C ( clk ), .D ( signal_10349 ), .Q ( signal_10350 ) ) ;
    buf_clk cell_4766 ( .C ( clk ), .D ( signal_10357 ), .Q ( signal_10358 ) ) ;
    buf_clk cell_4774 ( .C ( clk ), .D ( signal_10365 ), .Q ( signal_10366 ) ) ;
    buf_clk cell_4804 ( .C ( clk ), .D ( signal_10395 ), .Q ( signal_10396 ) ) ;
    buf_clk cell_4810 ( .C ( clk ), .D ( signal_10401 ), .Q ( signal_10402 ) ) ;
    buf_clk cell_4816 ( .C ( clk ), .D ( signal_10407 ), .Q ( signal_10408 ) ) ;
    buf_clk cell_4822 ( .C ( clk ), .D ( signal_10413 ), .Q ( signal_10414 ) ) ;
    buf_clk cell_4828 ( .C ( clk ), .D ( signal_10419 ), .Q ( signal_10420 ) ) ;
    buf_clk cell_4834 ( .C ( clk ), .D ( signal_10425 ), .Q ( signal_10426 ) ) ;
    buf_clk cell_4854 ( .C ( clk ), .D ( signal_10445 ), .Q ( signal_10446 ) ) ;
    buf_clk cell_4862 ( .C ( clk ), .D ( signal_10453 ), .Q ( signal_10454 ) ) ;
    buf_clk cell_4870 ( .C ( clk ), .D ( signal_10461 ), .Q ( signal_10462 ) ) ;
    buf_clk cell_4876 ( .C ( clk ), .D ( signal_10467 ), .Q ( signal_10468 ) ) ;
    buf_clk cell_4882 ( .C ( clk ), .D ( signal_10473 ), .Q ( signal_10474 ) ) ;
    buf_clk cell_4888 ( .C ( clk ), .D ( signal_10479 ), .Q ( signal_10480 ) ) ;
    buf_clk cell_4894 ( .C ( clk ), .D ( signal_10485 ), .Q ( signal_10486 ) ) ;
    buf_clk cell_4900 ( .C ( clk ), .D ( signal_10491 ), .Q ( signal_10492 ) ) ;
    buf_clk cell_4906 ( .C ( clk ), .D ( signal_10497 ), .Q ( signal_10498 ) ) ;
    buf_clk cell_4924 ( .C ( clk ), .D ( signal_10515 ), .Q ( signal_10516 ) ) ;
    buf_clk cell_4930 ( .C ( clk ), .D ( signal_10521 ), .Q ( signal_10522 ) ) ;
    buf_clk cell_4936 ( .C ( clk ), .D ( signal_10527 ), .Q ( signal_10528 ) ) ;
    buf_clk cell_4954 ( .C ( clk ), .D ( signal_10545 ), .Q ( signal_10546 ) ) ;
    buf_clk cell_4960 ( .C ( clk ), .D ( signal_10551 ), .Q ( signal_10552 ) ) ;
    buf_clk cell_4966 ( .C ( clk ), .D ( signal_10557 ), .Q ( signal_10558 ) ) ;
    buf_clk cell_4972 ( .C ( clk ), .D ( signal_10563 ), .Q ( signal_10564 ) ) ;
    buf_clk cell_4978 ( .C ( clk ), .D ( signal_10569 ), .Q ( signal_10570 ) ) ;
    buf_clk cell_4984 ( .C ( clk ), .D ( signal_10575 ), .Q ( signal_10576 ) ) ;
    buf_clk cell_5004 ( .C ( clk ), .D ( signal_10595 ), .Q ( signal_10596 ) ) ;
    buf_clk cell_5014 ( .C ( clk ), .D ( signal_10605 ), .Q ( signal_10606 ) ) ;
    buf_clk cell_5024 ( .C ( clk ), .D ( signal_10615 ), .Q ( signal_10616 ) ) ;
    buf_clk cell_5050 ( .C ( clk ), .D ( signal_10641 ), .Q ( signal_10642 ) ) ;
    buf_clk cell_5058 ( .C ( clk ), .D ( signal_10649 ), .Q ( signal_10650 ) ) ;
    buf_clk cell_5066 ( .C ( clk ), .D ( signal_10657 ), .Q ( signal_10658 ) ) ;
    buf_clk cell_5074 ( .C ( clk ), .D ( signal_10665 ), .Q ( signal_10666 ) ) ;
    buf_clk cell_5082 ( .C ( clk ), .D ( signal_10673 ), .Q ( signal_10674 ) ) ;
    buf_clk cell_5090 ( .C ( clk ), .D ( signal_10681 ), .Q ( signal_10682 ) ) ;
    buf_clk cell_5148 ( .C ( clk ), .D ( signal_10739 ), .Q ( signal_10740 ) ) ;
    buf_clk cell_5158 ( .C ( clk ), .D ( signal_10749 ), .Q ( signal_10750 ) ) ;
    buf_clk cell_5168 ( .C ( clk ), .D ( signal_10759 ), .Q ( signal_10760 ) ) ;
    buf_clk cell_5200 ( .C ( clk ), .D ( signal_10791 ), .Q ( signal_10792 ) ) ;
    buf_clk cell_5208 ( .C ( clk ), .D ( signal_10799 ), .Q ( signal_10800 ) ) ;
    buf_clk cell_5216 ( .C ( clk ), .D ( signal_10807 ), .Q ( signal_10808 ) ) ;
    buf_clk cell_5242 ( .C ( clk ), .D ( signal_10833 ), .Q ( signal_10834 ) ) ;
    buf_clk cell_5250 ( .C ( clk ), .D ( signal_10841 ), .Q ( signal_10842 ) ) ;
    buf_clk cell_5258 ( .C ( clk ), .D ( signal_10849 ), .Q ( signal_10850 ) ) ;
    buf_clk cell_5266 ( .C ( clk ), .D ( signal_10857 ), .Q ( signal_10858 ) ) ;
    buf_clk cell_5274 ( .C ( clk ), .D ( signal_10865 ), .Q ( signal_10866 ) ) ;
    buf_clk cell_5282 ( .C ( clk ), .D ( signal_10873 ), .Q ( signal_10874 ) ) ;
    buf_clk cell_5290 ( .C ( clk ), .D ( signal_10881 ), .Q ( signal_10882 ) ) ;
    buf_clk cell_5298 ( .C ( clk ), .D ( signal_10889 ), .Q ( signal_10890 ) ) ;
    buf_clk cell_5306 ( .C ( clk ), .D ( signal_10897 ), .Q ( signal_10898 ) ) ;
    buf_clk cell_5316 ( .C ( clk ), .D ( signal_10907 ), .Q ( signal_10908 ) ) ;
    buf_clk cell_5326 ( .C ( clk ), .D ( signal_10917 ), .Q ( signal_10918 ) ) ;
    buf_clk cell_5336 ( .C ( clk ), .D ( signal_10927 ), .Q ( signal_10928 ) ) ;
    buf_clk cell_5344 ( .C ( clk ), .D ( signal_10935 ), .Q ( signal_10936 ) ) ;
    buf_clk cell_5352 ( .C ( clk ), .D ( signal_10943 ), .Q ( signal_10944 ) ) ;
    buf_clk cell_5360 ( .C ( clk ), .D ( signal_10951 ), .Q ( signal_10952 ) ) ;
    buf_clk cell_5368 ( .C ( clk ), .D ( signal_10959 ), .Q ( signal_10960 ) ) ;
    buf_clk cell_5376 ( .C ( clk ), .D ( signal_10967 ), .Q ( signal_10968 ) ) ;
    buf_clk cell_5384 ( .C ( clk ), .D ( signal_10975 ), .Q ( signal_10976 ) ) ;
    buf_clk cell_5398 ( .C ( clk ), .D ( signal_10989 ), .Q ( signal_10990 ) ) ;
    buf_clk cell_5406 ( .C ( clk ), .D ( signal_10997 ), .Q ( signal_10998 ) ) ;
    buf_clk cell_5414 ( .C ( clk ), .D ( signal_11005 ), .Q ( signal_11006 ) ) ;
    buf_clk cell_5422 ( .C ( clk ), .D ( signal_11013 ), .Q ( signal_11014 ) ) ;
    buf_clk cell_5430 ( .C ( clk ), .D ( signal_11021 ), .Q ( signal_11022 ) ) ;
    buf_clk cell_5438 ( .C ( clk ), .D ( signal_11029 ), .Q ( signal_11030 ) ) ;
    buf_clk cell_5446 ( .C ( clk ), .D ( signal_11037 ), .Q ( signal_11038 ) ) ;
    buf_clk cell_5454 ( .C ( clk ), .D ( signal_11045 ), .Q ( signal_11046 ) ) ;
    buf_clk cell_5462 ( .C ( clk ), .D ( signal_11053 ), .Q ( signal_11054 ) ) ;
    buf_clk cell_5572 ( .C ( clk ), .D ( signal_11163 ), .Q ( signal_11164 ) ) ;
    buf_clk cell_5582 ( .C ( clk ), .D ( signal_11173 ), .Q ( signal_11174 ) ) ;
    buf_clk cell_5592 ( .C ( clk ), .D ( signal_11183 ), .Q ( signal_11184 ) ) ;
    buf_clk cell_5650 ( .C ( clk ), .D ( signal_11241 ), .Q ( signal_11242 ) ) ;
    buf_clk cell_5660 ( .C ( clk ), .D ( signal_11251 ), .Q ( signal_11252 ) ) ;
    buf_clk cell_5670 ( .C ( clk ), .D ( signal_11261 ), .Q ( signal_11262 ) ) ;
    buf_clk cell_6256 ( .C ( clk ), .D ( signal_11847 ), .Q ( signal_11848 ) ) ;
    buf_clk cell_6270 ( .C ( clk ), .D ( signal_11861 ), .Q ( signal_11862 ) ) ;
    buf_clk cell_6284 ( .C ( clk ), .D ( signal_11875 ), .Q ( signal_11876 ) ) ;
    buf_clk cell_6322 ( .C ( clk ), .D ( signal_11913 ), .Q ( signal_11914 ) ) ;
    buf_clk cell_6336 ( .C ( clk ), .D ( signal_11927 ), .Q ( signal_11928 ) ) ;
    buf_clk cell_6350 ( .C ( clk ), .D ( signal_11941 ), .Q ( signal_11942 ) ) ;
    buf_clk cell_6442 ( .C ( clk ), .D ( signal_12033 ), .Q ( signal_12034 ) ) ;
    buf_clk cell_6458 ( .C ( clk ), .D ( signal_12049 ), .Q ( signal_12050 ) ) ;
    buf_clk cell_6474 ( .C ( clk ), .D ( signal_12065 ), .Q ( signal_12066 ) ) ;
    buf_clk cell_6502 ( .C ( clk ), .D ( signal_12093 ), .Q ( signal_12094 ) ) ;
    buf_clk cell_6518 ( .C ( clk ), .D ( signal_12109 ), .Q ( signal_12110 ) ) ;
    buf_clk cell_6534 ( .C ( clk ), .D ( signal_12125 ), .Q ( signal_12126 ) ) ;
    buf_clk cell_6736 ( .C ( clk ), .D ( signal_12327 ), .Q ( signal_12328 ) ) ;
    buf_clk cell_6754 ( .C ( clk ), .D ( signal_12345 ), .Q ( signal_12346 ) ) ;
    buf_clk cell_6772 ( .C ( clk ), .D ( signal_12363 ), .Q ( signal_12364 ) ) ;
    buf_clk cell_6886 ( .C ( clk ), .D ( signal_12477 ), .Q ( signal_12478 ) ) ;
    buf_clk cell_6906 ( .C ( clk ), .D ( signal_12497 ), .Q ( signal_12498 ) ) ;
    buf_clk cell_6926 ( .C ( clk ), .D ( signal_12517 ), .Q ( signal_12518 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_3891 ( .C ( clk ), .D ( signal_9358 ), .Q ( signal_9483 ) ) ;
    buf_clk cell_3893 ( .C ( clk ), .D ( signal_9360 ), .Q ( signal_9485 ) ) ;
    buf_clk cell_3895 ( .C ( clk ), .D ( signal_9362 ), .Q ( signal_9487 ) ) ;
    buf_clk cell_3901 ( .C ( clk ), .D ( signal_9492 ), .Q ( signal_9493 ) ) ;
    buf_clk cell_3907 ( .C ( clk ), .D ( signal_9498 ), .Q ( signal_9499 ) ) ;
    buf_clk cell_3913 ( .C ( clk ), .D ( signal_9504 ), .Q ( signal_9505 ) ) ;
    buf_clk cell_3919 ( .C ( clk ), .D ( signal_9510 ), .Q ( signal_9511 ) ) ;
    buf_clk cell_3925 ( .C ( clk ), .D ( signal_9516 ), .Q ( signal_9517 ) ) ;
    buf_clk cell_3931 ( .C ( clk ), .D ( signal_9522 ), .Q ( signal_9523 ) ) ;
    buf_clk cell_3937 ( .C ( clk ), .D ( signal_9528 ), .Q ( signal_9529 ) ) ;
    buf_clk cell_3943 ( .C ( clk ), .D ( signal_9534 ), .Q ( signal_9535 ) ) ;
    buf_clk cell_3949 ( .C ( clk ), .D ( signal_9540 ), .Q ( signal_9541 ) ) ;
    buf_clk cell_3953 ( .C ( clk ), .D ( signal_9544 ), .Q ( signal_9545 ) ) ;
    buf_clk cell_3957 ( .C ( clk ), .D ( signal_9548 ), .Q ( signal_9549 ) ) ;
    buf_clk cell_3961 ( .C ( clk ), .D ( signal_9552 ), .Q ( signal_9553 ) ) ;
    buf_clk cell_3967 ( .C ( clk ), .D ( signal_9558 ), .Q ( signal_9559 ) ) ;
    buf_clk cell_3973 ( .C ( clk ), .D ( signal_9564 ), .Q ( signal_9565 ) ) ;
    buf_clk cell_3979 ( .C ( clk ), .D ( signal_9570 ), .Q ( signal_9571 ) ) ;
    buf_clk cell_3983 ( .C ( clk ), .D ( signal_9574 ), .Q ( signal_9575 ) ) ;
    buf_clk cell_3987 ( .C ( clk ), .D ( signal_9578 ), .Q ( signal_9579 ) ) ;
    buf_clk cell_3991 ( .C ( clk ), .D ( signal_9582 ), .Q ( signal_9583 ) ) ;
    buf_clk cell_3995 ( .C ( clk ), .D ( signal_9586 ), .Q ( signal_9587 ) ) ;
    buf_clk cell_3999 ( .C ( clk ), .D ( signal_9590 ), .Q ( signal_9591 ) ) ;
    buf_clk cell_4003 ( .C ( clk ), .D ( signal_9594 ), .Q ( signal_9595 ) ) ;
    buf_clk cell_4007 ( .C ( clk ), .D ( signal_9598 ), .Q ( signal_9599 ) ) ;
    buf_clk cell_4011 ( .C ( clk ), .D ( signal_9602 ), .Q ( signal_9603 ) ) ;
    buf_clk cell_4015 ( .C ( clk ), .D ( signal_9606 ), .Q ( signal_9607 ) ) ;
    buf_clk cell_4019 ( .C ( clk ), .D ( signal_9610 ), .Q ( signal_9611 ) ) ;
    buf_clk cell_4023 ( .C ( clk ), .D ( signal_9614 ), .Q ( signal_9615 ) ) ;
    buf_clk cell_4027 ( .C ( clk ), .D ( signal_9618 ), .Q ( signal_9619 ) ) ;
    buf_clk cell_4031 ( .C ( clk ), .D ( signal_9622 ), .Q ( signal_9623 ) ) ;
    buf_clk cell_4035 ( .C ( clk ), .D ( signal_9626 ), .Q ( signal_9627 ) ) ;
    buf_clk cell_4039 ( .C ( clk ), .D ( signal_9630 ), .Q ( signal_9631 ) ) ;
    buf_clk cell_4045 ( .C ( clk ), .D ( signal_9636 ), .Q ( signal_9637 ) ) ;
    buf_clk cell_4051 ( .C ( clk ), .D ( signal_9642 ), .Q ( signal_9643 ) ) ;
    buf_clk cell_4057 ( .C ( clk ), .D ( signal_9648 ), .Q ( signal_9649 ) ) ;
    buf_clk cell_4061 ( .C ( clk ), .D ( signal_9652 ), .Q ( signal_9653 ) ) ;
    buf_clk cell_4065 ( .C ( clk ), .D ( signal_9656 ), .Q ( signal_9657 ) ) ;
    buf_clk cell_4069 ( .C ( clk ), .D ( signal_9660 ), .Q ( signal_9661 ) ) ;
    buf_clk cell_4071 ( .C ( clk ), .D ( signal_1999 ), .Q ( signal_9663 ) ) ;
    buf_clk cell_4073 ( .C ( clk ), .D ( signal_4522 ), .Q ( signal_9665 ) ) ;
    buf_clk cell_4075 ( .C ( clk ), .D ( signal_4523 ), .Q ( signal_9667 ) ) ;
    buf_clk cell_4077 ( .C ( clk ), .D ( signal_9220 ), .Q ( signal_9669 ) ) ;
    buf_clk cell_4079 ( .C ( clk ), .D ( signal_9222 ), .Q ( signal_9671 ) ) ;
    buf_clk cell_4081 ( .C ( clk ), .D ( signal_9224 ), .Q ( signal_9673 ) ) ;
    buf_clk cell_4083 ( .C ( clk ), .D ( signal_1811 ), .Q ( signal_9675 ) ) ;
    buf_clk cell_4085 ( .C ( clk ), .D ( signal_4146 ), .Q ( signal_9677 ) ) ;
    buf_clk cell_4087 ( .C ( clk ), .D ( signal_4147 ), .Q ( signal_9679 ) ) ;
    buf_clk cell_4089 ( .C ( clk ), .D ( signal_1980 ), .Q ( signal_9681 ) ) ;
    buf_clk cell_4091 ( .C ( clk ), .D ( signal_4484 ), .Q ( signal_9683 ) ) ;
    buf_clk cell_4093 ( .C ( clk ), .D ( signal_4485 ), .Q ( signal_9685 ) ) ;
    buf_clk cell_4095 ( .C ( clk ), .D ( signal_1983 ), .Q ( signal_9687 ) ) ;
    buf_clk cell_4097 ( .C ( clk ), .D ( signal_4490 ), .Q ( signal_9689 ) ) ;
    buf_clk cell_4099 ( .C ( clk ), .D ( signal_4491 ), .Q ( signal_9691 ) ) ;
    buf_clk cell_4103 ( .C ( clk ), .D ( signal_9694 ), .Q ( signal_9695 ) ) ;
    buf_clk cell_4107 ( .C ( clk ), .D ( signal_9698 ), .Q ( signal_9699 ) ) ;
    buf_clk cell_4111 ( .C ( clk ), .D ( signal_9702 ), .Q ( signal_9703 ) ) ;
    buf_clk cell_4113 ( .C ( clk ), .D ( signal_1965 ), .Q ( signal_9705 ) ) ;
    buf_clk cell_4115 ( .C ( clk ), .D ( signal_4454 ), .Q ( signal_9707 ) ) ;
    buf_clk cell_4117 ( .C ( clk ), .D ( signal_4455 ), .Q ( signal_9709 ) ) ;
    buf_clk cell_4119 ( .C ( clk ), .D ( signal_1968 ), .Q ( signal_9711 ) ) ;
    buf_clk cell_4121 ( .C ( clk ), .D ( signal_4460 ), .Q ( signal_9713 ) ) ;
    buf_clk cell_4123 ( .C ( clk ), .D ( signal_4461 ), .Q ( signal_9715 ) ) ;
    buf_clk cell_4125 ( .C ( clk ), .D ( signal_9286 ), .Q ( signal_9717 ) ) ;
    buf_clk cell_4127 ( .C ( clk ), .D ( signal_9288 ), .Q ( signal_9719 ) ) ;
    buf_clk cell_4129 ( .C ( clk ), .D ( signal_9290 ), .Q ( signal_9721 ) ) ;
    buf_clk cell_4135 ( .C ( clk ), .D ( signal_9726 ), .Q ( signal_9727 ) ) ;
    buf_clk cell_4141 ( .C ( clk ), .D ( signal_9732 ), .Q ( signal_9733 ) ) ;
    buf_clk cell_4147 ( .C ( clk ), .D ( signal_9738 ), .Q ( signal_9739 ) ) ;
    buf_clk cell_4149 ( .C ( clk ), .D ( signal_1970 ), .Q ( signal_9741 ) ) ;
    buf_clk cell_4151 ( .C ( clk ), .D ( signal_4464 ), .Q ( signal_9743 ) ) ;
    buf_clk cell_4153 ( .C ( clk ), .D ( signal_4465 ), .Q ( signal_9745 ) ) ;
    buf_clk cell_4157 ( .C ( clk ), .D ( signal_9748 ), .Q ( signal_9749 ) ) ;
    buf_clk cell_4161 ( .C ( clk ), .D ( signal_9752 ), .Q ( signal_9753 ) ) ;
    buf_clk cell_4165 ( .C ( clk ), .D ( signal_9756 ), .Q ( signal_9757 ) ) ;
    buf_clk cell_4167 ( .C ( clk ), .D ( signal_9180 ), .Q ( signal_9759 ) ) ;
    buf_clk cell_4169 ( .C ( clk ), .D ( signal_9184 ), .Q ( signal_9761 ) ) ;
    buf_clk cell_4171 ( .C ( clk ), .D ( signal_9188 ), .Q ( signal_9763 ) ) ;
    buf_clk cell_4173 ( .C ( clk ), .D ( signal_9298 ), .Q ( signal_9765 ) ) ;
    buf_clk cell_4175 ( .C ( clk ), .D ( signal_9300 ), .Q ( signal_9767 ) ) ;
    buf_clk cell_4177 ( .C ( clk ), .D ( signal_9302 ), .Q ( signal_9769 ) ) ;
    buf_clk cell_4183 ( .C ( clk ), .D ( signal_9774 ), .Q ( signal_9775 ) ) ;
    buf_clk cell_4189 ( .C ( clk ), .D ( signal_9780 ), .Q ( signal_9781 ) ) ;
    buf_clk cell_4195 ( .C ( clk ), .D ( signal_9786 ), .Q ( signal_9787 ) ) ;
    buf_clk cell_4199 ( .C ( clk ), .D ( signal_9790 ), .Q ( signal_9791 ) ) ;
    buf_clk cell_4203 ( .C ( clk ), .D ( signal_9794 ), .Q ( signal_9795 ) ) ;
    buf_clk cell_4207 ( .C ( clk ), .D ( signal_9798 ), .Q ( signal_9799 ) ) ;
    buf_clk cell_4209 ( .C ( clk ), .D ( signal_1755 ), .Q ( signal_9801 ) ) ;
    buf_clk cell_4211 ( .C ( clk ), .D ( signal_4034 ), .Q ( signal_9803 ) ) ;
    buf_clk cell_4213 ( .C ( clk ), .D ( signal_4035 ), .Q ( signal_9805 ) ) ;
    buf_clk cell_4215 ( .C ( clk ), .D ( signal_1987 ), .Q ( signal_9807 ) ) ;
    buf_clk cell_4217 ( .C ( clk ), .D ( signal_4498 ), .Q ( signal_9809 ) ) ;
    buf_clk cell_4219 ( .C ( clk ), .D ( signal_4499 ), .Q ( signal_9811 ) ) ;
    buf_clk cell_4223 ( .C ( clk ), .D ( signal_9814 ), .Q ( signal_9815 ) ) ;
    buf_clk cell_4227 ( .C ( clk ), .D ( signal_9818 ), .Q ( signal_9819 ) ) ;
    buf_clk cell_4231 ( .C ( clk ), .D ( signal_9822 ), .Q ( signal_9823 ) ) ;
    buf_clk cell_4235 ( .C ( clk ), .D ( signal_9826 ), .Q ( signal_9827 ) ) ;
    buf_clk cell_4239 ( .C ( clk ), .D ( signal_9830 ), .Q ( signal_9831 ) ) ;
    buf_clk cell_4243 ( .C ( clk ), .D ( signal_9834 ), .Q ( signal_9835 ) ) ;
    buf_clk cell_4247 ( .C ( clk ), .D ( signal_9838 ), .Q ( signal_9839 ) ) ;
    buf_clk cell_4251 ( .C ( clk ), .D ( signal_9842 ), .Q ( signal_9843 ) ) ;
    buf_clk cell_4255 ( .C ( clk ), .D ( signal_9846 ), .Q ( signal_9847 ) ) ;
    buf_clk cell_4257 ( .C ( clk ), .D ( signal_9258 ), .Q ( signal_9849 ) ) ;
    buf_clk cell_4259 ( .C ( clk ), .D ( signal_9262 ), .Q ( signal_9851 ) ) ;
    buf_clk cell_4261 ( .C ( clk ), .D ( signal_9266 ), .Q ( signal_9853 ) ) ;
    buf_clk cell_4267 ( .C ( clk ), .D ( signal_9858 ), .Q ( signal_9859 ) ) ;
    buf_clk cell_4273 ( .C ( clk ), .D ( signal_9864 ), .Q ( signal_9865 ) ) ;
    buf_clk cell_4279 ( .C ( clk ), .D ( signal_9870 ), .Q ( signal_9871 ) ) ;
    buf_clk cell_4283 ( .C ( clk ), .D ( signal_9874 ), .Q ( signal_9875 ) ) ;
    buf_clk cell_4287 ( .C ( clk ), .D ( signal_9878 ), .Q ( signal_9879 ) ) ;
    buf_clk cell_4291 ( .C ( clk ), .D ( signal_9882 ), .Q ( signal_9883 ) ) ;
    buf_clk cell_4297 ( .C ( clk ), .D ( signal_9888 ), .Q ( signal_9889 ) ) ;
    buf_clk cell_4303 ( .C ( clk ), .D ( signal_9894 ), .Q ( signal_9895 ) ) ;
    buf_clk cell_4309 ( .C ( clk ), .D ( signal_9900 ), .Q ( signal_9901 ) ) ;
    buf_clk cell_4313 ( .C ( clk ), .D ( signal_9904 ), .Q ( signal_9905 ) ) ;
    buf_clk cell_4317 ( .C ( clk ), .D ( signal_9908 ), .Q ( signal_9909 ) ) ;
    buf_clk cell_4321 ( .C ( clk ), .D ( signal_9912 ), .Q ( signal_9913 ) ) ;
    buf_clk cell_4325 ( .C ( clk ), .D ( signal_9916 ), .Q ( signal_9917 ) ) ;
    buf_clk cell_4329 ( .C ( clk ), .D ( signal_9920 ), .Q ( signal_9921 ) ) ;
    buf_clk cell_4333 ( .C ( clk ), .D ( signal_9924 ), .Q ( signal_9925 ) ) ;
    buf_clk cell_4337 ( .C ( clk ), .D ( signal_9928 ), .Q ( signal_9929 ) ) ;
    buf_clk cell_4341 ( .C ( clk ), .D ( signal_9932 ), .Q ( signal_9933 ) ) ;
    buf_clk cell_4345 ( .C ( clk ), .D ( signal_9936 ), .Q ( signal_9937 ) ) ;
    buf_clk cell_4347 ( .C ( clk ), .D ( signal_1966 ), .Q ( signal_9939 ) ) ;
    buf_clk cell_4349 ( .C ( clk ), .D ( signal_4456 ), .Q ( signal_9941 ) ) ;
    buf_clk cell_4351 ( .C ( clk ), .D ( signal_4457 ), .Q ( signal_9943 ) ) ;
    buf_clk cell_4355 ( .C ( clk ), .D ( signal_9946 ), .Q ( signal_9947 ) ) ;
    buf_clk cell_4359 ( .C ( clk ), .D ( signal_9950 ), .Q ( signal_9951 ) ) ;
    buf_clk cell_4363 ( .C ( clk ), .D ( signal_9954 ), .Q ( signal_9955 ) ) ;
    buf_clk cell_4367 ( .C ( clk ), .D ( signal_9958 ), .Q ( signal_9959 ) ) ;
    buf_clk cell_4371 ( .C ( clk ), .D ( signal_9962 ), .Q ( signal_9963 ) ) ;
    buf_clk cell_4375 ( .C ( clk ), .D ( signal_9966 ), .Q ( signal_9967 ) ) ;
    buf_clk cell_4381 ( .C ( clk ), .D ( signal_9972 ), .Q ( signal_9973 ) ) ;
    buf_clk cell_4387 ( .C ( clk ), .D ( signal_9978 ), .Q ( signal_9979 ) ) ;
    buf_clk cell_4393 ( .C ( clk ), .D ( signal_9984 ), .Q ( signal_9985 ) ) ;
    buf_clk cell_4395 ( .C ( clk ), .D ( signal_2011 ), .Q ( signal_9987 ) ) ;
    buf_clk cell_4397 ( .C ( clk ), .D ( signal_4546 ), .Q ( signal_9989 ) ) ;
    buf_clk cell_4399 ( .C ( clk ), .D ( signal_4547 ), .Q ( signal_9991 ) ) ;
    buf_clk cell_4401 ( .C ( clk ), .D ( signal_1843 ), .Q ( signal_9993 ) ) ;
    buf_clk cell_4403 ( .C ( clk ), .D ( signal_4210 ), .Q ( signal_9995 ) ) ;
    buf_clk cell_4405 ( .C ( clk ), .D ( signal_4211 ), .Q ( signal_9997 ) ) ;
    buf_clk cell_4409 ( .C ( clk ), .D ( signal_10000 ), .Q ( signal_10001 ) ) ;
    buf_clk cell_4413 ( .C ( clk ), .D ( signal_10004 ), .Q ( signal_10005 ) ) ;
    buf_clk cell_4417 ( .C ( clk ), .D ( signal_10008 ), .Q ( signal_10009 ) ) ;
    buf_clk cell_4423 ( .C ( clk ), .D ( signal_10014 ), .Q ( signal_10015 ) ) ;
    buf_clk cell_4429 ( .C ( clk ), .D ( signal_10020 ), .Q ( signal_10021 ) ) ;
    buf_clk cell_4435 ( .C ( clk ), .D ( signal_10026 ), .Q ( signal_10027 ) ) ;
    buf_clk cell_4441 ( .C ( clk ), .D ( signal_10032 ), .Q ( signal_10033 ) ) ;
    buf_clk cell_4447 ( .C ( clk ), .D ( signal_10038 ), .Q ( signal_10039 ) ) ;
    buf_clk cell_4453 ( .C ( clk ), .D ( signal_10044 ), .Q ( signal_10045 ) ) ;
    buf_clk cell_4459 ( .C ( clk ), .D ( signal_10050 ), .Q ( signal_10051 ) ) ;
    buf_clk cell_4465 ( .C ( clk ), .D ( signal_10056 ), .Q ( signal_10057 ) ) ;
    buf_clk cell_4471 ( .C ( clk ), .D ( signal_10062 ), .Q ( signal_10063 ) ) ;
    buf_clk cell_4475 ( .C ( clk ), .D ( signal_10066 ), .Q ( signal_10067 ) ) ;
    buf_clk cell_4479 ( .C ( clk ), .D ( signal_10070 ), .Q ( signal_10071 ) ) ;
    buf_clk cell_4483 ( .C ( clk ), .D ( signal_10074 ), .Q ( signal_10075 ) ) ;
    buf_clk cell_4485 ( .C ( clk ), .D ( signal_9246 ), .Q ( signal_10077 ) ) ;
    buf_clk cell_4487 ( .C ( clk ), .D ( signal_9250 ), .Q ( signal_10079 ) ) ;
    buf_clk cell_4489 ( .C ( clk ), .D ( signal_9254 ), .Q ( signal_10081 ) ) ;
    buf_clk cell_4491 ( .C ( clk ), .D ( signal_9276 ), .Q ( signal_10083 ) ) ;
    buf_clk cell_4493 ( .C ( clk ), .D ( signal_9280 ), .Q ( signal_10085 ) ) ;
    buf_clk cell_4495 ( .C ( clk ), .D ( signal_9284 ), .Q ( signal_10087 ) ) ;
    buf_clk cell_4501 ( .C ( clk ), .D ( signal_10092 ), .Q ( signal_10093 ) ) ;
    buf_clk cell_4509 ( .C ( clk ), .D ( signal_10100 ), .Q ( signal_10101 ) ) ;
    buf_clk cell_4517 ( .C ( clk ), .D ( signal_10108 ), .Q ( signal_10109 ) ) ;
    buf_clk cell_4521 ( .C ( clk ), .D ( signal_1758 ), .Q ( signal_10113 ) ) ;
    buf_clk cell_4525 ( .C ( clk ), .D ( signal_4040 ), .Q ( signal_10117 ) ) ;
    buf_clk cell_4529 ( .C ( clk ), .D ( signal_4041 ), .Q ( signal_10121 ) ) ;
    buf_clk cell_4535 ( .C ( clk ), .D ( signal_10126 ), .Q ( signal_10127 ) ) ;
    buf_clk cell_4541 ( .C ( clk ), .D ( signal_10132 ), .Q ( signal_10133 ) ) ;
    buf_clk cell_4547 ( .C ( clk ), .D ( signal_10138 ), .Q ( signal_10139 ) ) ;
    buf_clk cell_4553 ( .C ( clk ), .D ( signal_10144 ), .Q ( signal_10145 ) ) ;
    buf_clk cell_4559 ( .C ( clk ), .D ( signal_10150 ), .Q ( signal_10151 ) ) ;
    buf_clk cell_4565 ( .C ( clk ), .D ( signal_10156 ), .Q ( signal_10157 ) ) ;
    buf_clk cell_4569 ( .C ( clk ), .D ( signal_1762 ), .Q ( signal_10161 ) ) ;
    buf_clk cell_4573 ( .C ( clk ), .D ( signal_4048 ), .Q ( signal_10165 ) ) ;
    buf_clk cell_4577 ( .C ( clk ), .D ( signal_4049 ), .Q ( signal_10169 ) ) ;
    buf_clk cell_4583 ( .C ( clk ), .D ( signal_10174 ), .Q ( signal_10175 ) ) ;
    buf_clk cell_4589 ( .C ( clk ), .D ( signal_10180 ), .Q ( signal_10181 ) ) ;
    buf_clk cell_4595 ( .C ( clk ), .D ( signal_10186 ), .Q ( signal_10187 ) ) ;
    buf_clk cell_4599 ( .C ( clk ), .D ( signal_9156 ), .Q ( signal_10191 ) ) ;
    buf_clk cell_4603 ( .C ( clk ), .D ( signal_9160 ), .Q ( signal_10195 ) ) ;
    buf_clk cell_4607 ( .C ( clk ), .D ( signal_9164 ), .Q ( signal_10199 ) ) ;
    buf_clk cell_4611 ( .C ( clk ), .D ( signal_1845 ), .Q ( signal_10203 ) ) ;
    buf_clk cell_4615 ( .C ( clk ), .D ( signal_4214 ), .Q ( signal_10207 ) ) ;
    buf_clk cell_4619 ( .C ( clk ), .D ( signal_4215 ), .Q ( signal_10211 ) ) ;
    buf_clk cell_4637 ( .C ( clk ), .D ( signal_10228 ), .Q ( signal_10229 ) ) ;
    buf_clk cell_4643 ( .C ( clk ), .D ( signal_10234 ), .Q ( signal_10235 ) ) ;
    buf_clk cell_4649 ( .C ( clk ), .D ( signal_10240 ), .Q ( signal_10241 ) ) ;
    buf_clk cell_4655 ( .C ( clk ), .D ( signal_10246 ), .Q ( signal_10247 ) ) ;
    buf_clk cell_4661 ( .C ( clk ), .D ( signal_10252 ), .Q ( signal_10253 ) ) ;
    buf_clk cell_4667 ( .C ( clk ), .D ( signal_10258 ), .Q ( signal_10259 ) ) ;
    buf_clk cell_4673 ( .C ( clk ), .D ( signal_10264 ), .Q ( signal_10265 ) ) ;
    buf_clk cell_4679 ( .C ( clk ), .D ( signal_10270 ), .Q ( signal_10271 ) ) ;
    buf_clk cell_4685 ( .C ( clk ), .D ( signal_10276 ), .Q ( signal_10277 ) ) ;
    buf_clk cell_4695 ( .C ( clk ), .D ( signal_1810 ), .Q ( signal_10287 ) ) ;
    buf_clk cell_4699 ( .C ( clk ), .D ( signal_4144 ), .Q ( signal_10291 ) ) ;
    buf_clk cell_4703 ( .C ( clk ), .D ( signal_4145 ), .Q ( signal_10295 ) ) ;
    buf_clk cell_4709 ( .C ( clk ), .D ( signal_10300 ), .Q ( signal_10301 ) ) ;
    buf_clk cell_4715 ( .C ( clk ), .D ( signal_10306 ), .Q ( signal_10307 ) ) ;
    buf_clk cell_4721 ( .C ( clk ), .D ( signal_10312 ), .Q ( signal_10313 ) ) ;
    buf_clk cell_4733 ( .C ( clk ), .D ( signal_10324 ), .Q ( signal_10325 ) ) ;
    buf_clk cell_4739 ( .C ( clk ), .D ( signal_10330 ), .Q ( signal_10331 ) ) ;
    buf_clk cell_4745 ( .C ( clk ), .D ( signal_10336 ), .Q ( signal_10337 ) ) ;
    buf_clk cell_4759 ( .C ( clk ), .D ( signal_10350 ), .Q ( signal_10351 ) ) ;
    buf_clk cell_4767 ( .C ( clk ), .D ( signal_10358 ), .Q ( signal_10359 ) ) ;
    buf_clk cell_4775 ( .C ( clk ), .D ( signal_10366 ), .Q ( signal_10367 ) ) ;
    buf_clk cell_4779 ( .C ( clk ), .D ( signal_1814 ), .Q ( signal_10371 ) ) ;
    buf_clk cell_4783 ( .C ( clk ), .D ( signal_4152 ), .Q ( signal_10375 ) ) ;
    buf_clk cell_4787 ( .C ( clk ), .D ( signal_4153 ), .Q ( signal_10379 ) ) ;
    buf_clk cell_4791 ( .C ( clk ), .D ( signal_1820 ), .Q ( signal_10383 ) ) ;
    buf_clk cell_4795 ( .C ( clk ), .D ( signal_4164 ), .Q ( signal_10387 ) ) ;
    buf_clk cell_4799 ( .C ( clk ), .D ( signal_4165 ), .Q ( signal_10391 ) ) ;
    buf_clk cell_4805 ( .C ( clk ), .D ( signal_10396 ), .Q ( signal_10397 ) ) ;
    buf_clk cell_4811 ( .C ( clk ), .D ( signal_10402 ), .Q ( signal_10403 ) ) ;
    buf_clk cell_4817 ( .C ( clk ), .D ( signal_10408 ), .Q ( signal_10409 ) ) ;
    buf_clk cell_4823 ( .C ( clk ), .D ( signal_10414 ), .Q ( signal_10415 ) ) ;
    buf_clk cell_4829 ( .C ( clk ), .D ( signal_10420 ), .Q ( signal_10421 ) ) ;
    buf_clk cell_4835 ( .C ( clk ), .D ( signal_10426 ), .Q ( signal_10427 ) ) ;
    buf_clk cell_4839 ( .C ( clk ), .D ( signal_2006 ), .Q ( signal_10431 ) ) ;
    buf_clk cell_4843 ( .C ( clk ), .D ( signal_4536 ), .Q ( signal_10435 ) ) ;
    buf_clk cell_4847 ( .C ( clk ), .D ( signal_4537 ), .Q ( signal_10439 ) ) ;
    buf_clk cell_4855 ( .C ( clk ), .D ( signal_10446 ), .Q ( signal_10447 ) ) ;
    buf_clk cell_4863 ( .C ( clk ), .D ( signal_10454 ), .Q ( signal_10455 ) ) ;
    buf_clk cell_4871 ( .C ( clk ), .D ( signal_10462 ), .Q ( signal_10463 ) ) ;
    buf_clk cell_4877 ( .C ( clk ), .D ( signal_10468 ), .Q ( signal_10469 ) ) ;
    buf_clk cell_4883 ( .C ( clk ), .D ( signal_10474 ), .Q ( signal_10475 ) ) ;
    buf_clk cell_4889 ( .C ( clk ), .D ( signal_10480 ), .Q ( signal_10481 ) ) ;
    buf_clk cell_4895 ( .C ( clk ), .D ( signal_10486 ), .Q ( signal_10487 ) ) ;
    buf_clk cell_4901 ( .C ( clk ), .D ( signal_10492 ), .Q ( signal_10493 ) ) ;
    buf_clk cell_4907 ( .C ( clk ), .D ( signal_10498 ), .Q ( signal_10499 ) ) ;
    buf_clk cell_4925 ( .C ( clk ), .D ( signal_10516 ), .Q ( signal_10517 ) ) ;
    buf_clk cell_4931 ( .C ( clk ), .D ( signal_10522 ), .Q ( signal_10523 ) ) ;
    buf_clk cell_4937 ( .C ( clk ), .D ( signal_10528 ), .Q ( signal_10529 ) ) ;
    buf_clk cell_4955 ( .C ( clk ), .D ( signal_10546 ), .Q ( signal_10547 ) ) ;
    buf_clk cell_4961 ( .C ( clk ), .D ( signal_10552 ), .Q ( signal_10553 ) ) ;
    buf_clk cell_4967 ( .C ( clk ), .D ( signal_10558 ), .Q ( signal_10559 ) ) ;
    buf_clk cell_4973 ( .C ( clk ), .D ( signal_10564 ), .Q ( signal_10565 ) ) ;
    buf_clk cell_4979 ( .C ( clk ), .D ( signal_10570 ), .Q ( signal_10571 ) ) ;
    buf_clk cell_4985 ( .C ( clk ), .D ( signal_10576 ), .Q ( signal_10577 ) ) ;
    buf_clk cell_4989 ( .C ( clk ), .D ( signal_1818 ), .Q ( signal_10581 ) ) ;
    buf_clk cell_4993 ( .C ( clk ), .D ( signal_4160 ), .Q ( signal_10585 ) ) ;
    buf_clk cell_4997 ( .C ( clk ), .D ( signal_4161 ), .Q ( signal_10589 ) ) ;
    buf_clk cell_5005 ( .C ( clk ), .D ( signal_10596 ), .Q ( signal_10597 ) ) ;
    buf_clk cell_5015 ( .C ( clk ), .D ( signal_10606 ), .Q ( signal_10607 ) ) ;
    buf_clk cell_5025 ( .C ( clk ), .D ( signal_10616 ), .Q ( signal_10617 ) ) ;
    buf_clk cell_5031 ( .C ( clk ), .D ( signal_1988 ), .Q ( signal_10623 ) ) ;
    buf_clk cell_5037 ( .C ( clk ), .D ( signal_4500 ), .Q ( signal_10629 ) ) ;
    buf_clk cell_5043 ( .C ( clk ), .D ( signal_4501 ), .Q ( signal_10635 ) ) ;
    buf_clk cell_5051 ( .C ( clk ), .D ( signal_10642 ), .Q ( signal_10643 ) ) ;
    buf_clk cell_5059 ( .C ( clk ), .D ( signal_10650 ), .Q ( signal_10651 ) ) ;
    buf_clk cell_5067 ( .C ( clk ), .D ( signal_10658 ), .Q ( signal_10659 ) ) ;
    buf_clk cell_5075 ( .C ( clk ), .D ( signal_10666 ), .Q ( signal_10667 ) ) ;
    buf_clk cell_5083 ( .C ( clk ), .D ( signal_10674 ), .Q ( signal_10675 ) ) ;
    buf_clk cell_5091 ( .C ( clk ), .D ( signal_10682 ), .Q ( signal_10683 ) ) ;
    buf_clk cell_5149 ( .C ( clk ), .D ( signal_10740 ), .Q ( signal_10741 ) ) ;
    buf_clk cell_5159 ( .C ( clk ), .D ( signal_10750 ), .Q ( signal_10751 ) ) ;
    buf_clk cell_5169 ( .C ( clk ), .D ( signal_10760 ), .Q ( signal_10761 ) ) ;
    buf_clk cell_5175 ( .C ( clk ), .D ( signal_2016 ), .Q ( signal_10767 ) ) ;
    buf_clk cell_5181 ( .C ( clk ), .D ( signal_4556 ), .Q ( signal_10773 ) ) ;
    buf_clk cell_5187 ( .C ( clk ), .D ( signal_4557 ), .Q ( signal_10779 ) ) ;
    buf_clk cell_5201 ( .C ( clk ), .D ( signal_10792 ), .Q ( signal_10793 ) ) ;
    buf_clk cell_5209 ( .C ( clk ), .D ( signal_10800 ), .Q ( signal_10801 ) ) ;
    buf_clk cell_5217 ( .C ( clk ), .D ( signal_10808 ), .Q ( signal_10809 ) ) ;
    buf_clk cell_5223 ( .C ( clk ), .D ( signal_1979 ), .Q ( signal_10815 ) ) ;
    buf_clk cell_5229 ( .C ( clk ), .D ( signal_4482 ), .Q ( signal_10821 ) ) ;
    buf_clk cell_5235 ( .C ( clk ), .D ( signal_4483 ), .Q ( signal_10827 ) ) ;
    buf_clk cell_5243 ( .C ( clk ), .D ( signal_10834 ), .Q ( signal_10835 ) ) ;
    buf_clk cell_5251 ( .C ( clk ), .D ( signal_10842 ), .Q ( signal_10843 ) ) ;
    buf_clk cell_5259 ( .C ( clk ), .D ( signal_10850 ), .Q ( signal_10851 ) ) ;
    buf_clk cell_5267 ( .C ( clk ), .D ( signal_10858 ), .Q ( signal_10859 ) ) ;
    buf_clk cell_5275 ( .C ( clk ), .D ( signal_10866 ), .Q ( signal_10867 ) ) ;
    buf_clk cell_5283 ( .C ( clk ), .D ( signal_10874 ), .Q ( signal_10875 ) ) ;
    buf_clk cell_5291 ( .C ( clk ), .D ( signal_10882 ), .Q ( signal_10883 ) ) ;
    buf_clk cell_5299 ( .C ( clk ), .D ( signal_10890 ), .Q ( signal_10891 ) ) ;
    buf_clk cell_5307 ( .C ( clk ), .D ( signal_10898 ), .Q ( signal_10899 ) ) ;
    buf_clk cell_5317 ( .C ( clk ), .D ( signal_10908 ), .Q ( signal_10909 ) ) ;
    buf_clk cell_5327 ( .C ( clk ), .D ( signal_10918 ), .Q ( signal_10919 ) ) ;
    buf_clk cell_5337 ( .C ( clk ), .D ( signal_10928 ), .Q ( signal_10929 ) ) ;
    buf_clk cell_5345 ( .C ( clk ), .D ( signal_10936 ), .Q ( signal_10937 ) ) ;
    buf_clk cell_5353 ( .C ( clk ), .D ( signal_10944 ), .Q ( signal_10945 ) ) ;
    buf_clk cell_5361 ( .C ( clk ), .D ( signal_10952 ), .Q ( signal_10953 ) ) ;
    buf_clk cell_5369 ( .C ( clk ), .D ( signal_10960 ), .Q ( signal_10961 ) ) ;
    buf_clk cell_5377 ( .C ( clk ), .D ( signal_10968 ), .Q ( signal_10969 ) ) ;
    buf_clk cell_5385 ( .C ( clk ), .D ( signal_10976 ), .Q ( signal_10977 ) ) ;
    buf_clk cell_5399 ( .C ( clk ), .D ( signal_10990 ), .Q ( signal_10991 ) ) ;
    buf_clk cell_5407 ( .C ( clk ), .D ( signal_10998 ), .Q ( signal_10999 ) ) ;
    buf_clk cell_5415 ( .C ( clk ), .D ( signal_11006 ), .Q ( signal_11007 ) ) ;
    buf_clk cell_5423 ( .C ( clk ), .D ( signal_11014 ), .Q ( signal_11015 ) ) ;
    buf_clk cell_5431 ( .C ( clk ), .D ( signal_11022 ), .Q ( signal_11023 ) ) ;
    buf_clk cell_5439 ( .C ( clk ), .D ( signal_11030 ), .Q ( signal_11031 ) ) ;
    buf_clk cell_5447 ( .C ( clk ), .D ( signal_11038 ), .Q ( signal_11039 ) ) ;
    buf_clk cell_5455 ( .C ( clk ), .D ( signal_11046 ), .Q ( signal_11047 ) ) ;
    buf_clk cell_5463 ( .C ( clk ), .D ( signal_11054 ), .Q ( signal_11055 ) ) ;
    buf_clk cell_5487 ( .C ( clk ), .D ( signal_2030 ), .Q ( signal_11079 ) ) ;
    buf_clk cell_5495 ( .C ( clk ), .D ( signal_4584 ), .Q ( signal_11087 ) ) ;
    buf_clk cell_5503 ( .C ( clk ), .D ( signal_4585 ), .Q ( signal_11095 ) ) ;
    buf_clk cell_5547 ( .C ( clk ), .D ( signal_9466 ), .Q ( signal_11139 ) ) ;
    buf_clk cell_5555 ( .C ( clk ), .D ( signal_9468 ), .Q ( signal_11147 ) ) ;
    buf_clk cell_5563 ( .C ( clk ), .D ( signal_9470 ), .Q ( signal_11155 ) ) ;
    buf_clk cell_5573 ( .C ( clk ), .D ( signal_11164 ), .Q ( signal_11165 ) ) ;
    buf_clk cell_5583 ( .C ( clk ), .D ( signal_11174 ), .Q ( signal_11175 ) ) ;
    buf_clk cell_5593 ( .C ( clk ), .D ( signal_11184 ), .Q ( signal_11185 ) ) ;
    buf_clk cell_5625 ( .C ( clk ), .D ( signal_1982 ), .Q ( signal_11217 ) ) ;
    buf_clk cell_5633 ( .C ( clk ), .D ( signal_4488 ), .Q ( signal_11225 ) ) ;
    buf_clk cell_5641 ( .C ( clk ), .D ( signal_4489 ), .Q ( signal_11233 ) ) ;
    buf_clk cell_5651 ( .C ( clk ), .D ( signal_11242 ), .Q ( signal_11243 ) ) ;
    buf_clk cell_5661 ( .C ( clk ), .D ( signal_11252 ), .Q ( signal_11253 ) ) ;
    buf_clk cell_5671 ( .C ( clk ), .D ( signal_11262 ), .Q ( signal_11263 ) ) ;
    buf_clk cell_5679 ( .C ( clk ), .D ( signal_1967 ), .Q ( signal_11271 ) ) ;
    buf_clk cell_5687 ( .C ( clk ), .D ( signal_4458 ), .Q ( signal_11279 ) ) ;
    buf_clk cell_5695 ( .C ( clk ), .D ( signal_4459 ), .Q ( signal_11287 ) ) ;
    buf_clk cell_5919 ( .C ( clk ), .D ( signal_1978 ), .Q ( signal_11511 ) ) ;
    buf_clk cell_5929 ( .C ( clk ), .D ( signal_4480 ), .Q ( signal_11521 ) ) ;
    buf_clk cell_5939 ( .C ( clk ), .D ( signal_4481 ), .Q ( signal_11531 ) ) ;
    buf_clk cell_6183 ( .C ( clk ), .D ( signal_1736 ), .Q ( signal_11775 ) ) ;
    buf_clk cell_6195 ( .C ( clk ), .D ( signal_3996 ), .Q ( signal_11787 ) ) ;
    buf_clk cell_6207 ( .C ( clk ), .D ( signal_3997 ), .Q ( signal_11799 ) ) ;
    buf_clk cell_6257 ( .C ( clk ), .D ( signal_11848 ), .Q ( signal_11849 ) ) ;
    buf_clk cell_6271 ( .C ( clk ), .D ( signal_11862 ), .Q ( signal_11863 ) ) ;
    buf_clk cell_6285 ( .C ( clk ), .D ( signal_11876 ), .Q ( signal_11877 ) ) ;
    buf_clk cell_6323 ( .C ( clk ), .D ( signal_11914 ), .Q ( signal_11915 ) ) ;
    buf_clk cell_6337 ( .C ( clk ), .D ( signal_11928 ), .Q ( signal_11929 ) ) ;
    buf_clk cell_6351 ( .C ( clk ), .D ( signal_11942 ), .Q ( signal_11943 ) ) ;
    buf_clk cell_6443 ( .C ( clk ), .D ( signal_12034 ), .Q ( signal_12035 ) ) ;
    buf_clk cell_6459 ( .C ( clk ), .D ( signal_12050 ), .Q ( signal_12051 ) ) ;
    buf_clk cell_6475 ( .C ( clk ), .D ( signal_12066 ), .Q ( signal_12067 ) ) ;
    buf_clk cell_6503 ( .C ( clk ), .D ( signal_12094 ), .Q ( signal_12095 ) ) ;
    buf_clk cell_6519 ( .C ( clk ), .D ( signal_12110 ), .Q ( signal_12111 ) ) ;
    buf_clk cell_6535 ( .C ( clk ), .D ( signal_12126 ), .Q ( signal_12127 ) ) ;
    buf_clk cell_6687 ( .C ( clk ), .D ( signal_1783 ), .Q ( signal_12279 ) ) ;
    buf_clk cell_6703 ( .C ( clk ), .D ( signal_4090 ), .Q ( signal_12295 ) ) ;
    buf_clk cell_6719 ( .C ( clk ), .D ( signal_4091 ), .Q ( signal_12311 ) ) ;
    buf_clk cell_6737 ( .C ( clk ), .D ( signal_12328 ), .Q ( signal_12329 ) ) ;
    buf_clk cell_6755 ( .C ( clk ), .D ( signal_12346 ), .Q ( signal_12347 ) ) ;
    buf_clk cell_6773 ( .C ( clk ), .D ( signal_12364 ), .Q ( signal_12365 ) ) ;
    buf_clk cell_6887 ( .C ( clk ), .D ( signal_12478 ), .Q ( signal_12479 ) ) ;
    buf_clk cell_6907 ( .C ( clk ), .D ( signal_12498 ), .Q ( signal_12499 ) ) ;
    buf_clk cell_6927 ( .C ( clk ), .D ( signal_12518 ), .Q ( signal_12519 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1819 ( .a ({signal_8930, signal_8928, signal_8926}), .b ({signal_3899, signal_3898, signal_1687}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743]}), .c ({signal_4193, signal_4192, signal_1834}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1834 ( .a ({signal_8936, signal_8934, signal_8932}), .b ({signal_3945, signal_3944, signal_1710}), .clk ( clk ), .r ({Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({signal_4223, signal_4222, signal_1849}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1872 ( .a ({signal_4193, signal_4192, signal_1834}), .b ({signal_4299, signal_4298, signal_1887}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1875 ( .a ({signal_4223, signal_4222, signal_1849}), .b ({signal_4305, signal_4304, signal_1890}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1893 ( .a ({signal_8948, signal_8944, signal_8940}), .b ({signal_3985, signal_3984, signal_1730}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749]}), .c ({signal_4341, signal_4340, signal_1908}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1902 ( .a ({signal_4059, signal_4058, signal_1767}), .b ({signal_4097, signal_4096, signal_1786}), .clk ( clk ), .r ({Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({signal_4359, signal_4358, signal_1917}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1904 ( .a ({signal_8948, signal_8944, signal_8940}), .b ({signal_4005, signal_4004, signal_1740}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755]}), .c ({signal_4363, signal_4362, signal_1919}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1911 ( .a ({signal_4105, signal_4104, signal_1790}), .b ({signal_8954, signal_8952, signal_8950}), .clk ( clk ), .r ({Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({signal_4377, signal_4376, signal_1926}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1912 ( .a ({signal_8966, signal_8962, signal_8958}), .b ({signal_4109, signal_4108, signal_1792}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761]}), .c ({signal_4379, signal_4378, signal_1927}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1918 ( .a ({signal_8978, signal_8974, signal_8970}), .b ({signal_4133, signal_4132, signal_1804}), .clk ( clk ), .r ({Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({signal_4391, signal_4390, signal_1933}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1921 ( .a ({signal_8990, signal_8986, signal_8982}), .b ({signal_4137, signal_4136, signal_1806}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767]}), .c ({signal_4397, signal_4396, signal_1936}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1922 ( .a ({signal_4141, signal_4140, signal_1808}), .b ({signal_4143, signal_4142, signal_1809}), .clk ( clk ), .r ({Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_4399, signal_4398, signal_1937}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1924 ( .a ({signal_9014, signal_9006, signal_8998}), .b ({signal_4029, signal_4028, signal_1752}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773]}), .c ({signal_4403, signal_4402, signal_1939}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1925 ( .a ({signal_9020, signal_9018, signal_9016}), .b ({signal_4155, signal_4154, signal_1815}), .clk ( clk ), .r ({Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({signal_4405, signal_4404, signal_1940}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1926 ( .a ({signal_9026, signal_9024, signal_9022}), .b ({signal_4031, signal_4030, signal_1753}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779]}), .c ({signal_4407, signal_4406, signal_1941}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1928 ( .a ({signal_9038, signal_9034, signal_9030}), .b ({signal_4163, signal_4162, signal_1819}), .clk ( clk ), .r ({Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({signal_4411, signal_4410, signal_1943}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1929 ( .a ({signal_4103, signal_4102, signal_1789}), .b ({signal_9044, signal_9042, signal_9040}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785]}), .c ({signal_4413, signal_4412, signal_1944}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1930 ( .a ({signal_4037, signal_4036, signal_1756}), .b ({signal_4039, signal_4038, signal_1757}), .clk ( clk ), .r ({Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({signal_4415, signal_4414, signal_1945}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1931 ( .a ({signal_9050, signal_9048, signal_9046}), .b ({signal_4043, signal_4042, signal_1759}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791]}), .c ({signal_4417, signal_4416, signal_1946}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1933 ( .a ({signal_9062, signal_9058, signal_9054}), .b ({signal_4179, signal_4178, signal_1827}), .clk ( clk ), .r ({Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({signal_4421, signal_4420, signal_1948}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1934 ( .a ({signal_9068, signal_9066, signal_9064}), .b ({signal_4191, signal_4190, signal_1833}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797]}), .c ({signal_4423, signal_4422, signal_1949}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1935 ( .a ({signal_9074, signal_9072, signal_9070}), .b ({signal_4195, signal_4194, signal_1835}), .clk ( clk ), .r ({Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_4425, signal_4424, signal_1950}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1936 ( .a ({signal_4047, signal_4046, signal_1761}), .b ({signal_4197, signal_4196, signal_1836}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803]}), .c ({signal_4427, signal_4426, signal_1951}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1937 ( .a ({signal_9080, signal_9078, signal_9076}), .b ({signal_4035, signal_4034, signal_1755}), .clk ( clk ), .r ({Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({signal_4429, signal_4428, signal_1952}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1938 ( .a ({signal_9086, signal_9084, signal_9082}), .b ({signal_4199, signal_4198, signal_1837}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809]}), .c ({signal_4431, signal_4430, signal_1953}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1939 ( .a ({signal_9092, signal_9090, signal_9088}), .b ({signal_4201, signal_4200, signal_1838}), .clk ( clk ), .r ({Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({signal_4433, signal_4432, signal_1954}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1940 ( .a ({signal_9104, signal_9100, signal_9096}), .b ({signal_4205, signal_4204, signal_1840}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815]}), .c ({signal_4435, signal_4434, signal_1955}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1941 ( .a ({signal_9110, signal_9108, signal_9106}), .b ({signal_4051, signal_4050, signal_1763}), .clk ( clk ), .r ({Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({signal_4437, signal_4436, signal_1956}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1942 ( .a ({signal_9116, signal_9114, signal_9112}), .b ({signal_4207, signal_4206, signal_1841}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821]}), .c ({signal_4439, signal_4438, signal_1957}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1943 ( .a ({signal_4131, signal_4130, signal_1803}), .b ({signal_9122, signal_9120, signal_9118}), .clk ( clk ), .r ({Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({signal_4441, signal_4440, signal_1958}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1945 ( .a ({signal_4175, signal_4174, signal_1825}), .b ({signal_4217, signal_4216, signal_1846}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827]}), .c ({signal_4445, signal_4444, signal_1960}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1946 ( .a ({signal_9128, signal_9126, signal_9124}), .b ({signal_4055, signal_4054, signal_1765}), .clk ( clk ), .r ({Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_4447, signal_4446, signal_1961}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1947 ( .a ({signal_4117, signal_4116, signal_1796}), .b ({signal_4219, signal_4218, signal_1847}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833]}), .c ({signal_4449, signal_4448, signal_1962}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1961 ( .a ({signal_4341, signal_4340, signal_1908}), .b ({signal_4477, signal_4476, signal_1976}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1969 ( .a ({signal_4359, signal_4358, signal_1917}), .b ({signal_4493, signal_4492, signal_1984}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1971 ( .a ({signal_4363, signal_4362, signal_1919}), .b ({signal_4497, signal_4496, signal_1986}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1978 ( .a ({signal_4379, signal_4378, signal_1927}), .b ({signal_4511, signal_4510, signal_1993}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1986 ( .a ({signal_4397, signal_4396, signal_1936}), .b ({signal_4527, signal_4526, signal_2001}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1987 ( .a ({signal_4399, signal_4398, signal_1937}), .b ({signal_4529, signal_4528, signal_2002}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1989 ( .a ({signal_4403, signal_4402, signal_1939}), .b ({signal_4533, signal_4532, signal_2004}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1992 ( .a ({signal_4423, signal_4422, signal_1949}), .b ({signal_4539, signal_4538, signal_2007}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1993 ( .a ({signal_4427, signal_4426, signal_1951}), .b ({signal_4541, signal_4540, signal_2008}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1994 ( .a ({signal_4439, signal_4438, signal_1957}), .b ({signal_4543, signal_4542, signal_2009}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1995 ( .a ({signal_4441, signal_4440, signal_1958}), .b ({signal_4545, signal_4544, signal_2010}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1997 ( .a ({signal_4445, signal_4444, signal_1960}), .b ({signal_4549, signal_4548, signal_2012}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_1998 ( .a ({signal_4449, signal_4448, signal_1962}), .b ({signal_4551, signal_4550, signal_2013}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_1999 ( .a ({signal_4239, signal_4238, signal_1857}), .b ({signal_9140, signal_9136, signal_9132}), .clk ( clk ), .r ({Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({signal_4553, signal_4552, signal_2014}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2002 ( .a ({signal_9146, signal_9144, signal_9142}), .b ({signal_4073, signal_4072, signal_1774}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839]}), .c ({signal_4559, signal_4558, signal_2017}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2007 ( .a ({signal_9152, signal_9150, signal_9148}), .b ({signal_4313, signal_4312, signal_1894}), .clk ( clk ), .r ({Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({signal_4569, signal_4568, signal_2022}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2009 ( .a ({signal_9164, signal_9160, signal_9156}), .b ({signal_4317, signal_4316, signal_1896}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845]}), .c ({signal_4573, signal_4572, signal_2024}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2010 ( .a ({signal_9176, signal_9172, signal_9168}), .b ({signal_4323, signal_4322, signal_1899}), .clk ( clk ), .r ({Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({signal_4575, signal_4574, signal_2025}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2013 ( .a ({signal_9188, signal_9184, signal_9180}), .b ({signal_4261, signal_4260, signal_1868}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851]}), .c ({signal_4581, signal_4580, signal_2028}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2016 ( .a ({signal_9200, signal_9196, signal_9192}), .b ({signal_4273, signal_4272, signal_1874}), .clk ( clk ), .r ({Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({signal_4587, signal_4586, signal_2031}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2017 ( .a ({signal_9206, signal_9204, signal_9202}), .b ({signal_4275, signal_4274, signal_1875}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857]}), .c ({signal_4589, signal_4588, signal_2032}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2018 ( .a ({signal_9212, signal_9210, signal_9208}), .b ({signal_4277, signal_4276, signal_1876}), .clk ( clk ), .r ({Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_4591, signal_4590, signal_2033}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2019 ( .a ({signal_9218, signal_9216, signal_9214}), .b ({signal_4151, signal_4150, signal_1813}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863]}), .c ({signal_4593, signal_4592, signal_2034}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2020 ( .a ({signal_9224, signal_9222, signal_9220}), .b ({signal_4279, signal_4278, signal_1877}), .clk ( clk ), .r ({Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({signal_4595, signal_4594, signal_2035}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2021 ( .a ({signal_9230, signal_9228, signal_9226}), .b ({signal_4281, signal_4280, signal_1878}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869]}), .c ({signal_4597, signal_4596, signal_2036}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2022 ( .a ({signal_9242, signal_9238, signal_9234}), .b ({signal_4283, signal_4282, signal_1879}), .clk ( clk ), .r ({Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({signal_4599, signal_4598, signal_2037}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2023 ( .a ({signal_9254, signal_9250, signal_9246}), .b ({signal_4285, signal_4284, signal_1880}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875]}), .c ({signal_4601, signal_4600, signal_2038}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2024 ( .a ({signal_9266, signal_9262, signal_9258}), .b ({signal_4287, signal_4286, signal_1881}), .clk ( clk ), .r ({Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({signal_4603, signal_4602, signal_2039}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2025 ( .a ({signal_9272, signal_9270, signal_9268}), .b ({signal_4289, signal_4288, signal_1882}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881]}), .c ({signal_4605, signal_4604, signal_2040}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2026 ( .a ({signal_4177, signal_4176, signal_1826}), .b ({signal_4357, signal_4356, signal_1916}), .clk ( clk ), .r ({Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({signal_4607, signal_4606, signal_2041}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2028 ( .a ({signal_9284, signal_9280, signal_9276}), .b ({signal_4291, signal_4290, signal_1883}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887]}), .c ({signal_4611, signal_4610, signal_2043}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2029 ( .a ({signal_9290, signal_9288, signal_9286}), .b ({signal_4293, signal_4292, signal_1884}), .clk ( clk ), .r ({Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_4613, signal_4612, signal_2044}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2030 ( .a ({signal_9296, signal_9294, signal_9292}), .b ({signal_4185, signal_4184, signal_1830}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893]}), .c ({signal_4615, signal_4614, signal_2045}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2031 ( .a ({signal_9302, signal_9300, signal_9298}), .b ({signal_4297, signal_4296, signal_1886}), .clk ( clk ), .r ({Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({signal_4617, signal_4616, signal_2046}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2033 ( .a ({signal_9308, signal_9306, signal_9304}), .b ({signal_4203, signal_4202, signal_1839}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899]}), .c ({signal_4621, signal_4620, signal_2048}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2034 ( .a ({signal_9314, signal_9312, signal_9310}), .b ({signal_4161, signal_4160, signal_1818}), .clk ( clk ), .r ({Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({signal_4623, signal_4622, signal_2049}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2035 ( .a ({signal_9326, signal_9322, signal_9318}), .b ({signal_4301, signal_4300, signal_1888}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905]}), .c ({signal_4625, signal_4624, signal_2050}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2036 ( .a ({signal_9164, signal_9160, signal_9156}), .b ({signal_4303, signal_4302, signal_1889}), .clk ( clk ), .r ({Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({signal_4627, signal_4626, signal_2051}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2046 ( .a ({signal_4553, signal_4552, signal_2014}), .b ({signal_4647, signal_4646, signal_2061}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2047 ( .a ({signal_4559, signal_4558, signal_2017}), .b ({signal_4649, signal_4648, signal_2062}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2049 ( .a ({signal_4569, signal_4568, signal_2022}), .b ({signal_4653, signal_4652, signal_2064}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2050 ( .a ({signal_4573, signal_4572, signal_2024}), .b ({signal_4655, signal_4654, signal_2065}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2051 ( .a ({signal_4575, signal_4574, signal_2025}), .b ({signal_4657, signal_4656, signal_2066}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2053 ( .a ({signal_4581, signal_4580, signal_2028}), .b ({signal_4661, signal_4660, signal_2068}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2054 ( .a ({signal_4587, signal_4586, signal_2031}), .b ({signal_4663, signal_4662, signal_2069}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2055 ( .a ({signal_4589, signal_4588, signal_2032}), .b ({signal_4665, signal_4664, signal_2070}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2056 ( .a ({signal_4591, signal_4590, signal_2033}), .b ({signal_4667, signal_4666, signal_2071}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2057 ( .a ({signal_4593, signal_4592, signal_2034}), .b ({signal_4669, signal_4668, signal_2072}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2058 ( .a ({signal_4595, signal_4594, signal_2035}), .b ({signal_4671, signal_4670, signal_2073}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2059 ( .a ({signal_4597, signal_4596, signal_2036}), .b ({signal_4673, signal_4672, signal_2074}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2060 ( .a ({signal_4599, signal_4598, signal_2037}), .b ({signal_4675, signal_4674, signal_2075}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2061 ( .a ({signal_4601, signal_4600, signal_2038}), .b ({signal_4677, signal_4676, signal_2076}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2062 ( .a ({signal_4603, signal_4602, signal_2039}), .b ({signal_4679, signal_4678, signal_2077}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2063 ( .a ({signal_4607, signal_4606, signal_2041}), .b ({signal_4681, signal_4680, signal_2078}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2065 ( .a ({signal_4611, signal_4610, signal_2043}), .b ({signal_4685, signal_4684, signal_2080}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2066 ( .a ({signal_4613, signal_4612, signal_2044}), .b ({signal_4687, signal_4686, signal_2081}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2067 ( .a ({signal_4617, signal_4616, signal_2046}), .b ({signal_4689, signal_4688, signal_2082}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2069 ( .a ({signal_4621, signal_4620, signal_2048}), .b ({signal_4693, signal_4692, signal_2084}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2070 ( .a ({signal_4625, signal_4624, signal_2050}), .b ({signal_4695, signal_4694, signal_2085}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2071 ( .a ({signal_4627, signal_4626, signal_2051}), .b ({signal_4697, signal_4696, signal_2086}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2074 ( .a ({signal_4479, signal_4478, signal_1977}), .b ({signal_9338, signal_9334, signal_9330}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911]}), .c ({signal_4703, signal_4702, signal_2089}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2075 ( .a ({signal_9344, signal_9342, signal_9340}), .b ({signal_4453, signal_4452, signal_1964}), .clk ( clk ), .r ({Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({signal_4705, signal_4704, signal_2090}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2076 ( .a ({signal_9356, signal_9352, signal_9348}), .b ({signal_4555, signal_4554, signal_2015}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917]}), .c ({signal_4707, signal_4706, signal_2091}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2077 ( .a ({signal_9362, signal_9360, signal_9358}), .b ({signal_4463, signal_4462, signal_1969}), .clk ( clk ), .r ({Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_4709, signal_4708, signal_2092}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2078 ( .a ({signal_4451, signal_4450, signal_1963}), .b ({signal_9368, signal_9366, signal_9364}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923]}), .c ({signal_4711, signal_4710, signal_2093}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2079 ( .a ({signal_4471, signal_4470, signal_1973}), .b ({signal_4473, signal_4472, signal_1974}), .clk ( clk ), .r ({Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({signal_4713, signal_4712, signal_2094}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2080 ( .a ({signal_9380, signal_9376, signal_9372}), .b ({signal_4561, signal_4560, signal_2018}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929]}), .c ({signal_4715, signal_4714, signal_2095}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2081 ( .a ({signal_9392, signal_9388, signal_9384}), .b ({signal_4565, signal_4564, signal_2020}), .clk ( clk ), .r ({Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({signal_4717, signal_4716, signal_2096}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2082 ( .a ({signal_9404, signal_9400, signal_9396}), .b ({signal_4567, signal_4566, signal_2021}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935]}), .c ({signal_4719, signal_4718, signal_2097}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2083 ( .a ({signal_9410, signal_9408, signal_9406}), .b ({signal_4487, signal_4486, signal_1981}), .clk ( clk ), .r ({Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({signal_4721, signal_4720, signal_2098}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2085 ( .a ({signal_9422, signal_9418, signal_9414}), .b ({signal_4495, signal_4494, signal_1985}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941]}), .c ({signal_4725, signal_4724, signal_2100}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2086 ( .a ({signal_9434, signal_9430, signal_9426}), .b ({signal_4571, signal_4570, signal_2023}), .clk ( clk ), .r ({Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({signal_4727, signal_4726, signal_2101}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2087 ( .a ({signal_4307, signal_4306, signal_1891}), .b ({signal_4503, signal_4502, signal_1989}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947]}), .c ({signal_4729, signal_4728, signal_2102}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2088 ( .a ({signal_4505, signal_4504, signal_1990}), .b ({signal_4507, signal_4506, signal_1991}), .clk ( clk ), .r ({Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_4731, signal_4730, signal_2103}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2089 ( .a ({signal_9440, signal_9438, signal_9436}), .b ({signal_4509, signal_4508, signal_1992}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953]}), .c ({signal_4733, signal_4732, signal_2104}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2091 ( .a ({signal_4579, signal_4578, signal_2027}), .b ({signal_4295, signal_4294, signal_1885}), .clk ( clk ), .r ({Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({signal_4737, signal_4736, signal_2106}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2092 ( .a ({signal_9452, signal_9448, signal_9444}), .b ({signal_4513, signal_4512, signal_1994}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959]}), .c ({signal_4739, signal_4738, signal_2107}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2093 ( .a ({signal_9458, signal_9456, signal_9454}), .b ({signal_4515, signal_4514, signal_1995}), .clk ( clk ), .r ({Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({signal_4741, signal_4740, signal_2108}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2094 ( .a ({signal_4129, signal_4128, signal_1802}), .b ({signal_4517, signal_4516, signal_1996}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965]}), .c ({signal_4743, signal_4742, signal_2109}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2095 ( .a ({signal_4467, signal_4466, signal_1971}), .b ({signal_4519, signal_4518, signal_1997}), .clk ( clk ), .r ({Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({signal_4745, signal_4744, signal_2110}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2096 ( .a ({signal_4037, signal_4036, signal_1756}), .b ({signal_4521, signal_4520, signal_1998}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971]}), .c ({signal_4747, signal_4746, signal_2111}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2097 ( .a ({signal_4469, signal_4468, signal_1972}), .b ({signal_9044, signal_9042, signal_9040}), .clk ( clk ), .r ({Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({signal_4749, signal_4748, signal_2112}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2099 ( .a ({signal_3921, signal_3920, signal_1698}), .b ({signal_4525, signal_4524, signal_2000}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977]}), .c ({signal_4753, signal_4752, signal_2114}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2101 ( .a ({signal_4475, signal_4474, signal_1975}), .b ({signal_4531, signal_4530, signal_2003}), .clk ( clk ), .r ({Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_4757, signal_4756, signal_2116}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2104 ( .a ({signal_9464, signal_9462, signal_9460}), .b ({signal_4535, signal_4534, signal_2005}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983]}), .c ({signal_4763, signal_4762, signal_2119}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2110 ( .a ({signal_4583, signal_4582, signal_2029}), .b ({signal_4221, signal_4220, signal_1848}), .clk ( clk ), .r ({Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({signal_4775, signal_4774, signal_2125}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2124 ( .a ({signal_4703, signal_4702, signal_2089}), .b ({signal_4803, signal_4802, signal_2139}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2125 ( .a ({signal_4707, signal_4706, signal_2091}), .b ({signal_4805, signal_4804, signal_2140}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2126 ( .a ({signal_4709, signal_4708, signal_2092}), .b ({signal_4807, signal_4806, signal_2141}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2127 ( .a ({signal_4717, signal_4716, signal_2096}), .b ({signal_4809, signal_4808, signal_2142}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2128 ( .a ({signal_4719, signal_4718, signal_2097}), .b ({signal_4811, signal_4810, signal_2143}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2130 ( .a ({signal_4727, signal_4726, signal_2101}), .b ({signal_4815, signal_4814, signal_2145}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2133 ( .a ({signal_4763, signal_4762, signal_2119}), .b ({signal_4821, signal_4820, signal_2148}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2135 ( .a ({signal_4775, signal_4774, signal_2125}), .b ({signal_4825, signal_4824, signal_2150}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2144 ( .a ({signal_9470, signal_9468, signal_9466}), .b ({signal_4651, signal_4650, signal_2063}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989]}), .c ({signal_4843, signal_4842, signal_2159}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2148 ( .a ({signal_9482, signal_9478, signal_9474}), .b ({signal_4659, signal_4658, signal_2067}), .clk ( clk ), .r ({Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({signal_4851, signal_4850, signal_2163}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2185 ( .a ({signal_4843, signal_4842, signal_2159}), .b ({signal_4925, signal_4924, signal_2200}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2186 ( .a ({signal_4851, signal_4850, signal_2163}), .b ({signal_4927, signal_4926, signal_2201}) ) ;
    buf_clk cell_3892 ( .C ( clk ), .D ( signal_9483 ), .Q ( signal_9484 ) ) ;
    buf_clk cell_3894 ( .C ( clk ), .D ( signal_9485 ), .Q ( signal_9486 ) ) ;
    buf_clk cell_3896 ( .C ( clk ), .D ( signal_9487 ), .Q ( signal_9488 ) ) ;
    buf_clk cell_3902 ( .C ( clk ), .D ( signal_9493 ), .Q ( signal_9494 ) ) ;
    buf_clk cell_3908 ( .C ( clk ), .D ( signal_9499 ), .Q ( signal_9500 ) ) ;
    buf_clk cell_3914 ( .C ( clk ), .D ( signal_9505 ), .Q ( signal_9506 ) ) ;
    buf_clk cell_3920 ( .C ( clk ), .D ( signal_9511 ), .Q ( signal_9512 ) ) ;
    buf_clk cell_3926 ( .C ( clk ), .D ( signal_9517 ), .Q ( signal_9518 ) ) ;
    buf_clk cell_3932 ( .C ( clk ), .D ( signal_9523 ), .Q ( signal_9524 ) ) ;
    buf_clk cell_3938 ( .C ( clk ), .D ( signal_9529 ), .Q ( signal_9530 ) ) ;
    buf_clk cell_3944 ( .C ( clk ), .D ( signal_9535 ), .Q ( signal_9536 ) ) ;
    buf_clk cell_3950 ( .C ( clk ), .D ( signal_9541 ), .Q ( signal_9542 ) ) ;
    buf_clk cell_3954 ( .C ( clk ), .D ( signal_9545 ), .Q ( signal_9546 ) ) ;
    buf_clk cell_3958 ( .C ( clk ), .D ( signal_9549 ), .Q ( signal_9550 ) ) ;
    buf_clk cell_3962 ( .C ( clk ), .D ( signal_9553 ), .Q ( signal_9554 ) ) ;
    buf_clk cell_3968 ( .C ( clk ), .D ( signal_9559 ), .Q ( signal_9560 ) ) ;
    buf_clk cell_3974 ( .C ( clk ), .D ( signal_9565 ), .Q ( signal_9566 ) ) ;
    buf_clk cell_3980 ( .C ( clk ), .D ( signal_9571 ), .Q ( signal_9572 ) ) ;
    buf_clk cell_3984 ( .C ( clk ), .D ( signal_9575 ), .Q ( signal_9576 ) ) ;
    buf_clk cell_3988 ( .C ( clk ), .D ( signal_9579 ), .Q ( signal_9580 ) ) ;
    buf_clk cell_3992 ( .C ( clk ), .D ( signal_9583 ), .Q ( signal_9584 ) ) ;
    buf_clk cell_3996 ( .C ( clk ), .D ( signal_9587 ), .Q ( signal_9588 ) ) ;
    buf_clk cell_4000 ( .C ( clk ), .D ( signal_9591 ), .Q ( signal_9592 ) ) ;
    buf_clk cell_4004 ( .C ( clk ), .D ( signal_9595 ), .Q ( signal_9596 ) ) ;
    buf_clk cell_4008 ( .C ( clk ), .D ( signal_9599 ), .Q ( signal_9600 ) ) ;
    buf_clk cell_4012 ( .C ( clk ), .D ( signal_9603 ), .Q ( signal_9604 ) ) ;
    buf_clk cell_4016 ( .C ( clk ), .D ( signal_9607 ), .Q ( signal_9608 ) ) ;
    buf_clk cell_4020 ( .C ( clk ), .D ( signal_9611 ), .Q ( signal_9612 ) ) ;
    buf_clk cell_4024 ( .C ( clk ), .D ( signal_9615 ), .Q ( signal_9616 ) ) ;
    buf_clk cell_4028 ( .C ( clk ), .D ( signal_9619 ), .Q ( signal_9620 ) ) ;
    buf_clk cell_4032 ( .C ( clk ), .D ( signal_9623 ), .Q ( signal_9624 ) ) ;
    buf_clk cell_4036 ( .C ( clk ), .D ( signal_9627 ), .Q ( signal_9628 ) ) ;
    buf_clk cell_4040 ( .C ( clk ), .D ( signal_9631 ), .Q ( signal_9632 ) ) ;
    buf_clk cell_4046 ( .C ( clk ), .D ( signal_9637 ), .Q ( signal_9638 ) ) ;
    buf_clk cell_4052 ( .C ( clk ), .D ( signal_9643 ), .Q ( signal_9644 ) ) ;
    buf_clk cell_4058 ( .C ( clk ), .D ( signal_9649 ), .Q ( signal_9650 ) ) ;
    buf_clk cell_4062 ( .C ( clk ), .D ( signal_9653 ), .Q ( signal_9654 ) ) ;
    buf_clk cell_4066 ( .C ( clk ), .D ( signal_9657 ), .Q ( signal_9658 ) ) ;
    buf_clk cell_4070 ( .C ( clk ), .D ( signal_9661 ), .Q ( signal_9662 ) ) ;
    buf_clk cell_4072 ( .C ( clk ), .D ( signal_9663 ), .Q ( signal_9664 ) ) ;
    buf_clk cell_4074 ( .C ( clk ), .D ( signal_9665 ), .Q ( signal_9666 ) ) ;
    buf_clk cell_4076 ( .C ( clk ), .D ( signal_9667 ), .Q ( signal_9668 ) ) ;
    buf_clk cell_4078 ( .C ( clk ), .D ( signal_9669 ), .Q ( signal_9670 ) ) ;
    buf_clk cell_4080 ( .C ( clk ), .D ( signal_9671 ), .Q ( signal_9672 ) ) ;
    buf_clk cell_4082 ( .C ( clk ), .D ( signal_9673 ), .Q ( signal_9674 ) ) ;
    buf_clk cell_4084 ( .C ( clk ), .D ( signal_9675 ), .Q ( signal_9676 ) ) ;
    buf_clk cell_4086 ( .C ( clk ), .D ( signal_9677 ), .Q ( signal_9678 ) ) ;
    buf_clk cell_4088 ( .C ( clk ), .D ( signal_9679 ), .Q ( signal_9680 ) ) ;
    buf_clk cell_4090 ( .C ( clk ), .D ( signal_9681 ), .Q ( signal_9682 ) ) ;
    buf_clk cell_4092 ( .C ( clk ), .D ( signal_9683 ), .Q ( signal_9684 ) ) ;
    buf_clk cell_4094 ( .C ( clk ), .D ( signal_9685 ), .Q ( signal_9686 ) ) ;
    buf_clk cell_4096 ( .C ( clk ), .D ( signal_9687 ), .Q ( signal_9688 ) ) ;
    buf_clk cell_4098 ( .C ( clk ), .D ( signal_9689 ), .Q ( signal_9690 ) ) ;
    buf_clk cell_4100 ( .C ( clk ), .D ( signal_9691 ), .Q ( signal_9692 ) ) ;
    buf_clk cell_4104 ( .C ( clk ), .D ( signal_9695 ), .Q ( signal_9696 ) ) ;
    buf_clk cell_4108 ( .C ( clk ), .D ( signal_9699 ), .Q ( signal_9700 ) ) ;
    buf_clk cell_4112 ( .C ( clk ), .D ( signal_9703 ), .Q ( signal_9704 ) ) ;
    buf_clk cell_4114 ( .C ( clk ), .D ( signal_9705 ), .Q ( signal_9706 ) ) ;
    buf_clk cell_4116 ( .C ( clk ), .D ( signal_9707 ), .Q ( signal_9708 ) ) ;
    buf_clk cell_4118 ( .C ( clk ), .D ( signal_9709 ), .Q ( signal_9710 ) ) ;
    buf_clk cell_4120 ( .C ( clk ), .D ( signal_9711 ), .Q ( signal_9712 ) ) ;
    buf_clk cell_4122 ( .C ( clk ), .D ( signal_9713 ), .Q ( signal_9714 ) ) ;
    buf_clk cell_4124 ( .C ( clk ), .D ( signal_9715 ), .Q ( signal_9716 ) ) ;
    buf_clk cell_4126 ( .C ( clk ), .D ( signal_9717 ), .Q ( signal_9718 ) ) ;
    buf_clk cell_4128 ( .C ( clk ), .D ( signal_9719 ), .Q ( signal_9720 ) ) ;
    buf_clk cell_4130 ( .C ( clk ), .D ( signal_9721 ), .Q ( signal_9722 ) ) ;
    buf_clk cell_4136 ( .C ( clk ), .D ( signal_9727 ), .Q ( signal_9728 ) ) ;
    buf_clk cell_4142 ( .C ( clk ), .D ( signal_9733 ), .Q ( signal_9734 ) ) ;
    buf_clk cell_4148 ( .C ( clk ), .D ( signal_9739 ), .Q ( signal_9740 ) ) ;
    buf_clk cell_4150 ( .C ( clk ), .D ( signal_9741 ), .Q ( signal_9742 ) ) ;
    buf_clk cell_4152 ( .C ( clk ), .D ( signal_9743 ), .Q ( signal_9744 ) ) ;
    buf_clk cell_4154 ( .C ( clk ), .D ( signal_9745 ), .Q ( signal_9746 ) ) ;
    buf_clk cell_4158 ( .C ( clk ), .D ( signal_9749 ), .Q ( signal_9750 ) ) ;
    buf_clk cell_4162 ( .C ( clk ), .D ( signal_9753 ), .Q ( signal_9754 ) ) ;
    buf_clk cell_4166 ( .C ( clk ), .D ( signal_9757 ), .Q ( signal_9758 ) ) ;
    buf_clk cell_4168 ( .C ( clk ), .D ( signal_9759 ), .Q ( signal_9760 ) ) ;
    buf_clk cell_4170 ( .C ( clk ), .D ( signal_9761 ), .Q ( signal_9762 ) ) ;
    buf_clk cell_4172 ( .C ( clk ), .D ( signal_9763 ), .Q ( signal_9764 ) ) ;
    buf_clk cell_4174 ( .C ( clk ), .D ( signal_9765 ), .Q ( signal_9766 ) ) ;
    buf_clk cell_4176 ( .C ( clk ), .D ( signal_9767 ), .Q ( signal_9768 ) ) ;
    buf_clk cell_4178 ( .C ( clk ), .D ( signal_9769 ), .Q ( signal_9770 ) ) ;
    buf_clk cell_4184 ( .C ( clk ), .D ( signal_9775 ), .Q ( signal_9776 ) ) ;
    buf_clk cell_4190 ( .C ( clk ), .D ( signal_9781 ), .Q ( signal_9782 ) ) ;
    buf_clk cell_4196 ( .C ( clk ), .D ( signal_9787 ), .Q ( signal_9788 ) ) ;
    buf_clk cell_4200 ( .C ( clk ), .D ( signal_9791 ), .Q ( signal_9792 ) ) ;
    buf_clk cell_4204 ( .C ( clk ), .D ( signal_9795 ), .Q ( signal_9796 ) ) ;
    buf_clk cell_4208 ( .C ( clk ), .D ( signal_9799 ), .Q ( signal_9800 ) ) ;
    buf_clk cell_4210 ( .C ( clk ), .D ( signal_9801 ), .Q ( signal_9802 ) ) ;
    buf_clk cell_4212 ( .C ( clk ), .D ( signal_9803 ), .Q ( signal_9804 ) ) ;
    buf_clk cell_4214 ( .C ( clk ), .D ( signal_9805 ), .Q ( signal_9806 ) ) ;
    buf_clk cell_4216 ( .C ( clk ), .D ( signal_9807 ), .Q ( signal_9808 ) ) ;
    buf_clk cell_4218 ( .C ( clk ), .D ( signal_9809 ), .Q ( signal_9810 ) ) ;
    buf_clk cell_4220 ( .C ( clk ), .D ( signal_9811 ), .Q ( signal_9812 ) ) ;
    buf_clk cell_4224 ( .C ( clk ), .D ( signal_9815 ), .Q ( signal_9816 ) ) ;
    buf_clk cell_4228 ( .C ( clk ), .D ( signal_9819 ), .Q ( signal_9820 ) ) ;
    buf_clk cell_4232 ( .C ( clk ), .D ( signal_9823 ), .Q ( signal_9824 ) ) ;
    buf_clk cell_4236 ( .C ( clk ), .D ( signal_9827 ), .Q ( signal_9828 ) ) ;
    buf_clk cell_4240 ( .C ( clk ), .D ( signal_9831 ), .Q ( signal_9832 ) ) ;
    buf_clk cell_4244 ( .C ( clk ), .D ( signal_9835 ), .Q ( signal_9836 ) ) ;
    buf_clk cell_4248 ( .C ( clk ), .D ( signal_9839 ), .Q ( signal_9840 ) ) ;
    buf_clk cell_4252 ( .C ( clk ), .D ( signal_9843 ), .Q ( signal_9844 ) ) ;
    buf_clk cell_4256 ( .C ( clk ), .D ( signal_9847 ), .Q ( signal_9848 ) ) ;
    buf_clk cell_4258 ( .C ( clk ), .D ( signal_9849 ), .Q ( signal_9850 ) ) ;
    buf_clk cell_4260 ( .C ( clk ), .D ( signal_9851 ), .Q ( signal_9852 ) ) ;
    buf_clk cell_4262 ( .C ( clk ), .D ( signal_9853 ), .Q ( signal_9854 ) ) ;
    buf_clk cell_4268 ( .C ( clk ), .D ( signal_9859 ), .Q ( signal_9860 ) ) ;
    buf_clk cell_4274 ( .C ( clk ), .D ( signal_9865 ), .Q ( signal_9866 ) ) ;
    buf_clk cell_4280 ( .C ( clk ), .D ( signal_9871 ), .Q ( signal_9872 ) ) ;
    buf_clk cell_4284 ( .C ( clk ), .D ( signal_9875 ), .Q ( signal_9876 ) ) ;
    buf_clk cell_4288 ( .C ( clk ), .D ( signal_9879 ), .Q ( signal_9880 ) ) ;
    buf_clk cell_4292 ( .C ( clk ), .D ( signal_9883 ), .Q ( signal_9884 ) ) ;
    buf_clk cell_4298 ( .C ( clk ), .D ( signal_9889 ), .Q ( signal_9890 ) ) ;
    buf_clk cell_4304 ( .C ( clk ), .D ( signal_9895 ), .Q ( signal_9896 ) ) ;
    buf_clk cell_4310 ( .C ( clk ), .D ( signal_9901 ), .Q ( signal_9902 ) ) ;
    buf_clk cell_4314 ( .C ( clk ), .D ( signal_9905 ), .Q ( signal_9906 ) ) ;
    buf_clk cell_4318 ( .C ( clk ), .D ( signal_9909 ), .Q ( signal_9910 ) ) ;
    buf_clk cell_4322 ( .C ( clk ), .D ( signal_9913 ), .Q ( signal_9914 ) ) ;
    buf_clk cell_4326 ( .C ( clk ), .D ( signal_9917 ), .Q ( signal_9918 ) ) ;
    buf_clk cell_4330 ( .C ( clk ), .D ( signal_9921 ), .Q ( signal_9922 ) ) ;
    buf_clk cell_4334 ( .C ( clk ), .D ( signal_9925 ), .Q ( signal_9926 ) ) ;
    buf_clk cell_4338 ( .C ( clk ), .D ( signal_9929 ), .Q ( signal_9930 ) ) ;
    buf_clk cell_4342 ( .C ( clk ), .D ( signal_9933 ), .Q ( signal_9934 ) ) ;
    buf_clk cell_4346 ( .C ( clk ), .D ( signal_9937 ), .Q ( signal_9938 ) ) ;
    buf_clk cell_4348 ( .C ( clk ), .D ( signal_9939 ), .Q ( signal_9940 ) ) ;
    buf_clk cell_4350 ( .C ( clk ), .D ( signal_9941 ), .Q ( signal_9942 ) ) ;
    buf_clk cell_4352 ( .C ( clk ), .D ( signal_9943 ), .Q ( signal_9944 ) ) ;
    buf_clk cell_4356 ( .C ( clk ), .D ( signal_9947 ), .Q ( signal_9948 ) ) ;
    buf_clk cell_4360 ( .C ( clk ), .D ( signal_9951 ), .Q ( signal_9952 ) ) ;
    buf_clk cell_4364 ( .C ( clk ), .D ( signal_9955 ), .Q ( signal_9956 ) ) ;
    buf_clk cell_4368 ( .C ( clk ), .D ( signal_9959 ), .Q ( signal_9960 ) ) ;
    buf_clk cell_4372 ( .C ( clk ), .D ( signal_9963 ), .Q ( signal_9964 ) ) ;
    buf_clk cell_4376 ( .C ( clk ), .D ( signal_9967 ), .Q ( signal_9968 ) ) ;
    buf_clk cell_4382 ( .C ( clk ), .D ( signal_9973 ), .Q ( signal_9974 ) ) ;
    buf_clk cell_4388 ( .C ( clk ), .D ( signal_9979 ), .Q ( signal_9980 ) ) ;
    buf_clk cell_4394 ( .C ( clk ), .D ( signal_9985 ), .Q ( signal_9986 ) ) ;
    buf_clk cell_4396 ( .C ( clk ), .D ( signal_9987 ), .Q ( signal_9988 ) ) ;
    buf_clk cell_4398 ( .C ( clk ), .D ( signal_9989 ), .Q ( signal_9990 ) ) ;
    buf_clk cell_4400 ( .C ( clk ), .D ( signal_9991 ), .Q ( signal_9992 ) ) ;
    buf_clk cell_4402 ( .C ( clk ), .D ( signal_9993 ), .Q ( signal_9994 ) ) ;
    buf_clk cell_4404 ( .C ( clk ), .D ( signal_9995 ), .Q ( signal_9996 ) ) ;
    buf_clk cell_4406 ( .C ( clk ), .D ( signal_9997 ), .Q ( signal_9998 ) ) ;
    buf_clk cell_4410 ( .C ( clk ), .D ( signal_10001 ), .Q ( signal_10002 ) ) ;
    buf_clk cell_4414 ( .C ( clk ), .D ( signal_10005 ), .Q ( signal_10006 ) ) ;
    buf_clk cell_4418 ( .C ( clk ), .D ( signal_10009 ), .Q ( signal_10010 ) ) ;
    buf_clk cell_4424 ( .C ( clk ), .D ( signal_10015 ), .Q ( signal_10016 ) ) ;
    buf_clk cell_4430 ( .C ( clk ), .D ( signal_10021 ), .Q ( signal_10022 ) ) ;
    buf_clk cell_4436 ( .C ( clk ), .D ( signal_10027 ), .Q ( signal_10028 ) ) ;
    buf_clk cell_4442 ( .C ( clk ), .D ( signal_10033 ), .Q ( signal_10034 ) ) ;
    buf_clk cell_4448 ( .C ( clk ), .D ( signal_10039 ), .Q ( signal_10040 ) ) ;
    buf_clk cell_4454 ( .C ( clk ), .D ( signal_10045 ), .Q ( signal_10046 ) ) ;
    buf_clk cell_4460 ( .C ( clk ), .D ( signal_10051 ), .Q ( signal_10052 ) ) ;
    buf_clk cell_4466 ( .C ( clk ), .D ( signal_10057 ), .Q ( signal_10058 ) ) ;
    buf_clk cell_4472 ( .C ( clk ), .D ( signal_10063 ), .Q ( signal_10064 ) ) ;
    buf_clk cell_4476 ( .C ( clk ), .D ( signal_10067 ), .Q ( signal_10068 ) ) ;
    buf_clk cell_4480 ( .C ( clk ), .D ( signal_10071 ), .Q ( signal_10072 ) ) ;
    buf_clk cell_4484 ( .C ( clk ), .D ( signal_10075 ), .Q ( signal_10076 ) ) ;
    buf_clk cell_4486 ( .C ( clk ), .D ( signal_10077 ), .Q ( signal_10078 ) ) ;
    buf_clk cell_4488 ( .C ( clk ), .D ( signal_10079 ), .Q ( signal_10080 ) ) ;
    buf_clk cell_4490 ( .C ( clk ), .D ( signal_10081 ), .Q ( signal_10082 ) ) ;
    buf_clk cell_4492 ( .C ( clk ), .D ( signal_10083 ), .Q ( signal_10084 ) ) ;
    buf_clk cell_4494 ( .C ( clk ), .D ( signal_10085 ), .Q ( signal_10086 ) ) ;
    buf_clk cell_4496 ( .C ( clk ), .D ( signal_10087 ), .Q ( signal_10088 ) ) ;
    buf_clk cell_4502 ( .C ( clk ), .D ( signal_10093 ), .Q ( signal_10094 ) ) ;
    buf_clk cell_4510 ( .C ( clk ), .D ( signal_10101 ), .Q ( signal_10102 ) ) ;
    buf_clk cell_4518 ( .C ( clk ), .D ( signal_10109 ), .Q ( signal_10110 ) ) ;
    buf_clk cell_4522 ( .C ( clk ), .D ( signal_10113 ), .Q ( signal_10114 ) ) ;
    buf_clk cell_4526 ( .C ( clk ), .D ( signal_10117 ), .Q ( signal_10118 ) ) ;
    buf_clk cell_4530 ( .C ( clk ), .D ( signal_10121 ), .Q ( signal_10122 ) ) ;
    buf_clk cell_4536 ( .C ( clk ), .D ( signal_10127 ), .Q ( signal_10128 ) ) ;
    buf_clk cell_4542 ( .C ( clk ), .D ( signal_10133 ), .Q ( signal_10134 ) ) ;
    buf_clk cell_4548 ( .C ( clk ), .D ( signal_10139 ), .Q ( signal_10140 ) ) ;
    buf_clk cell_4554 ( .C ( clk ), .D ( signal_10145 ), .Q ( signal_10146 ) ) ;
    buf_clk cell_4560 ( .C ( clk ), .D ( signal_10151 ), .Q ( signal_10152 ) ) ;
    buf_clk cell_4566 ( .C ( clk ), .D ( signal_10157 ), .Q ( signal_10158 ) ) ;
    buf_clk cell_4570 ( .C ( clk ), .D ( signal_10161 ), .Q ( signal_10162 ) ) ;
    buf_clk cell_4574 ( .C ( clk ), .D ( signal_10165 ), .Q ( signal_10166 ) ) ;
    buf_clk cell_4578 ( .C ( clk ), .D ( signal_10169 ), .Q ( signal_10170 ) ) ;
    buf_clk cell_4584 ( .C ( clk ), .D ( signal_10175 ), .Q ( signal_10176 ) ) ;
    buf_clk cell_4590 ( .C ( clk ), .D ( signal_10181 ), .Q ( signal_10182 ) ) ;
    buf_clk cell_4596 ( .C ( clk ), .D ( signal_10187 ), .Q ( signal_10188 ) ) ;
    buf_clk cell_4600 ( .C ( clk ), .D ( signal_10191 ), .Q ( signal_10192 ) ) ;
    buf_clk cell_4604 ( .C ( clk ), .D ( signal_10195 ), .Q ( signal_10196 ) ) ;
    buf_clk cell_4608 ( .C ( clk ), .D ( signal_10199 ), .Q ( signal_10200 ) ) ;
    buf_clk cell_4612 ( .C ( clk ), .D ( signal_10203 ), .Q ( signal_10204 ) ) ;
    buf_clk cell_4616 ( .C ( clk ), .D ( signal_10207 ), .Q ( signal_10208 ) ) ;
    buf_clk cell_4620 ( .C ( clk ), .D ( signal_10211 ), .Q ( signal_10212 ) ) ;
    buf_clk cell_4638 ( .C ( clk ), .D ( signal_10229 ), .Q ( signal_10230 ) ) ;
    buf_clk cell_4644 ( .C ( clk ), .D ( signal_10235 ), .Q ( signal_10236 ) ) ;
    buf_clk cell_4650 ( .C ( clk ), .D ( signal_10241 ), .Q ( signal_10242 ) ) ;
    buf_clk cell_4656 ( .C ( clk ), .D ( signal_10247 ), .Q ( signal_10248 ) ) ;
    buf_clk cell_4662 ( .C ( clk ), .D ( signal_10253 ), .Q ( signal_10254 ) ) ;
    buf_clk cell_4668 ( .C ( clk ), .D ( signal_10259 ), .Q ( signal_10260 ) ) ;
    buf_clk cell_4674 ( .C ( clk ), .D ( signal_10265 ), .Q ( signal_10266 ) ) ;
    buf_clk cell_4680 ( .C ( clk ), .D ( signal_10271 ), .Q ( signal_10272 ) ) ;
    buf_clk cell_4686 ( .C ( clk ), .D ( signal_10277 ), .Q ( signal_10278 ) ) ;
    buf_clk cell_4696 ( .C ( clk ), .D ( signal_10287 ), .Q ( signal_10288 ) ) ;
    buf_clk cell_4700 ( .C ( clk ), .D ( signal_10291 ), .Q ( signal_10292 ) ) ;
    buf_clk cell_4704 ( .C ( clk ), .D ( signal_10295 ), .Q ( signal_10296 ) ) ;
    buf_clk cell_4710 ( .C ( clk ), .D ( signal_10301 ), .Q ( signal_10302 ) ) ;
    buf_clk cell_4716 ( .C ( clk ), .D ( signal_10307 ), .Q ( signal_10308 ) ) ;
    buf_clk cell_4722 ( .C ( clk ), .D ( signal_10313 ), .Q ( signal_10314 ) ) ;
    buf_clk cell_4734 ( .C ( clk ), .D ( signal_10325 ), .Q ( signal_10326 ) ) ;
    buf_clk cell_4740 ( .C ( clk ), .D ( signal_10331 ), .Q ( signal_10332 ) ) ;
    buf_clk cell_4746 ( .C ( clk ), .D ( signal_10337 ), .Q ( signal_10338 ) ) ;
    buf_clk cell_4760 ( .C ( clk ), .D ( signal_10351 ), .Q ( signal_10352 ) ) ;
    buf_clk cell_4768 ( .C ( clk ), .D ( signal_10359 ), .Q ( signal_10360 ) ) ;
    buf_clk cell_4776 ( .C ( clk ), .D ( signal_10367 ), .Q ( signal_10368 ) ) ;
    buf_clk cell_4780 ( .C ( clk ), .D ( signal_10371 ), .Q ( signal_10372 ) ) ;
    buf_clk cell_4784 ( .C ( clk ), .D ( signal_10375 ), .Q ( signal_10376 ) ) ;
    buf_clk cell_4788 ( .C ( clk ), .D ( signal_10379 ), .Q ( signal_10380 ) ) ;
    buf_clk cell_4792 ( .C ( clk ), .D ( signal_10383 ), .Q ( signal_10384 ) ) ;
    buf_clk cell_4796 ( .C ( clk ), .D ( signal_10387 ), .Q ( signal_10388 ) ) ;
    buf_clk cell_4800 ( .C ( clk ), .D ( signal_10391 ), .Q ( signal_10392 ) ) ;
    buf_clk cell_4806 ( .C ( clk ), .D ( signal_10397 ), .Q ( signal_10398 ) ) ;
    buf_clk cell_4812 ( .C ( clk ), .D ( signal_10403 ), .Q ( signal_10404 ) ) ;
    buf_clk cell_4818 ( .C ( clk ), .D ( signal_10409 ), .Q ( signal_10410 ) ) ;
    buf_clk cell_4824 ( .C ( clk ), .D ( signal_10415 ), .Q ( signal_10416 ) ) ;
    buf_clk cell_4830 ( .C ( clk ), .D ( signal_10421 ), .Q ( signal_10422 ) ) ;
    buf_clk cell_4836 ( .C ( clk ), .D ( signal_10427 ), .Q ( signal_10428 ) ) ;
    buf_clk cell_4840 ( .C ( clk ), .D ( signal_10431 ), .Q ( signal_10432 ) ) ;
    buf_clk cell_4844 ( .C ( clk ), .D ( signal_10435 ), .Q ( signal_10436 ) ) ;
    buf_clk cell_4848 ( .C ( clk ), .D ( signal_10439 ), .Q ( signal_10440 ) ) ;
    buf_clk cell_4856 ( .C ( clk ), .D ( signal_10447 ), .Q ( signal_10448 ) ) ;
    buf_clk cell_4864 ( .C ( clk ), .D ( signal_10455 ), .Q ( signal_10456 ) ) ;
    buf_clk cell_4872 ( .C ( clk ), .D ( signal_10463 ), .Q ( signal_10464 ) ) ;
    buf_clk cell_4878 ( .C ( clk ), .D ( signal_10469 ), .Q ( signal_10470 ) ) ;
    buf_clk cell_4884 ( .C ( clk ), .D ( signal_10475 ), .Q ( signal_10476 ) ) ;
    buf_clk cell_4890 ( .C ( clk ), .D ( signal_10481 ), .Q ( signal_10482 ) ) ;
    buf_clk cell_4896 ( .C ( clk ), .D ( signal_10487 ), .Q ( signal_10488 ) ) ;
    buf_clk cell_4902 ( .C ( clk ), .D ( signal_10493 ), .Q ( signal_10494 ) ) ;
    buf_clk cell_4908 ( .C ( clk ), .D ( signal_10499 ), .Q ( signal_10500 ) ) ;
    buf_clk cell_4926 ( .C ( clk ), .D ( signal_10517 ), .Q ( signal_10518 ) ) ;
    buf_clk cell_4932 ( .C ( clk ), .D ( signal_10523 ), .Q ( signal_10524 ) ) ;
    buf_clk cell_4938 ( .C ( clk ), .D ( signal_10529 ), .Q ( signal_10530 ) ) ;
    buf_clk cell_4956 ( .C ( clk ), .D ( signal_10547 ), .Q ( signal_10548 ) ) ;
    buf_clk cell_4962 ( .C ( clk ), .D ( signal_10553 ), .Q ( signal_10554 ) ) ;
    buf_clk cell_4968 ( .C ( clk ), .D ( signal_10559 ), .Q ( signal_10560 ) ) ;
    buf_clk cell_4974 ( .C ( clk ), .D ( signal_10565 ), .Q ( signal_10566 ) ) ;
    buf_clk cell_4980 ( .C ( clk ), .D ( signal_10571 ), .Q ( signal_10572 ) ) ;
    buf_clk cell_4986 ( .C ( clk ), .D ( signal_10577 ), .Q ( signal_10578 ) ) ;
    buf_clk cell_4990 ( .C ( clk ), .D ( signal_10581 ), .Q ( signal_10582 ) ) ;
    buf_clk cell_4994 ( .C ( clk ), .D ( signal_10585 ), .Q ( signal_10586 ) ) ;
    buf_clk cell_4998 ( .C ( clk ), .D ( signal_10589 ), .Q ( signal_10590 ) ) ;
    buf_clk cell_5006 ( .C ( clk ), .D ( signal_10597 ), .Q ( signal_10598 ) ) ;
    buf_clk cell_5016 ( .C ( clk ), .D ( signal_10607 ), .Q ( signal_10608 ) ) ;
    buf_clk cell_5026 ( .C ( clk ), .D ( signal_10617 ), .Q ( signal_10618 ) ) ;
    buf_clk cell_5032 ( .C ( clk ), .D ( signal_10623 ), .Q ( signal_10624 ) ) ;
    buf_clk cell_5038 ( .C ( clk ), .D ( signal_10629 ), .Q ( signal_10630 ) ) ;
    buf_clk cell_5044 ( .C ( clk ), .D ( signal_10635 ), .Q ( signal_10636 ) ) ;
    buf_clk cell_5052 ( .C ( clk ), .D ( signal_10643 ), .Q ( signal_10644 ) ) ;
    buf_clk cell_5060 ( .C ( clk ), .D ( signal_10651 ), .Q ( signal_10652 ) ) ;
    buf_clk cell_5068 ( .C ( clk ), .D ( signal_10659 ), .Q ( signal_10660 ) ) ;
    buf_clk cell_5076 ( .C ( clk ), .D ( signal_10667 ), .Q ( signal_10668 ) ) ;
    buf_clk cell_5084 ( .C ( clk ), .D ( signal_10675 ), .Q ( signal_10676 ) ) ;
    buf_clk cell_5092 ( .C ( clk ), .D ( signal_10683 ), .Q ( signal_10684 ) ) ;
    buf_clk cell_5150 ( .C ( clk ), .D ( signal_10741 ), .Q ( signal_10742 ) ) ;
    buf_clk cell_5160 ( .C ( clk ), .D ( signal_10751 ), .Q ( signal_10752 ) ) ;
    buf_clk cell_5170 ( .C ( clk ), .D ( signal_10761 ), .Q ( signal_10762 ) ) ;
    buf_clk cell_5176 ( .C ( clk ), .D ( signal_10767 ), .Q ( signal_10768 ) ) ;
    buf_clk cell_5182 ( .C ( clk ), .D ( signal_10773 ), .Q ( signal_10774 ) ) ;
    buf_clk cell_5188 ( .C ( clk ), .D ( signal_10779 ), .Q ( signal_10780 ) ) ;
    buf_clk cell_5202 ( .C ( clk ), .D ( signal_10793 ), .Q ( signal_10794 ) ) ;
    buf_clk cell_5210 ( .C ( clk ), .D ( signal_10801 ), .Q ( signal_10802 ) ) ;
    buf_clk cell_5218 ( .C ( clk ), .D ( signal_10809 ), .Q ( signal_10810 ) ) ;
    buf_clk cell_5224 ( .C ( clk ), .D ( signal_10815 ), .Q ( signal_10816 ) ) ;
    buf_clk cell_5230 ( .C ( clk ), .D ( signal_10821 ), .Q ( signal_10822 ) ) ;
    buf_clk cell_5236 ( .C ( clk ), .D ( signal_10827 ), .Q ( signal_10828 ) ) ;
    buf_clk cell_5244 ( .C ( clk ), .D ( signal_10835 ), .Q ( signal_10836 ) ) ;
    buf_clk cell_5252 ( .C ( clk ), .D ( signal_10843 ), .Q ( signal_10844 ) ) ;
    buf_clk cell_5260 ( .C ( clk ), .D ( signal_10851 ), .Q ( signal_10852 ) ) ;
    buf_clk cell_5268 ( .C ( clk ), .D ( signal_10859 ), .Q ( signal_10860 ) ) ;
    buf_clk cell_5276 ( .C ( clk ), .D ( signal_10867 ), .Q ( signal_10868 ) ) ;
    buf_clk cell_5284 ( .C ( clk ), .D ( signal_10875 ), .Q ( signal_10876 ) ) ;
    buf_clk cell_5292 ( .C ( clk ), .D ( signal_10883 ), .Q ( signal_10884 ) ) ;
    buf_clk cell_5300 ( .C ( clk ), .D ( signal_10891 ), .Q ( signal_10892 ) ) ;
    buf_clk cell_5308 ( .C ( clk ), .D ( signal_10899 ), .Q ( signal_10900 ) ) ;
    buf_clk cell_5318 ( .C ( clk ), .D ( signal_10909 ), .Q ( signal_10910 ) ) ;
    buf_clk cell_5328 ( .C ( clk ), .D ( signal_10919 ), .Q ( signal_10920 ) ) ;
    buf_clk cell_5338 ( .C ( clk ), .D ( signal_10929 ), .Q ( signal_10930 ) ) ;
    buf_clk cell_5346 ( .C ( clk ), .D ( signal_10937 ), .Q ( signal_10938 ) ) ;
    buf_clk cell_5354 ( .C ( clk ), .D ( signal_10945 ), .Q ( signal_10946 ) ) ;
    buf_clk cell_5362 ( .C ( clk ), .D ( signal_10953 ), .Q ( signal_10954 ) ) ;
    buf_clk cell_5370 ( .C ( clk ), .D ( signal_10961 ), .Q ( signal_10962 ) ) ;
    buf_clk cell_5378 ( .C ( clk ), .D ( signal_10969 ), .Q ( signal_10970 ) ) ;
    buf_clk cell_5386 ( .C ( clk ), .D ( signal_10977 ), .Q ( signal_10978 ) ) ;
    buf_clk cell_5400 ( .C ( clk ), .D ( signal_10991 ), .Q ( signal_10992 ) ) ;
    buf_clk cell_5408 ( .C ( clk ), .D ( signal_10999 ), .Q ( signal_11000 ) ) ;
    buf_clk cell_5416 ( .C ( clk ), .D ( signal_11007 ), .Q ( signal_11008 ) ) ;
    buf_clk cell_5424 ( .C ( clk ), .D ( signal_11015 ), .Q ( signal_11016 ) ) ;
    buf_clk cell_5432 ( .C ( clk ), .D ( signal_11023 ), .Q ( signal_11024 ) ) ;
    buf_clk cell_5440 ( .C ( clk ), .D ( signal_11031 ), .Q ( signal_11032 ) ) ;
    buf_clk cell_5448 ( .C ( clk ), .D ( signal_11039 ), .Q ( signal_11040 ) ) ;
    buf_clk cell_5456 ( .C ( clk ), .D ( signal_11047 ), .Q ( signal_11048 ) ) ;
    buf_clk cell_5464 ( .C ( clk ), .D ( signal_11055 ), .Q ( signal_11056 ) ) ;
    buf_clk cell_5488 ( .C ( clk ), .D ( signal_11079 ), .Q ( signal_11080 ) ) ;
    buf_clk cell_5496 ( .C ( clk ), .D ( signal_11087 ), .Q ( signal_11088 ) ) ;
    buf_clk cell_5504 ( .C ( clk ), .D ( signal_11095 ), .Q ( signal_11096 ) ) ;
    buf_clk cell_5548 ( .C ( clk ), .D ( signal_11139 ), .Q ( signal_11140 ) ) ;
    buf_clk cell_5556 ( .C ( clk ), .D ( signal_11147 ), .Q ( signal_11148 ) ) ;
    buf_clk cell_5564 ( .C ( clk ), .D ( signal_11155 ), .Q ( signal_11156 ) ) ;
    buf_clk cell_5574 ( .C ( clk ), .D ( signal_11165 ), .Q ( signal_11166 ) ) ;
    buf_clk cell_5584 ( .C ( clk ), .D ( signal_11175 ), .Q ( signal_11176 ) ) ;
    buf_clk cell_5594 ( .C ( clk ), .D ( signal_11185 ), .Q ( signal_11186 ) ) ;
    buf_clk cell_5626 ( .C ( clk ), .D ( signal_11217 ), .Q ( signal_11218 ) ) ;
    buf_clk cell_5634 ( .C ( clk ), .D ( signal_11225 ), .Q ( signal_11226 ) ) ;
    buf_clk cell_5642 ( .C ( clk ), .D ( signal_11233 ), .Q ( signal_11234 ) ) ;
    buf_clk cell_5652 ( .C ( clk ), .D ( signal_11243 ), .Q ( signal_11244 ) ) ;
    buf_clk cell_5662 ( .C ( clk ), .D ( signal_11253 ), .Q ( signal_11254 ) ) ;
    buf_clk cell_5672 ( .C ( clk ), .D ( signal_11263 ), .Q ( signal_11264 ) ) ;
    buf_clk cell_5680 ( .C ( clk ), .D ( signal_11271 ), .Q ( signal_11272 ) ) ;
    buf_clk cell_5688 ( .C ( clk ), .D ( signal_11279 ), .Q ( signal_11280 ) ) ;
    buf_clk cell_5696 ( .C ( clk ), .D ( signal_11287 ), .Q ( signal_11288 ) ) ;
    buf_clk cell_5920 ( .C ( clk ), .D ( signal_11511 ), .Q ( signal_11512 ) ) ;
    buf_clk cell_5930 ( .C ( clk ), .D ( signal_11521 ), .Q ( signal_11522 ) ) ;
    buf_clk cell_5940 ( .C ( clk ), .D ( signal_11531 ), .Q ( signal_11532 ) ) ;
    buf_clk cell_6184 ( .C ( clk ), .D ( signal_11775 ), .Q ( signal_11776 ) ) ;
    buf_clk cell_6196 ( .C ( clk ), .D ( signal_11787 ), .Q ( signal_11788 ) ) ;
    buf_clk cell_6208 ( .C ( clk ), .D ( signal_11799 ), .Q ( signal_11800 ) ) ;
    buf_clk cell_6258 ( .C ( clk ), .D ( signal_11849 ), .Q ( signal_11850 ) ) ;
    buf_clk cell_6272 ( .C ( clk ), .D ( signal_11863 ), .Q ( signal_11864 ) ) ;
    buf_clk cell_6286 ( .C ( clk ), .D ( signal_11877 ), .Q ( signal_11878 ) ) ;
    buf_clk cell_6324 ( .C ( clk ), .D ( signal_11915 ), .Q ( signal_11916 ) ) ;
    buf_clk cell_6338 ( .C ( clk ), .D ( signal_11929 ), .Q ( signal_11930 ) ) ;
    buf_clk cell_6352 ( .C ( clk ), .D ( signal_11943 ), .Q ( signal_11944 ) ) ;
    buf_clk cell_6444 ( .C ( clk ), .D ( signal_12035 ), .Q ( signal_12036 ) ) ;
    buf_clk cell_6460 ( .C ( clk ), .D ( signal_12051 ), .Q ( signal_12052 ) ) ;
    buf_clk cell_6476 ( .C ( clk ), .D ( signal_12067 ), .Q ( signal_12068 ) ) ;
    buf_clk cell_6504 ( .C ( clk ), .D ( signal_12095 ), .Q ( signal_12096 ) ) ;
    buf_clk cell_6520 ( .C ( clk ), .D ( signal_12111 ), .Q ( signal_12112 ) ) ;
    buf_clk cell_6536 ( .C ( clk ), .D ( signal_12127 ), .Q ( signal_12128 ) ) ;
    buf_clk cell_6688 ( .C ( clk ), .D ( signal_12279 ), .Q ( signal_12280 ) ) ;
    buf_clk cell_6704 ( .C ( clk ), .D ( signal_12295 ), .Q ( signal_12296 ) ) ;
    buf_clk cell_6720 ( .C ( clk ), .D ( signal_12311 ), .Q ( signal_12312 ) ) ;
    buf_clk cell_6738 ( .C ( clk ), .D ( signal_12329 ), .Q ( signal_12330 ) ) ;
    buf_clk cell_6756 ( .C ( clk ), .D ( signal_12347 ), .Q ( signal_12348 ) ) ;
    buf_clk cell_6774 ( .C ( clk ), .D ( signal_12365 ), .Q ( signal_12366 ) ) ;
    buf_clk cell_6888 ( .C ( clk ), .D ( signal_12479 ), .Q ( signal_12480 ) ) ;
    buf_clk cell_6908 ( .C ( clk ), .D ( signal_12499 ), .Q ( signal_12500 ) ) ;
    buf_clk cell_6928 ( .C ( clk ), .D ( signal_12519 ), .Q ( signal_12520 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_4503 ( .C ( clk ), .D ( signal_10094 ), .Q ( signal_10095 ) ) ;
    buf_clk cell_4511 ( .C ( clk ), .D ( signal_10102 ), .Q ( signal_10103 ) ) ;
    buf_clk cell_4519 ( .C ( clk ), .D ( signal_10110 ), .Q ( signal_10111 ) ) ;
    buf_clk cell_4523 ( .C ( clk ), .D ( signal_10114 ), .Q ( signal_10115 ) ) ;
    buf_clk cell_4527 ( .C ( clk ), .D ( signal_10118 ), .Q ( signal_10119 ) ) ;
    buf_clk cell_4531 ( .C ( clk ), .D ( signal_10122 ), .Q ( signal_10123 ) ) ;
    buf_clk cell_4537 ( .C ( clk ), .D ( signal_10128 ), .Q ( signal_10129 ) ) ;
    buf_clk cell_4543 ( .C ( clk ), .D ( signal_10134 ), .Q ( signal_10135 ) ) ;
    buf_clk cell_4549 ( .C ( clk ), .D ( signal_10140 ), .Q ( signal_10141 ) ) ;
    buf_clk cell_4555 ( .C ( clk ), .D ( signal_10146 ), .Q ( signal_10147 ) ) ;
    buf_clk cell_4561 ( .C ( clk ), .D ( signal_10152 ), .Q ( signal_10153 ) ) ;
    buf_clk cell_4567 ( .C ( clk ), .D ( signal_10158 ), .Q ( signal_10159 ) ) ;
    buf_clk cell_4571 ( .C ( clk ), .D ( signal_10162 ), .Q ( signal_10163 ) ) ;
    buf_clk cell_4575 ( .C ( clk ), .D ( signal_10166 ), .Q ( signal_10167 ) ) ;
    buf_clk cell_4579 ( .C ( clk ), .D ( signal_10170 ), .Q ( signal_10171 ) ) ;
    buf_clk cell_4585 ( .C ( clk ), .D ( signal_10176 ), .Q ( signal_10177 ) ) ;
    buf_clk cell_4591 ( .C ( clk ), .D ( signal_10182 ), .Q ( signal_10183 ) ) ;
    buf_clk cell_4597 ( .C ( clk ), .D ( signal_10188 ), .Q ( signal_10189 ) ) ;
    buf_clk cell_4601 ( .C ( clk ), .D ( signal_10192 ), .Q ( signal_10193 ) ) ;
    buf_clk cell_4605 ( .C ( clk ), .D ( signal_10196 ), .Q ( signal_10197 ) ) ;
    buf_clk cell_4609 ( .C ( clk ), .D ( signal_10200 ), .Q ( signal_10201 ) ) ;
    buf_clk cell_4613 ( .C ( clk ), .D ( signal_10204 ), .Q ( signal_10205 ) ) ;
    buf_clk cell_4617 ( .C ( clk ), .D ( signal_10208 ), .Q ( signal_10209 ) ) ;
    buf_clk cell_4621 ( .C ( clk ), .D ( signal_10212 ), .Q ( signal_10213 ) ) ;
    buf_clk cell_4623 ( .C ( clk ), .D ( signal_2071 ), .Q ( signal_10215 ) ) ;
    buf_clk cell_4625 ( .C ( clk ), .D ( signal_4666 ), .Q ( signal_10217 ) ) ;
    buf_clk cell_4627 ( .C ( clk ), .D ( signal_4667 ), .Q ( signal_10219 ) ) ;
    buf_clk cell_4629 ( .C ( clk ), .D ( signal_9850 ), .Q ( signal_10221 ) ) ;
    buf_clk cell_4631 ( .C ( clk ), .D ( signal_9852 ), .Q ( signal_10223 ) ) ;
    buf_clk cell_4633 ( .C ( clk ), .D ( signal_9854 ), .Q ( signal_10225 ) ) ;
    buf_clk cell_4639 ( .C ( clk ), .D ( signal_10230 ), .Q ( signal_10231 ) ) ;
    buf_clk cell_4645 ( .C ( clk ), .D ( signal_10236 ), .Q ( signal_10237 ) ) ;
    buf_clk cell_4651 ( .C ( clk ), .D ( signal_10242 ), .Q ( signal_10243 ) ) ;
    buf_clk cell_4657 ( .C ( clk ), .D ( signal_10248 ), .Q ( signal_10249 ) ) ;
    buf_clk cell_4663 ( .C ( clk ), .D ( signal_10254 ), .Q ( signal_10255 ) ) ;
    buf_clk cell_4669 ( .C ( clk ), .D ( signal_10260 ), .Q ( signal_10261 ) ) ;
    buf_clk cell_4675 ( .C ( clk ), .D ( signal_10266 ), .Q ( signal_10267 ) ) ;
    buf_clk cell_4681 ( .C ( clk ), .D ( signal_10272 ), .Q ( signal_10273 ) ) ;
    buf_clk cell_4687 ( .C ( clk ), .D ( signal_10278 ), .Q ( signal_10279 ) ) ;
    buf_clk cell_4689 ( .C ( clk ), .D ( signal_9654 ), .Q ( signal_10281 ) ) ;
    buf_clk cell_4691 ( .C ( clk ), .D ( signal_9658 ), .Q ( signal_10283 ) ) ;
    buf_clk cell_4693 ( .C ( clk ), .D ( signal_9662 ), .Q ( signal_10285 ) ) ;
    buf_clk cell_4697 ( .C ( clk ), .D ( signal_10288 ), .Q ( signal_10289 ) ) ;
    buf_clk cell_4701 ( .C ( clk ), .D ( signal_10292 ), .Q ( signal_10293 ) ) ;
    buf_clk cell_4705 ( .C ( clk ), .D ( signal_10296 ), .Q ( signal_10297 ) ) ;
    buf_clk cell_4711 ( .C ( clk ), .D ( signal_10302 ), .Q ( signal_10303 ) ) ;
    buf_clk cell_4717 ( .C ( clk ), .D ( signal_10308 ), .Q ( signal_10309 ) ) ;
    buf_clk cell_4723 ( .C ( clk ), .D ( signal_10314 ), .Q ( signal_10315 ) ) ;
    buf_clk cell_4725 ( .C ( clk ), .D ( signal_2081 ), .Q ( signal_10317 ) ) ;
    buf_clk cell_4727 ( .C ( clk ), .D ( signal_4686 ), .Q ( signal_10319 ) ) ;
    buf_clk cell_4729 ( .C ( clk ), .D ( signal_4687 ), .Q ( signal_10321 ) ) ;
    buf_clk cell_4735 ( .C ( clk ), .D ( signal_10326 ), .Q ( signal_10327 ) ) ;
    buf_clk cell_4741 ( .C ( clk ), .D ( signal_10332 ), .Q ( signal_10333 ) ) ;
    buf_clk cell_4747 ( .C ( clk ), .D ( signal_10338 ), .Q ( signal_10339 ) ) ;
    buf_clk cell_4749 ( .C ( clk ), .D ( signal_2069 ), .Q ( signal_10341 ) ) ;
    buf_clk cell_4751 ( .C ( clk ), .D ( signal_4662 ), .Q ( signal_10343 ) ) ;
    buf_clk cell_4753 ( .C ( clk ), .D ( signal_4663 ), .Q ( signal_10345 ) ) ;
    buf_clk cell_4761 ( .C ( clk ), .D ( signal_10352 ), .Q ( signal_10353 ) ) ;
    buf_clk cell_4769 ( .C ( clk ), .D ( signal_10360 ), .Q ( signal_10361 ) ) ;
    buf_clk cell_4777 ( .C ( clk ), .D ( signal_10368 ), .Q ( signal_10369 ) ) ;
    buf_clk cell_4781 ( .C ( clk ), .D ( signal_10372 ), .Q ( signal_10373 ) ) ;
    buf_clk cell_4785 ( .C ( clk ), .D ( signal_10376 ), .Q ( signal_10377 ) ) ;
    buf_clk cell_4789 ( .C ( clk ), .D ( signal_10380 ), .Q ( signal_10381 ) ) ;
    buf_clk cell_4793 ( .C ( clk ), .D ( signal_10384 ), .Q ( signal_10385 ) ) ;
    buf_clk cell_4797 ( .C ( clk ), .D ( signal_10388 ), .Q ( signal_10389 ) ) ;
    buf_clk cell_4801 ( .C ( clk ), .D ( signal_10392 ), .Q ( signal_10393 ) ) ;
    buf_clk cell_4807 ( .C ( clk ), .D ( signal_10398 ), .Q ( signal_10399 ) ) ;
    buf_clk cell_4813 ( .C ( clk ), .D ( signal_10404 ), .Q ( signal_10405 ) ) ;
    buf_clk cell_4819 ( .C ( clk ), .D ( signal_10410 ), .Q ( signal_10411 ) ) ;
    buf_clk cell_4825 ( .C ( clk ), .D ( signal_10416 ), .Q ( signal_10417 ) ) ;
    buf_clk cell_4831 ( .C ( clk ), .D ( signal_10422 ), .Q ( signal_10423 ) ) ;
    buf_clk cell_4837 ( .C ( clk ), .D ( signal_10428 ), .Q ( signal_10429 ) ) ;
    buf_clk cell_4841 ( .C ( clk ), .D ( signal_10432 ), .Q ( signal_10433 ) ) ;
    buf_clk cell_4845 ( .C ( clk ), .D ( signal_10436 ), .Q ( signal_10437 ) ) ;
    buf_clk cell_4849 ( .C ( clk ), .D ( signal_10440 ), .Q ( signal_10441 ) ) ;
    buf_clk cell_4857 ( .C ( clk ), .D ( signal_10448 ), .Q ( signal_10449 ) ) ;
    buf_clk cell_4865 ( .C ( clk ), .D ( signal_10456 ), .Q ( signal_10457 ) ) ;
    buf_clk cell_4873 ( .C ( clk ), .D ( signal_10464 ), .Q ( signal_10465 ) ) ;
    buf_clk cell_4879 ( .C ( clk ), .D ( signal_10470 ), .Q ( signal_10471 ) ) ;
    buf_clk cell_4885 ( .C ( clk ), .D ( signal_10476 ), .Q ( signal_10477 ) ) ;
    buf_clk cell_4891 ( .C ( clk ), .D ( signal_10482 ), .Q ( signal_10483 ) ) ;
    buf_clk cell_4897 ( .C ( clk ), .D ( signal_10488 ), .Q ( signal_10489 ) ) ;
    buf_clk cell_4903 ( .C ( clk ), .D ( signal_10494 ), .Q ( signal_10495 ) ) ;
    buf_clk cell_4909 ( .C ( clk ), .D ( signal_10500 ), .Q ( signal_10501 ) ) ;
    buf_clk cell_4911 ( .C ( clk ), .D ( signal_2201 ), .Q ( signal_10503 ) ) ;
    buf_clk cell_4913 ( .C ( clk ), .D ( signal_4926 ), .Q ( signal_10505 ) ) ;
    buf_clk cell_4915 ( .C ( clk ), .D ( signal_4927 ), .Q ( signal_10507 ) ) ;
    buf_clk cell_4917 ( .C ( clk ), .D ( signal_9766 ), .Q ( signal_10509 ) ) ;
    buf_clk cell_4919 ( .C ( clk ), .D ( signal_9768 ), .Q ( signal_10511 ) ) ;
    buf_clk cell_4921 ( .C ( clk ), .D ( signal_9770 ), .Q ( signal_10513 ) ) ;
    buf_clk cell_4927 ( .C ( clk ), .D ( signal_10518 ), .Q ( signal_10519 ) ) ;
    buf_clk cell_4933 ( .C ( clk ), .D ( signal_10524 ), .Q ( signal_10525 ) ) ;
    buf_clk cell_4939 ( .C ( clk ), .D ( signal_10530 ), .Q ( signal_10531 ) ) ;
    buf_clk cell_4941 ( .C ( clk ), .D ( signal_9760 ), .Q ( signal_10533 ) ) ;
    buf_clk cell_4943 ( .C ( clk ), .D ( signal_9762 ), .Q ( signal_10535 ) ) ;
    buf_clk cell_4945 ( .C ( clk ), .D ( signal_9764 ), .Q ( signal_10537 ) ) ;
    buf_clk cell_4947 ( .C ( clk ), .D ( signal_9494 ), .Q ( signal_10539 ) ) ;
    buf_clk cell_4949 ( .C ( clk ), .D ( signal_9500 ), .Q ( signal_10541 ) ) ;
    buf_clk cell_4951 ( .C ( clk ), .D ( signal_9506 ), .Q ( signal_10543 ) ) ;
    buf_clk cell_4957 ( .C ( clk ), .D ( signal_10548 ), .Q ( signal_10549 ) ) ;
    buf_clk cell_4963 ( .C ( clk ), .D ( signal_10554 ), .Q ( signal_10555 ) ) ;
    buf_clk cell_4969 ( .C ( clk ), .D ( signal_10560 ), .Q ( signal_10561 ) ) ;
    buf_clk cell_4975 ( .C ( clk ), .D ( signal_10566 ), .Q ( signal_10567 ) ) ;
    buf_clk cell_4981 ( .C ( clk ), .D ( signal_10572 ), .Q ( signal_10573 ) ) ;
    buf_clk cell_4987 ( .C ( clk ), .D ( signal_10578 ), .Q ( signal_10579 ) ) ;
    buf_clk cell_4991 ( .C ( clk ), .D ( signal_10582 ), .Q ( signal_10583 ) ) ;
    buf_clk cell_4995 ( .C ( clk ), .D ( signal_10586 ), .Q ( signal_10587 ) ) ;
    buf_clk cell_4999 ( .C ( clk ), .D ( signal_10590 ), .Q ( signal_10591 ) ) ;
    buf_clk cell_5007 ( .C ( clk ), .D ( signal_10598 ), .Q ( signal_10599 ) ) ;
    buf_clk cell_5017 ( .C ( clk ), .D ( signal_10608 ), .Q ( signal_10609 ) ) ;
    buf_clk cell_5027 ( .C ( clk ), .D ( signal_10618 ), .Q ( signal_10619 ) ) ;
    buf_clk cell_5033 ( .C ( clk ), .D ( signal_10624 ), .Q ( signal_10625 ) ) ;
    buf_clk cell_5039 ( .C ( clk ), .D ( signal_10630 ), .Q ( signal_10631 ) ) ;
    buf_clk cell_5045 ( .C ( clk ), .D ( signal_10636 ), .Q ( signal_10637 ) ) ;
    buf_clk cell_5053 ( .C ( clk ), .D ( signal_10644 ), .Q ( signal_10645 ) ) ;
    buf_clk cell_5061 ( .C ( clk ), .D ( signal_10652 ), .Q ( signal_10653 ) ) ;
    buf_clk cell_5069 ( .C ( clk ), .D ( signal_10660 ), .Q ( signal_10661 ) ) ;
    buf_clk cell_5077 ( .C ( clk ), .D ( signal_10668 ), .Q ( signal_10669 ) ) ;
    buf_clk cell_5085 ( .C ( clk ), .D ( signal_10676 ), .Q ( signal_10677 ) ) ;
    buf_clk cell_5093 ( .C ( clk ), .D ( signal_10684 ), .Q ( signal_10685 ) ) ;
    buf_clk cell_5097 ( .C ( clk ), .D ( signal_9718 ), .Q ( signal_10689 ) ) ;
    buf_clk cell_5101 ( .C ( clk ), .D ( signal_9720 ), .Q ( signal_10693 ) ) ;
    buf_clk cell_5105 ( .C ( clk ), .D ( signal_9722 ), .Q ( signal_10697 ) ) ;
    buf_clk cell_5109 ( .C ( clk ), .D ( signal_2116 ), .Q ( signal_10701 ) ) ;
    buf_clk cell_5113 ( .C ( clk ), .D ( signal_4756 ), .Q ( signal_10705 ) ) ;
    buf_clk cell_5117 ( .C ( clk ), .D ( signal_4757 ), .Q ( signal_10709 ) ) ;
    buf_clk cell_5133 ( .C ( clk ), .D ( signal_2109 ), .Q ( signal_10725 ) ) ;
    buf_clk cell_5137 ( .C ( clk ), .D ( signal_4742 ), .Q ( signal_10729 ) ) ;
    buf_clk cell_5141 ( .C ( clk ), .D ( signal_4743 ), .Q ( signal_10733 ) ) ;
    buf_clk cell_5151 ( .C ( clk ), .D ( signal_10742 ), .Q ( signal_10743 ) ) ;
    buf_clk cell_5161 ( .C ( clk ), .D ( signal_10752 ), .Q ( signal_10753 ) ) ;
    buf_clk cell_5171 ( .C ( clk ), .D ( signal_10762 ), .Q ( signal_10763 ) ) ;
    buf_clk cell_5177 ( .C ( clk ), .D ( signal_10768 ), .Q ( signal_10769 ) ) ;
    buf_clk cell_5183 ( .C ( clk ), .D ( signal_10774 ), .Q ( signal_10775 ) ) ;
    buf_clk cell_5189 ( .C ( clk ), .D ( signal_10780 ), .Q ( signal_10781 ) ) ;
    buf_clk cell_5203 ( .C ( clk ), .D ( signal_10794 ), .Q ( signal_10795 ) ) ;
    buf_clk cell_5211 ( .C ( clk ), .D ( signal_10802 ), .Q ( signal_10803 ) ) ;
    buf_clk cell_5219 ( .C ( clk ), .D ( signal_10810 ), .Q ( signal_10811 ) ) ;
    buf_clk cell_5225 ( .C ( clk ), .D ( signal_10816 ), .Q ( signal_10817 ) ) ;
    buf_clk cell_5231 ( .C ( clk ), .D ( signal_10822 ), .Q ( signal_10823 ) ) ;
    buf_clk cell_5237 ( .C ( clk ), .D ( signal_10828 ), .Q ( signal_10829 ) ) ;
    buf_clk cell_5245 ( .C ( clk ), .D ( signal_10836 ), .Q ( signal_10837 ) ) ;
    buf_clk cell_5253 ( .C ( clk ), .D ( signal_10844 ), .Q ( signal_10845 ) ) ;
    buf_clk cell_5261 ( .C ( clk ), .D ( signal_10852 ), .Q ( signal_10853 ) ) ;
    buf_clk cell_5269 ( .C ( clk ), .D ( signal_10860 ), .Q ( signal_10861 ) ) ;
    buf_clk cell_5277 ( .C ( clk ), .D ( signal_10868 ), .Q ( signal_10869 ) ) ;
    buf_clk cell_5285 ( .C ( clk ), .D ( signal_10876 ), .Q ( signal_10877 ) ) ;
    buf_clk cell_5293 ( .C ( clk ), .D ( signal_10884 ), .Q ( signal_10885 ) ) ;
    buf_clk cell_5301 ( .C ( clk ), .D ( signal_10892 ), .Q ( signal_10893 ) ) ;
    buf_clk cell_5309 ( .C ( clk ), .D ( signal_10900 ), .Q ( signal_10901 ) ) ;
    buf_clk cell_5319 ( .C ( clk ), .D ( signal_10910 ), .Q ( signal_10911 ) ) ;
    buf_clk cell_5329 ( .C ( clk ), .D ( signal_10920 ), .Q ( signal_10921 ) ) ;
    buf_clk cell_5339 ( .C ( clk ), .D ( signal_10930 ), .Q ( signal_10931 ) ) ;
    buf_clk cell_5347 ( .C ( clk ), .D ( signal_10938 ), .Q ( signal_10939 ) ) ;
    buf_clk cell_5355 ( .C ( clk ), .D ( signal_10946 ), .Q ( signal_10947 ) ) ;
    buf_clk cell_5363 ( .C ( clk ), .D ( signal_10954 ), .Q ( signal_10955 ) ) ;
    buf_clk cell_5371 ( .C ( clk ), .D ( signal_10962 ), .Q ( signal_10963 ) ) ;
    buf_clk cell_5379 ( .C ( clk ), .D ( signal_10970 ), .Q ( signal_10971 ) ) ;
    buf_clk cell_5387 ( .C ( clk ), .D ( signal_10978 ), .Q ( signal_10979 ) ) ;
    buf_clk cell_5401 ( .C ( clk ), .D ( signal_10992 ), .Q ( signal_10993 ) ) ;
    buf_clk cell_5409 ( .C ( clk ), .D ( signal_11000 ), .Q ( signal_11001 ) ) ;
    buf_clk cell_5417 ( .C ( clk ), .D ( signal_11008 ), .Q ( signal_11009 ) ) ;
    buf_clk cell_5425 ( .C ( clk ), .D ( signal_11016 ), .Q ( signal_11017 ) ) ;
    buf_clk cell_5433 ( .C ( clk ), .D ( signal_11024 ), .Q ( signal_11025 ) ) ;
    buf_clk cell_5441 ( .C ( clk ), .D ( signal_11032 ), .Q ( signal_11033 ) ) ;
    buf_clk cell_5449 ( .C ( clk ), .D ( signal_11040 ), .Q ( signal_11041 ) ) ;
    buf_clk cell_5457 ( .C ( clk ), .D ( signal_11048 ), .Q ( signal_11049 ) ) ;
    buf_clk cell_5465 ( .C ( clk ), .D ( signal_11056 ), .Q ( signal_11057 ) ) ;
    buf_clk cell_5469 ( .C ( clk ), .D ( signal_1945 ), .Q ( signal_11061 ) ) ;
    buf_clk cell_5475 ( .C ( clk ), .D ( signal_4414 ), .Q ( signal_11067 ) ) ;
    buf_clk cell_5481 ( .C ( clk ), .D ( signal_4415 ), .Q ( signal_11073 ) ) ;
    buf_clk cell_5489 ( .C ( clk ), .D ( signal_11080 ), .Q ( signal_11081 ) ) ;
    buf_clk cell_5497 ( .C ( clk ), .D ( signal_11088 ), .Q ( signal_11089 ) ) ;
    buf_clk cell_5505 ( .C ( clk ), .D ( signal_11096 ), .Q ( signal_11097 ) ) ;
    buf_clk cell_5511 ( .C ( clk ), .D ( signal_2111 ), .Q ( signal_11103 ) ) ;
    buf_clk cell_5517 ( .C ( clk ), .D ( signal_4746 ), .Q ( signal_11109 ) ) ;
    buf_clk cell_5523 ( .C ( clk ), .D ( signal_4747 ), .Q ( signal_11115 ) ) ;
    buf_clk cell_5529 ( .C ( clk ), .D ( signal_1976 ), .Q ( signal_11121 ) ) ;
    buf_clk cell_5535 ( .C ( clk ), .D ( signal_4476 ), .Q ( signal_11127 ) ) ;
    buf_clk cell_5541 ( .C ( clk ), .D ( signal_4477 ), .Q ( signal_11133 ) ) ;
    buf_clk cell_5549 ( .C ( clk ), .D ( signal_11140 ), .Q ( signal_11141 ) ) ;
    buf_clk cell_5557 ( .C ( clk ), .D ( signal_11148 ), .Q ( signal_11149 ) ) ;
    buf_clk cell_5565 ( .C ( clk ), .D ( signal_11156 ), .Q ( signal_11157 ) ) ;
    buf_clk cell_5575 ( .C ( clk ), .D ( signal_11166 ), .Q ( signal_11167 ) ) ;
    buf_clk cell_5585 ( .C ( clk ), .D ( signal_11176 ), .Q ( signal_11177 ) ) ;
    buf_clk cell_5595 ( .C ( clk ), .D ( signal_11186 ), .Q ( signal_11187 ) ) ;
    buf_clk cell_5607 ( .C ( clk ), .D ( signal_2070 ), .Q ( signal_11199 ) ) ;
    buf_clk cell_5613 ( .C ( clk ), .D ( signal_4664 ), .Q ( signal_11205 ) ) ;
    buf_clk cell_5619 ( .C ( clk ), .D ( signal_4665 ), .Q ( signal_11211 ) ) ;
    buf_clk cell_5627 ( .C ( clk ), .D ( signal_11218 ), .Q ( signal_11219 ) ) ;
    buf_clk cell_5635 ( .C ( clk ), .D ( signal_11226 ), .Q ( signal_11227 ) ) ;
    buf_clk cell_5643 ( .C ( clk ), .D ( signal_11234 ), .Q ( signal_11235 ) ) ;
    buf_clk cell_5653 ( .C ( clk ), .D ( signal_11244 ), .Q ( signal_11245 ) ) ;
    buf_clk cell_5663 ( .C ( clk ), .D ( signal_11254 ), .Q ( signal_11255 ) ) ;
    buf_clk cell_5673 ( .C ( clk ), .D ( signal_11264 ), .Q ( signal_11265 ) ) ;
    buf_clk cell_5681 ( .C ( clk ), .D ( signal_11272 ), .Q ( signal_11273 ) ) ;
    buf_clk cell_5689 ( .C ( clk ), .D ( signal_11280 ), .Q ( signal_11281 ) ) ;
    buf_clk cell_5697 ( .C ( clk ), .D ( signal_11288 ), .Q ( signal_11289 ) ) ;
    buf_clk cell_5703 ( .C ( clk ), .D ( signal_1890 ), .Q ( signal_11295 ) ) ;
    buf_clk cell_5709 ( .C ( clk ), .D ( signal_4304 ), .Q ( signal_11301 ) ) ;
    buf_clk cell_5715 ( .C ( clk ), .D ( signal_4305 ), .Q ( signal_11307 ) ) ;
    buf_clk cell_5721 ( .C ( clk ), .D ( signal_2002 ), .Q ( signal_11313 ) ) ;
    buf_clk cell_5727 ( .C ( clk ), .D ( signal_4528 ), .Q ( signal_11319 ) ) ;
    buf_clk cell_5733 ( .C ( clk ), .D ( signal_4529 ), .Q ( signal_11325 ) ) ;
    buf_clk cell_5769 ( .C ( clk ), .D ( signal_2106 ), .Q ( signal_11361 ) ) ;
    buf_clk cell_5775 ( .C ( clk ), .D ( signal_4736 ), .Q ( signal_11367 ) ) ;
    buf_clk cell_5781 ( .C ( clk ), .D ( signal_4737 ), .Q ( signal_11373 ) ) ;
    buf_clk cell_5793 ( .C ( clk ), .D ( signal_2068 ), .Q ( signal_11385 ) ) ;
    buf_clk cell_5799 ( .C ( clk ), .D ( signal_4660 ), .Q ( signal_11391 ) ) ;
    buf_clk cell_5805 ( .C ( clk ), .D ( signal_4661 ), .Q ( signal_11397 ) ) ;
    buf_clk cell_5823 ( .C ( clk ), .D ( signal_2073 ), .Q ( signal_11415 ) ) ;
    buf_clk cell_5829 ( .C ( clk ), .D ( signal_4670 ), .Q ( signal_11421 ) ) ;
    buf_clk cell_5835 ( .C ( clk ), .D ( signal_4671 ), .Q ( signal_11427 ) ) ;
    buf_clk cell_5877 ( .C ( clk ), .D ( signal_2110 ), .Q ( signal_11469 ) ) ;
    buf_clk cell_5885 ( .C ( clk ), .D ( signal_4744 ), .Q ( signal_11477 ) ) ;
    buf_clk cell_5893 ( .C ( clk ), .D ( signal_4745 ), .Q ( signal_11485 ) ) ;
    buf_clk cell_5921 ( .C ( clk ), .D ( signal_11512 ), .Q ( signal_11513 ) ) ;
    buf_clk cell_5931 ( .C ( clk ), .D ( signal_11522 ), .Q ( signal_11523 ) ) ;
    buf_clk cell_5941 ( .C ( clk ), .D ( signal_11532 ), .Q ( signal_11533 ) ) ;
    buf_clk cell_5979 ( .C ( clk ), .D ( signal_9792 ), .Q ( signal_11571 ) ) ;
    buf_clk cell_5987 ( .C ( clk ), .D ( signal_9796 ), .Q ( signal_11579 ) ) ;
    buf_clk cell_5995 ( .C ( clk ), .D ( signal_9800 ), .Q ( signal_11587 ) ) ;
    buf_clk cell_6021 ( .C ( clk ), .D ( signal_1986 ), .Q ( signal_11613 ) ) ;
    buf_clk cell_6029 ( .C ( clk ), .D ( signal_4496 ), .Q ( signal_11621 ) ) ;
    buf_clk cell_6037 ( .C ( clk ), .D ( signal_4497 ), .Q ( signal_11629 ) ) ;
    buf_clk cell_6063 ( .C ( clk ), .D ( signal_2082 ), .Q ( signal_11655 ) ) ;
    buf_clk cell_6071 ( .C ( clk ), .D ( signal_4688 ), .Q ( signal_11663 ) ) ;
    buf_clk cell_6079 ( .C ( clk ), .D ( signal_4689 ), .Q ( signal_11671 ) ) ;
    buf_clk cell_6185 ( .C ( clk ), .D ( signal_11776 ), .Q ( signal_11777 ) ) ;
    buf_clk cell_6197 ( .C ( clk ), .D ( signal_11788 ), .Q ( signal_11789 ) ) ;
    buf_clk cell_6209 ( .C ( clk ), .D ( signal_11800 ), .Q ( signal_11801 ) ) ;
    buf_clk cell_6259 ( .C ( clk ), .D ( signal_11850 ), .Q ( signal_11851 ) ) ;
    buf_clk cell_6273 ( .C ( clk ), .D ( signal_11864 ), .Q ( signal_11865 ) ) ;
    buf_clk cell_6287 ( .C ( clk ), .D ( signal_11878 ), .Q ( signal_11879 ) ) ;
    buf_clk cell_6325 ( .C ( clk ), .D ( signal_11916 ), .Q ( signal_11917 ) ) ;
    buf_clk cell_6339 ( .C ( clk ), .D ( signal_11930 ), .Q ( signal_11931 ) ) ;
    buf_clk cell_6353 ( .C ( clk ), .D ( signal_11944 ), .Q ( signal_11945 ) ) ;
    buf_clk cell_6445 ( .C ( clk ), .D ( signal_12036 ), .Q ( signal_12037 ) ) ;
    buf_clk cell_6461 ( .C ( clk ), .D ( signal_12052 ), .Q ( signal_12053 ) ) ;
    buf_clk cell_6477 ( .C ( clk ), .D ( signal_12068 ), .Q ( signal_12069 ) ) ;
    buf_clk cell_6505 ( .C ( clk ), .D ( signal_12096 ), .Q ( signal_12097 ) ) ;
    buf_clk cell_6521 ( .C ( clk ), .D ( signal_12112 ), .Q ( signal_12113 ) ) ;
    buf_clk cell_6537 ( .C ( clk ), .D ( signal_12128 ), .Q ( signal_12129 ) ) ;
    buf_clk cell_6689 ( .C ( clk ), .D ( signal_12280 ), .Q ( signal_12281 ) ) ;
    buf_clk cell_6705 ( .C ( clk ), .D ( signal_12296 ), .Q ( signal_12297 ) ) ;
    buf_clk cell_6721 ( .C ( clk ), .D ( signal_12312 ), .Q ( signal_12313 ) ) ;
    buf_clk cell_6739 ( .C ( clk ), .D ( signal_12330 ), .Q ( signal_12331 ) ) ;
    buf_clk cell_6757 ( .C ( clk ), .D ( signal_12348 ), .Q ( signal_12349 ) ) ;
    buf_clk cell_6775 ( .C ( clk ), .D ( signal_12366 ), .Q ( signal_12367 ) ) ;
    buf_clk cell_6889 ( .C ( clk ), .D ( signal_12480 ), .Q ( signal_12481 ) ) ;
    buf_clk cell_6909 ( .C ( clk ), .D ( signal_12500 ), .Q ( signal_12501 ) ) ;
    buf_clk cell_6929 ( .C ( clk ), .D ( signal_12520 ), .Q ( signal_12521 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2027 ( .a ({signal_9488, signal_9486, signal_9484}), .b ({signal_4377, signal_4376, signal_1926}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995]}), .c ({signal_4609, signal_4608, signal_2042}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2032 ( .a ({signal_9506, signal_9500, signal_9494}), .b ({signal_4299, signal_4298, signal_1887}), .clk ( clk ), .r ({Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({signal_4619, signal_4618, signal_2047}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2037 ( .a ({signal_9524, signal_9518, signal_9512}), .b ({signal_4405, signal_4404, signal_1940}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001]}), .c ({signal_4629, signal_4628, signal_2052}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2038 ( .a ({signal_9542, signal_9536, signal_9530}), .b ({signal_4411, signal_4410, signal_1943}), .clk ( clk ), .r ({Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({signal_4631, signal_4630, signal_2053}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2039 ( .a ({signal_9554, signal_9550, signal_9546}), .b ({signal_4417, signal_4416, signal_1946}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007]}), .c ({signal_4633, signal_4632, signal_2054}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2040 ( .a ({signal_9572, signal_9566, signal_9560}), .b ({signal_4421, signal_4420, signal_1948}), .clk ( clk ), .r ({Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_4635, signal_4634, signal_2055}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2041 ( .a ({signal_9584, signal_9580, signal_9576}), .b ({signal_4425, signal_4424, signal_1950}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013]}), .c ({signal_4637, signal_4636, signal_2056}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2042 ( .a ({signal_9596, signal_9592, signal_9588}), .b ({signal_4433, signal_4432, signal_1954}), .clk ( clk ), .r ({Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({signal_4639, signal_4638, signal_2057}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2043 ( .a ({signal_9608, signal_9604, signal_9600}), .b ({signal_4435, signal_4434, signal_1955}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019]}), .c ({signal_4641, signal_4640, signal_2058}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2044 ( .a ({signal_9620, signal_9616, signal_9612}), .b ({signal_4437, signal_4436, signal_1956}), .clk ( clk ), .r ({Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({signal_4643, signal_4642, signal_2059}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2045 ( .a ({signal_9632, signal_9628, signal_9624}), .b ({signal_4447, signal_4446, signal_1961}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025]}), .c ({signal_4645, signal_4644, signal_2060}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2064 ( .a ({signal_4609, signal_4608, signal_2042}), .b ({signal_4683, signal_4682, signal_2079}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2068 ( .a ({signal_4619, signal_4618, signal_2047}), .b ({signal_4691, signal_4690, signal_2083}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2072 ( .a ({signal_4629, signal_4628, signal_2052}), .b ({signal_4699, signal_4698, signal_2087}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2073 ( .a ({signal_4641, signal_4640, signal_2058}), .b ({signal_4701, signal_4700, signal_2088}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2084 ( .a ({signal_9650, signal_9644, signal_9638}), .b ({signal_4493, signal_4492, signal_1984}), .clk ( clk ), .r ({Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({signal_4723, signal_4722, signal_2099}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2090 ( .a ({signal_9662, signal_9658, signal_9654}), .b ({signal_4511, signal_4510, signal_1993}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031]}), .c ({signal_4735, signal_4734, signal_2105}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2098 ( .a ({signal_4391, signal_4390, signal_1933}), .b ({signal_9668, signal_9666, signal_9664}), .clk ( clk ), .r ({Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({signal_4751, signal_4750, signal_2113}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2100 ( .a ({signal_9674, signal_9672, signal_9670}), .b ({signal_4527, signal_4526, signal_2001}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037]}), .c ({signal_4755, signal_4754, signal_2115}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2102 ( .a ({signal_9680, signal_9678, signal_9676}), .b ({signal_4533, signal_4532, signal_2004}), .clk ( clk ), .r ({Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_4759, signal_4758, signal_2117}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2103 ( .a ({signal_9686, signal_9684, signal_9682}), .b ({signal_4407, signal_4406, signal_1941}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043]}), .c ({signal_4761, signal_4760, signal_2118}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2105 ( .a ({signal_9692, signal_9690, signal_9688}), .b ({signal_4407, signal_4406, signal_1941}), .clk ( clk ), .r ({Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({signal_4765, signal_4764, signal_2120}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2106 ( .a ({signal_9704, signal_9700, signal_9696}), .b ({signal_4605, signal_4604, signal_2040}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049]}), .c ({signal_4767, signal_4766, signal_2121}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2107 ( .a ({signal_9710, signal_9708, signal_9706}), .b ({signal_4413, signal_4412, signal_1944}), .clk ( clk ), .r ({Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({signal_4769, signal_4768, signal_2122}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2108 ( .a ({signal_9716, signal_9714, signal_9712}), .b ({signal_4615, signal_4614, signal_2045}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055]}), .c ({signal_4771, signal_4770, signal_2123}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2109 ( .a ({signal_9722, signal_9720, signal_9718}), .b ({signal_4539, signal_4538, signal_2007}), .clk ( clk ), .r ({Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({signal_4773, signal_4772, signal_2124}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2111 ( .a ({signal_9740, signal_9734, signal_9728}), .b ({signal_4541, signal_4540, signal_2008}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061]}), .c ({signal_4777, signal_4776, signal_2126}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2112 ( .a ({signal_9746, signal_9744, signal_9742}), .b ({signal_4429, signal_4428, signal_1952}), .clk ( clk ), .r ({Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({signal_4779, signal_4778, signal_2127}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2113 ( .a ({signal_9758, signal_9754, signal_9750}), .b ({signal_4623, signal_4622, signal_2049}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067]}), .c ({signal_4781, signal_4780, signal_2128}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2114 ( .a ({signal_9764, signal_9762, signal_9760}), .b ({signal_4543, signal_4542, signal_2009}), .clk ( clk ), .r ({Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_4783, signal_4782, signal_2129}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2115 ( .a ({signal_9650, signal_9644, signal_9638}), .b ({signal_4545, signal_4544, signal_2010}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073]}), .c ({signal_4785, signal_4784, signal_2130}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2117 ( .a ({signal_9770, signal_9768, signal_9766}), .b ({signal_4549, signal_4548, signal_2012}), .clk ( clk ), .r ({Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({signal_4789, signal_4788, signal_2132}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2120 ( .a ({signal_9662, signal_9658, signal_9654}), .b ({signal_4551, signal_4550, signal_2013}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079]}), .c ({signal_4795, signal_4794, signal_2135}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2129 ( .a ({signal_4723, signal_4722, signal_2099}), .b ({signal_4813, signal_4812, signal_2144}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2131 ( .a ({signal_4735, signal_4734, signal_2105}), .b ({signal_4817, signal_4816, signal_2146}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2132 ( .a ({signal_4755, signal_4754, signal_2115}), .b ({signal_4819, signal_4818, signal_2147}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2134 ( .a ({signal_4773, signal_4772, signal_2124}), .b ({signal_4823, signal_4822, signal_2149}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2136 ( .a ({signal_4777, signal_4776, signal_2126}), .b ({signal_4827, signal_4826, signal_2151}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2137 ( .a ({signal_4783, signal_4782, signal_2129}), .b ({signal_4829, signal_4828, signal_2152}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2138 ( .a ({signal_4785, signal_4784, signal_2130}), .b ({signal_4831, signal_4830, signal_2153}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2139 ( .a ({signal_4789, signal_4788, signal_2132}), .b ({signal_4833, signal_4832, signal_2154}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2141 ( .a ({signal_4795, signal_4794, signal_2135}), .b ({signal_4837, signal_4836, signal_2156}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2142 ( .a ({signal_9788, signal_9782, signal_9776}), .b ({signal_4647, signal_4646, signal_2061}), .clk ( clk ), .r ({Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({signal_4839, signal_4838, signal_2157}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2143 ( .a ({signal_9800, signal_9796, signal_9792}), .b ({signal_4649, signal_4648, signal_2062}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085]}), .c ({signal_4841, signal_4840, signal_2158}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2145 ( .a ({signal_9806, signal_9804, signal_9802}), .b ({signal_4705, signal_4704, signal_2090}), .clk ( clk ), .r ({Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({signal_4845, signal_4844, signal_2160}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2146 ( .a ({signal_4655, signal_4654, signal_2065}), .b ({signal_9812, signal_9810, signal_9808}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091]}), .c ({signal_4847, signal_4846, signal_2161}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2147 ( .a ({signal_9824, signal_9820, signal_9816}), .b ({signal_4657, signal_4656, signal_2066}), .clk ( clk ), .r ({Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({signal_4849, signal_4848, signal_2162}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2149 ( .a ({signal_9836, signal_9832, signal_9828}), .b ({signal_4711, signal_4710, signal_2093}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097]}), .c ({signal_4853, signal_4852, signal_2164}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2150 ( .a ({signal_9848, signal_9844, signal_9840}), .b ({signal_4713, signal_4712, signal_2094}), .clk ( clk ), .r ({Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_4855, signal_4854, signal_2165}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2151 ( .a ({signal_9854, signal_9852, signal_9850}), .b ({signal_4669, signal_4668, signal_2072}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103]}), .c ({signal_4857, signal_4856, signal_2166}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2152 ( .a ({signal_9872, signal_9866, signal_9860}), .b ({signal_4715, signal_4714, signal_2095}), .clk ( clk ), .r ({Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({signal_4859, signal_4858, signal_2167}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2153 ( .a ({signal_9884, signal_9880, signal_9876}), .b ({signal_4721, signal_4720, signal_2098}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109]}), .c ({signal_4861, signal_4860, signal_2168}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2154 ( .a ({signal_9902, signal_9896, signal_9890}), .b ({signal_4675, signal_4674, signal_2075}), .clk ( clk ), .r ({Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({signal_4863, signal_4862, signal_2169}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2155 ( .a ({signal_4653, signal_4652, signal_2064}), .b ({signal_4677, signal_4676, signal_2076}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115]}), .c ({signal_4865, signal_4864, signal_2170}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2156 ( .a ({signal_9914, signal_9910, signal_9906}), .b ({signal_4679, signal_4678, signal_2077}), .clk ( clk ), .r ({Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({signal_4867, signal_4866, signal_2171}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2157 ( .a ({signal_9506, signal_9500, signal_9494}), .b ({signal_4681, signal_4680, signal_2078}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121]}), .c ({signal_4869, signal_4868, signal_2172}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2158 ( .a ({signal_9926, signal_9922, signal_9918}), .b ({signal_4725, signal_4724, signal_2100}), .clk ( clk ), .r ({Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({signal_4871, signal_4870, signal_2173}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2159 ( .a ({signal_9938, signal_9934, signal_9930}), .b ({signal_4729, signal_4728, signal_2102}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127]}), .c ({signal_4873, signal_4872, signal_2174}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2160 ( .a ({signal_9944, signal_9942, signal_9940}), .b ({signal_4731, signal_4730, signal_2103}), .clk ( clk ), .r ({Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_4875, signal_4874, signal_2175}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2161 ( .a ({signal_9956, signal_9952, signal_9948}), .b ({signal_4733, signal_4732, signal_2104}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133]}), .c ({signal_4877, signal_4876, signal_2176}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2163 ( .a ({signal_9968, signal_9964, signal_9960}), .b ({signal_4685, signal_4684, signal_2080}), .clk ( clk ), .r ({Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({signal_4881, signal_4880, signal_2178}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2164 ( .a ({signal_9986, signal_9980, signal_9974}), .b ({signal_4739, signal_4738, signal_2107}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139]}), .c ({signal_4883, signal_4882, signal_2179}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2165 ( .a ({signal_4741, signal_4740, signal_2108}), .b ({signal_4431, signal_4430, signal_1953}), .clk ( clk ), .r ({Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({signal_4885, signal_4884, signal_2180}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2166 ( .a ({signal_9506, signal_9500, signal_9494}), .b ({signal_4693, signal_4692, signal_2084}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145]}), .c ({signal_4887, signal_4886, signal_2181}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2167 ( .a ({signal_4695, signal_4694, signal_2085}), .b ({signal_9992, signal_9990, signal_9988}), .clk ( clk ), .r ({Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({signal_4889, signal_4888, signal_2182}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2168 ( .a ({signal_9998, signal_9996, signal_9994}), .b ({signal_4749, signal_4748, signal_2112}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151]}), .c ({signal_4891, signal_4890, signal_2183}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2169 ( .a ({signal_10010, signal_10006, signal_10002}), .b ({signal_4697, signal_4696, signal_2086}), .clk ( clk ), .r ({Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({signal_4893, signal_4892, signal_2184}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2171 ( .a ({signal_10028, signal_10022, signal_10016}), .b ({signal_4753, signal_4752, signal_2114}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157]}), .c ({signal_4897, signal_4896, signal_2186}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2184 ( .a ({signal_4841, signal_4840, signal_2158}), .b ({signal_4923, signal_4922, signal_2199}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2187 ( .a ({signal_4857, signal_4856, signal_2166}), .b ({signal_4929, signal_4928, signal_2202}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2188 ( .a ({signal_4869, signal_4868, signal_2172}), .b ({signal_4931, signal_4930, signal_2203}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2189 ( .a ({signal_4873, signal_4872, signal_2174}), .b ({signal_4933, signal_4932, signal_2204}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2191 ( .a ({signal_4883, signal_4882, signal_2179}), .b ({signal_4937, signal_4936, signal_2206}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2192 ( .a ({signal_4885, signal_4884, signal_2180}), .b ({signal_4939, signal_4938, signal_2207}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2193 ( .a ({signal_4887, signal_4886, signal_2181}), .b ({signal_4941, signal_4940, signal_2208}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2194 ( .a ({signal_4897, signal_4896, signal_2186}), .b ({signal_4943, signal_4942, signal_2209}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2201 ( .a ({signal_10046, signal_10040, signal_10034}), .b ({signal_4803, signal_4802, signal_2139}), .clk ( clk ), .r ({Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_4957, signal_4956, signal_2216}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2202 ( .a ({signal_10064, signal_10058, signal_10052}), .b ({signal_4805, signal_4804, signal_2140}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163]}), .c ({signal_4959, signal_4958, signal_2217}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2203 ( .a ({signal_10076, signal_10072, signal_10068}), .b ({signal_4807, signal_4806, signal_2141}), .clk ( clk ), .r ({Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({signal_4961, signal_4960, signal_2218}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2204 ( .a ({signal_9506, signal_9500, signal_9494}), .b ({signal_4809, signal_4808, signal_2142}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169]}), .c ({signal_4963, signal_4962, signal_2219}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2205 ( .a ({signal_10082, signal_10080, signal_10078}), .b ({signal_4811, signal_4810, signal_2143}), .clk ( clk ), .r ({Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({signal_4965, signal_4964, signal_2220}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2206 ( .a ({signal_9764, signal_9762, signal_9760}), .b ({signal_4815, signal_4814, signal_2145}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175]}), .c ({signal_4967, signal_4966, signal_2221}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2213 ( .a ({signal_10088, signal_10086, signal_10084}), .b ({signal_4821, signal_4820, signal_2148}), .clk ( clk ), .r ({Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({signal_4981, signal_4980, signal_2228}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2221 ( .a ({signal_10064, signal_10058, signal_10052}), .b ({signal_4825, signal_4824, signal_2150}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181]}), .c ({signal_4997, signal_4996, signal_2236}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2233 ( .a ({signal_4957, signal_4956, signal_2216}), .b ({signal_5021, signal_5020, signal_2248}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2234 ( .a ({signal_4959, signal_4958, signal_2217}), .b ({signal_5023, signal_5022, signal_2249}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2235 ( .a ({signal_4961, signal_4960, signal_2218}), .b ({signal_5025, signal_5024, signal_2250}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2236 ( .a ({signal_4963, signal_4962, signal_2219}), .b ({signal_5027, signal_5026, signal_2251}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2237 ( .a ({signal_4965, signal_4964, signal_2220}), .b ({signal_5029, signal_5028, signal_2252}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2238 ( .a ({signal_4967, signal_4966, signal_2221}), .b ({signal_5031, signal_5030, signal_2253}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2240 ( .a ({signal_4981, signal_4980, signal_2228}), .b ({signal_5035, signal_5034, signal_2255}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2242 ( .a ({signal_4997, signal_4996, signal_2236}), .b ({signal_5039, signal_5038, signal_2257}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2248 ( .a ({signal_4673, signal_4672, signal_2074}), .b ({signal_4925, signal_4924, signal_2200}), .clk ( clk ), .r ({Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({signal_5051, signal_5050, signal_2263}) ) ;
    buf_clk cell_4504 ( .C ( clk ), .D ( signal_10095 ), .Q ( signal_10096 ) ) ;
    buf_clk cell_4512 ( .C ( clk ), .D ( signal_10103 ), .Q ( signal_10104 ) ) ;
    buf_clk cell_4520 ( .C ( clk ), .D ( signal_10111 ), .Q ( signal_10112 ) ) ;
    buf_clk cell_4524 ( .C ( clk ), .D ( signal_10115 ), .Q ( signal_10116 ) ) ;
    buf_clk cell_4528 ( .C ( clk ), .D ( signal_10119 ), .Q ( signal_10120 ) ) ;
    buf_clk cell_4532 ( .C ( clk ), .D ( signal_10123 ), .Q ( signal_10124 ) ) ;
    buf_clk cell_4538 ( .C ( clk ), .D ( signal_10129 ), .Q ( signal_10130 ) ) ;
    buf_clk cell_4544 ( .C ( clk ), .D ( signal_10135 ), .Q ( signal_10136 ) ) ;
    buf_clk cell_4550 ( .C ( clk ), .D ( signal_10141 ), .Q ( signal_10142 ) ) ;
    buf_clk cell_4556 ( .C ( clk ), .D ( signal_10147 ), .Q ( signal_10148 ) ) ;
    buf_clk cell_4562 ( .C ( clk ), .D ( signal_10153 ), .Q ( signal_10154 ) ) ;
    buf_clk cell_4568 ( .C ( clk ), .D ( signal_10159 ), .Q ( signal_10160 ) ) ;
    buf_clk cell_4572 ( .C ( clk ), .D ( signal_10163 ), .Q ( signal_10164 ) ) ;
    buf_clk cell_4576 ( .C ( clk ), .D ( signal_10167 ), .Q ( signal_10168 ) ) ;
    buf_clk cell_4580 ( .C ( clk ), .D ( signal_10171 ), .Q ( signal_10172 ) ) ;
    buf_clk cell_4586 ( .C ( clk ), .D ( signal_10177 ), .Q ( signal_10178 ) ) ;
    buf_clk cell_4592 ( .C ( clk ), .D ( signal_10183 ), .Q ( signal_10184 ) ) ;
    buf_clk cell_4598 ( .C ( clk ), .D ( signal_10189 ), .Q ( signal_10190 ) ) ;
    buf_clk cell_4602 ( .C ( clk ), .D ( signal_10193 ), .Q ( signal_10194 ) ) ;
    buf_clk cell_4606 ( .C ( clk ), .D ( signal_10197 ), .Q ( signal_10198 ) ) ;
    buf_clk cell_4610 ( .C ( clk ), .D ( signal_10201 ), .Q ( signal_10202 ) ) ;
    buf_clk cell_4614 ( .C ( clk ), .D ( signal_10205 ), .Q ( signal_10206 ) ) ;
    buf_clk cell_4618 ( .C ( clk ), .D ( signal_10209 ), .Q ( signal_10210 ) ) ;
    buf_clk cell_4622 ( .C ( clk ), .D ( signal_10213 ), .Q ( signal_10214 ) ) ;
    buf_clk cell_4624 ( .C ( clk ), .D ( signal_10215 ), .Q ( signal_10216 ) ) ;
    buf_clk cell_4626 ( .C ( clk ), .D ( signal_10217 ), .Q ( signal_10218 ) ) ;
    buf_clk cell_4628 ( .C ( clk ), .D ( signal_10219 ), .Q ( signal_10220 ) ) ;
    buf_clk cell_4630 ( .C ( clk ), .D ( signal_10221 ), .Q ( signal_10222 ) ) ;
    buf_clk cell_4632 ( .C ( clk ), .D ( signal_10223 ), .Q ( signal_10224 ) ) ;
    buf_clk cell_4634 ( .C ( clk ), .D ( signal_10225 ), .Q ( signal_10226 ) ) ;
    buf_clk cell_4640 ( .C ( clk ), .D ( signal_10231 ), .Q ( signal_10232 ) ) ;
    buf_clk cell_4646 ( .C ( clk ), .D ( signal_10237 ), .Q ( signal_10238 ) ) ;
    buf_clk cell_4652 ( .C ( clk ), .D ( signal_10243 ), .Q ( signal_10244 ) ) ;
    buf_clk cell_4658 ( .C ( clk ), .D ( signal_10249 ), .Q ( signal_10250 ) ) ;
    buf_clk cell_4664 ( .C ( clk ), .D ( signal_10255 ), .Q ( signal_10256 ) ) ;
    buf_clk cell_4670 ( .C ( clk ), .D ( signal_10261 ), .Q ( signal_10262 ) ) ;
    buf_clk cell_4676 ( .C ( clk ), .D ( signal_10267 ), .Q ( signal_10268 ) ) ;
    buf_clk cell_4682 ( .C ( clk ), .D ( signal_10273 ), .Q ( signal_10274 ) ) ;
    buf_clk cell_4688 ( .C ( clk ), .D ( signal_10279 ), .Q ( signal_10280 ) ) ;
    buf_clk cell_4690 ( .C ( clk ), .D ( signal_10281 ), .Q ( signal_10282 ) ) ;
    buf_clk cell_4692 ( .C ( clk ), .D ( signal_10283 ), .Q ( signal_10284 ) ) ;
    buf_clk cell_4694 ( .C ( clk ), .D ( signal_10285 ), .Q ( signal_10286 ) ) ;
    buf_clk cell_4698 ( .C ( clk ), .D ( signal_10289 ), .Q ( signal_10290 ) ) ;
    buf_clk cell_4702 ( .C ( clk ), .D ( signal_10293 ), .Q ( signal_10294 ) ) ;
    buf_clk cell_4706 ( .C ( clk ), .D ( signal_10297 ), .Q ( signal_10298 ) ) ;
    buf_clk cell_4712 ( .C ( clk ), .D ( signal_10303 ), .Q ( signal_10304 ) ) ;
    buf_clk cell_4718 ( .C ( clk ), .D ( signal_10309 ), .Q ( signal_10310 ) ) ;
    buf_clk cell_4724 ( .C ( clk ), .D ( signal_10315 ), .Q ( signal_10316 ) ) ;
    buf_clk cell_4726 ( .C ( clk ), .D ( signal_10317 ), .Q ( signal_10318 ) ) ;
    buf_clk cell_4728 ( .C ( clk ), .D ( signal_10319 ), .Q ( signal_10320 ) ) ;
    buf_clk cell_4730 ( .C ( clk ), .D ( signal_10321 ), .Q ( signal_10322 ) ) ;
    buf_clk cell_4736 ( .C ( clk ), .D ( signal_10327 ), .Q ( signal_10328 ) ) ;
    buf_clk cell_4742 ( .C ( clk ), .D ( signal_10333 ), .Q ( signal_10334 ) ) ;
    buf_clk cell_4748 ( .C ( clk ), .D ( signal_10339 ), .Q ( signal_10340 ) ) ;
    buf_clk cell_4750 ( .C ( clk ), .D ( signal_10341 ), .Q ( signal_10342 ) ) ;
    buf_clk cell_4752 ( .C ( clk ), .D ( signal_10343 ), .Q ( signal_10344 ) ) ;
    buf_clk cell_4754 ( .C ( clk ), .D ( signal_10345 ), .Q ( signal_10346 ) ) ;
    buf_clk cell_4762 ( .C ( clk ), .D ( signal_10353 ), .Q ( signal_10354 ) ) ;
    buf_clk cell_4770 ( .C ( clk ), .D ( signal_10361 ), .Q ( signal_10362 ) ) ;
    buf_clk cell_4778 ( .C ( clk ), .D ( signal_10369 ), .Q ( signal_10370 ) ) ;
    buf_clk cell_4782 ( .C ( clk ), .D ( signal_10373 ), .Q ( signal_10374 ) ) ;
    buf_clk cell_4786 ( .C ( clk ), .D ( signal_10377 ), .Q ( signal_10378 ) ) ;
    buf_clk cell_4790 ( .C ( clk ), .D ( signal_10381 ), .Q ( signal_10382 ) ) ;
    buf_clk cell_4794 ( .C ( clk ), .D ( signal_10385 ), .Q ( signal_10386 ) ) ;
    buf_clk cell_4798 ( .C ( clk ), .D ( signal_10389 ), .Q ( signal_10390 ) ) ;
    buf_clk cell_4802 ( .C ( clk ), .D ( signal_10393 ), .Q ( signal_10394 ) ) ;
    buf_clk cell_4808 ( .C ( clk ), .D ( signal_10399 ), .Q ( signal_10400 ) ) ;
    buf_clk cell_4814 ( .C ( clk ), .D ( signal_10405 ), .Q ( signal_10406 ) ) ;
    buf_clk cell_4820 ( .C ( clk ), .D ( signal_10411 ), .Q ( signal_10412 ) ) ;
    buf_clk cell_4826 ( .C ( clk ), .D ( signal_10417 ), .Q ( signal_10418 ) ) ;
    buf_clk cell_4832 ( .C ( clk ), .D ( signal_10423 ), .Q ( signal_10424 ) ) ;
    buf_clk cell_4838 ( .C ( clk ), .D ( signal_10429 ), .Q ( signal_10430 ) ) ;
    buf_clk cell_4842 ( .C ( clk ), .D ( signal_10433 ), .Q ( signal_10434 ) ) ;
    buf_clk cell_4846 ( .C ( clk ), .D ( signal_10437 ), .Q ( signal_10438 ) ) ;
    buf_clk cell_4850 ( .C ( clk ), .D ( signal_10441 ), .Q ( signal_10442 ) ) ;
    buf_clk cell_4858 ( .C ( clk ), .D ( signal_10449 ), .Q ( signal_10450 ) ) ;
    buf_clk cell_4866 ( .C ( clk ), .D ( signal_10457 ), .Q ( signal_10458 ) ) ;
    buf_clk cell_4874 ( .C ( clk ), .D ( signal_10465 ), .Q ( signal_10466 ) ) ;
    buf_clk cell_4880 ( .C ( clk ), .D ( signal_10471 ), .Q ( signal_10472 ) ) ;
    buf_clk cell_4886 ( .C ( clk ), .D ( signal_10477 ), .Q ( signal_10478 ) ) ;
    buf_clk cell_4892 ( .C ( clk ), .D ( signal_10483 ), .Q ( signal_10484 ) ) ;
    buf_clk cell_4898 ( .C ( clk ), .D ( signal_10489 ), .Q ( signal_10490 ) ) ;
    buf_clk cell_4904 ( .C ( clk ), .D ( signal_10495 ), .Q ( signal_10496 ) ) ;
    buf_clk cell_4910 ( .C ( clk ), .D ( signal_10501 ), .Q ( signal_10502 ) ) ;
    buf_clk cell_4912 ( .C ( clk ), .D ( signal_10503 ), .Q ( signal_10504 ) ) ;
    buf_clk cell_4914 ( .C ( clk ), .D ( signal_10505 ), .Q ( signal_10506 ) ) ;
    buf_clk cell_4916 ( .C ( clk ), .D ( signal_10507 ), .Q ( signal_10508 ) ) ;
    buf_clk cell_4918 ( .C ( clk ), .D ( signal_10509 ), .Q ( signal_10510 ) ) ;
    buf_clk cell_4920 ( .C ( clk ), .D ( signal_10511 ), .Q ( signal_10512 ) ) ;
    buf_clk cell_4922 ( .C ( clk ), .D ( signal_10513 ), .Q ( signal_10514 ) ) ;
    buf_clk cell_4928 ( .C ( clk ), .D ( signal_10519 ), .Q ( signal_10520 ) ) ;
    buf_clk cell_4934 ( .C ( clk ), .D ( signal_10525 ), .Q ( signal_10526 ) ) ;
    buf_clk cell_4940 ( .C ( clk ), .D ( signal_10531 ), .Q ( signal_10532 ) ) ;
    buf_clk cell_4942 ( .C ( clk ), .D ( signal_10533 ), .Q ( signal_10534 ) ) ;
    buf_clk cell_4944 ( .C ( clk ), .D ( signal_10535 ), .Q ( signal_10536 ) ) ;
    buf_clk cell_4946 ( .C ( clk ), .D ( signal_10537 ), .Q ( signal_10538 ) ) ;
    buf_clk cell_4948 ( .C ( clk ), .D ( signal_10539 ), .Q ( signal_10540 ) ) ;
    buf_clk cell_4950 ( .C ( clk ), .D ( signal_10541 ), .Q ( signal_10542 ) ) ;
    buf_clk cell_4952 ( .C ( clk ), .D ( signal_10543 ), .Q ( signal_10544 ) ) ;
    buf_clk cell_4958 ( .C ( clk ), .D ( signal_10549 ), .Q ( signal_10550 ) ) ;
    buf_clk cell_4964 ( .C ( clk ), .D ( signal_10555 ), .Q ( signal_10556 ) ) ;
    buf_clk cell_4970 ( .C ( clk ), .D ( signal_10561 ), .Q ( signal_10562 ) ) ;
    buf_clk cell_4976 ( .C ( clk ), .D ( signal_10567 ), .Q ( signal_10568 ) ) ;
    buf_clk cell_4982 ( .C ( clk ), .D ( signal_10573 ), .Q ( signal_10574 ) ) ;
    buf_clk cell_4988 ( .C ( clk ), .D ( signal_10579 ), .Q ( signal_10580 ) ) ;
    buf_clk cell_4992 ( .C ( clk ), .D ( signal_10583 ), .Q ( signal_10584 ) ) ;
    buf_clk cell_4996 ( .C ( clk ), .D ( signal_10587 ), .Q ( signal_10588 ) ) ;
    buf_clk cell_5000 ( .C ( clk ), .D ( signal_10591 ), .Q ( signal_10592 ) ) ;
    buf_clk cell_5008 ( .C ( clk ), .D ( signal_10599 ), .Q ( signal_10600 ) ) ;
    buf_clk cell_5018 ( .C ( clk ), .D ( signal_10609 ), .Q ( signal_10610 ) ) ;
    buf_clk cell_5028 ( .C ( clk ), .D ( signal_10619 ), .Q ( signal_10620 ) ) ;
    buf_clk cell_5034 ( .C ( clk ), .D ( signal_10625 ), .Q ( signal_10626 ) ) ;
    buf_clk cell_5040 ( .C ( clk ), .D ( signal_10631 ), .Q ( signal_10632 ) ) ;
    buf_clk cell_5046 ( .C ( clk ), .D ( signal_10637 ), .Q ( signal_10638 ) ) ;
    buf_clk cell_5054 ( .C ( clk ), .D ( signal_10645 ), .Q ( signal_10646 ) ) ;
    buf_clk cell_5062 ( .C ( clk ), .D ( signal_10653 ), .Q ( signal_10654 ) ) ;
    buf_clk cell_5070 ( .C ( clk ), .D ( signal_10661 ), .Q ( signal_10662 ) ) ;
    buf_clk cell_5078 ( .C ( clk ), .D ( signal_10669 ), .Q ( signal_10670 ) ) ;
    buf_clk cell_5086 ( .C ( clk ), .D ( signal_10677 ), .Q ( signal_10678 ) ) ;
    buf_clk cell_5094 ( .C ( clk ), .D ( signal_10685 ), .Q ( signal_10686 ) ) ;
    buf_clk cell_5098 ( .C ( clk ), .D ( signal_10689 ), .Q ( signal_10690 ) ) ;
    buf_clk cell_5102 ( .C ( clk ), .D ( signal_10693 ), .Q ( signal_10694 ) ) ;
    buf_clk cell_5106 ( .C ( clk ), .D ( signal_10697 ), .Q ( signal_10698 ) ) ;
    buf_clk cell_5110 ( .C ( clk ), .D ( signal_10701 ), .Q ( signal_10702 ) ) ;
    buf_clk cell_5114 ( .C ( clk ), .D ( signal_10705 ), .Q ( signal_10706 ) ) ;
    buf_clk cell_5118 ( .C ( clk ), .D ( signal_10709 ), .Q ( signal_10710 ) ) ;
    buf_clk cell_5134 ( .C ( clk ), .D ( signal_10725 ), .Q ( signal_10726 ) ) ;
    buf_clk cell_5138 ( .C ( clk ), .D ( signal_10729 ), .Q ( signal_10730 ) ) ;
    buf_clk cell_5142 ( .C ( clk ), .D ( signal_10733 ), .Q ( signal_10734 ) ) ;
    buf_clk cell_5152 ( .C ( clk ), .D ( signal_10743 ), .Q ( signal_10744 ) ) ;
    buf_clk cell_5162 ( .C ( clk ), .D ( signal_10753 ), .Q ( signal_10754 ) ) ;
    buf_clk cell_5172 ( .C ( clk ), .D ( signal_10763 ), .Q ( signal_10764 ) ) ;
    buf_clk cell_5178 ( .C ( clk ), .D ( signal_10769 ), .Q ( signal_10770 ) ) ;
    buf_clk cell_5184 ( .C ( clk ), .D ( signal_10775 ), .Q ( signal_10776 ) ) ;
    buf_clk cell_5190 ( .C ( clk ), .D ( signal_10781 ), .Q ( signal_10782 ) ) ;
    buf_clk cell_5204 ( .C ( clk ), .D ( signal_10795 ), .Q ( signal_10796 ) ) ;
    buf_clk cell_5212 ( .C ( clk ), .D ( signal_10803 ), .Q ( signal_10804 ) ) ;
    buf_clk cell_5220 ( .C ( clk ), .D ( signal_10811 ), .Q ( signal_10812 ) ) ;
    buf_clk cell_5226 ( .C ( clk ), .D ( signal_10817 ), .Q ( signal_10818 ) ) ;
    buf_clk cell_5232 ( .C ( clk ), .D ( signal_10823 ), .Q ( signal_10824 ) ) ;
    buf_clk cell_5238 ( .C ( clk ), .D ( signal_10829 ), .Q ( signal_10830 ) ) ;
    buf_clk cell_5246 ( .C ( clk ), .D ( signal_10837 ), .Q ( signal_10838 ) ) ;
    buf_clk cell_5254 ( .C ( clk ), .D ( signal_10845 ), .Q ( signal_10846 ) ) ;
    buf_clk cell_5262 ( .C ( clk ), .D ( signal_10853 ), .Q ( signal_10854 ) ) ;
    buf_clk cell_5270 ( .C ( clk ), .D ( signal_10861 ), .Q ( signal_10862 ) ) ;
    buf_clk cell_5278 ( .C ( clk ), .D ( signal_10869 ), .Q ( signal_10870 ) ) ;
    buf_clk cell_5286 ( .C ( clk ), .D ( signal_10877 ), .Q ( signal_10878 ) ) ;
    buf_clk cell_5294 ( .C ( clk ), .D ( signal_10885 ), .Q ( signal_10886 ) ) ;
    buf_clk cell_5302 ( .C ( clk ), .D ( signal_10893 ), .Q ( signal_10894 ) ) ;
    buf_clk cell_5310 ( .C ( clk ), .D ( signal_10901 ), .Q ( signal_10902 ) ) ;
    buf_clk cell_5320 ( .C ( clk ), .D ( signal_10911 ), .Q ( signal_10912 ) ) ;
    buf_clk cell_5330 ( .C ( clk ), .D ( signal_10921 ), .Q ( signal_10922 ) ) ;
    buf_clk cell_5340 ( .C ( clk ), .D ( signal_10931 ), .Q ( signal_10932 ) ) ;
    buf_clk cell_5348 ( .C ( clk ), .D ( signal_10939 ), .Q ( signal_10940 ) ) ;
    buf_clk cell_5356 ( .C ( clk ), .D ( signal_10947 ), .Q ( signal_10948 ) ) ;
    buf_clk cell_5364 ( .C ( clk ), .D ( signal_10955 ), .Q ( signal_10956 ) ) ;
    buf_clk cell_5372 ( .C ( clk ), .D ( signal_10963 ), .Q ( signal_10964 ) ) ;
    buf_clk cell_5380 ( .C ( clk ), .D ( signal_10971 ), .Q ( signal_10972 ) ) ;
    buf_clk cell_5388 ( .C ( clk ), .D ( signal_10979 ), .Q ( signal_10980 ) ) ;
    buf_clk cell_5402 ( .C ( clk ), .D ( signal_10993 ), .Q ( signal_10994 ) ) ;
    buf_clk cell_5410 ( .C ( clk ), .D ( signal_11001 ), .Q ( signal_11002 ) ) ;
    buf_clk cell_5418 ( .C ( clk ), .D ( signal_11009 ), .Q ( signal_11010 ) ) ;
    buf_clk cell_5426 ( .C ( clk ), .D ( signal_11017 ), .Q ( signal_11018 ) ) ;
    buf_clk cell_5434 ( .C ( clk ), .D ( signal_11025 ), .Q ( signal_11026 ) ) ;
    buf_clk cell_5442 ( .C ( clk ), .D ( signal_11033 ), .Q ( signal_11034 ) ) ;
    buf_clk cell_5450 ( .C ( clk ), .D ( signal_11041 ), .Q ( signal_11042 ) ) ;
    buf_clk cell_5458 ( .C ( clk ), .D ( signal_11049 ), .Q ( signal_11050 ) ) ;
    buf_clk cell_5466 ( .C ( clk ), .D ( signal_11057 ), .Q ( signal_11058 ) ) ;
    buf_clk cell_5470 ( .C ( clk ), .D ( signal_11061 ), .Q ( signal_11062 ) ) ;
    buf_clk cell_5476 ( .C ( clk ), .D ( signal_11067 ), .Q ( signal_11068 ) ) ;
    buf_clk cell_5482 ( .C ( clk ), .D ( signal_11073 ), .Q ( signal_11074 ) ) ;
    buf_clk cell_5490 ( .C ( clk ), .D ( signal_11081 ), .Q ( signal_11082 ) ) ;
    buf_clk cell_5498 ( .C ( clk ), .D ( signal_11089 ), .Q ( signal_11090 ) ) ;
    buf_clk cell_5506 ( .C ( clk ), .D ( signal_11097 ), .Q ( signal_11098 ) ) ;
    buf_clk cell_5512 ( .C ( clk ), .D ( signal_11103 ), .Q ( signal_11104 ) ) ;
    buf_clk cell_5518 ( .C ( clk ), .D ( signal_11109 ), .Q ( signal_11110 ) ) ;
    buf_clk cell_5524 ( .C ( clk ), .D ( signal_11115 ), .Q ( signal_11116 ) ) ;
    buf_clk cell_5530 ( .C ( clk ), .D ( signal_11121 ), .Q ( signal_11122 ) ) ;
    buf_clk cell_5536 ( .C ( clk ), .D ( signal_11127 ), .Q ( signal_11128 ) ) ;
    buf_clk cell_5542 ( .C ( clk ), .D ( signal_11133 ), .Q ( signal_11134 ) ) ;
    buf_clk cell_5550 ( .C ( clk ), .D ( signal_11141 ), .Q ( signal_11142 ) ) ;
    buf_clk cell_5558 ( .C ( clk ), .D ( signal_11149 ), .Q ( signal_11150 ) ) ;
    buf_clk cell_5566 ( .C ( clk ), .D ( signal_11157 ), .Q ( signal_11158 ) ) ;
    buf_clk cell_5576 ( .C ( clk ), .D ( signal_11167 ), .Q ( signal_11168 ) ) ;
    buf_clk cell_5586 ( .C ( clk ), .D ( signal_11177 ), .Q ( signal_11178 ) ) ;
    buf_clk cell_5596 ( .C ( clk ), .D ( signal_11187 ), .Q ( signal_11188 ) ) ;
    buf_clk cell_5608 ( .C ( clk ), .D ( signal_11199 ), .Q ( signal_11200 ) ) ;
    buf_clk cell_5614 ( .C ( clk ), .D ( signal_11205 ), .Q ( signal_11206 ) ) ;
    buf_clk cell_5620 ( .C ( clk ), .D ( signal_11211 ), .Q ( signal_11212 ) ) ;
    buf_clk cell_5628 ( .C ( clk ), .D ( signal_11219 ), .Q ( signal_11220 ) ) ;
    buf_clk cell_5636 ( .C ( clk ), .D ( signal_11227 ), .Q ( signal_11228 ) ) ;
    buf_clk cell_5644 ( .C ( clk ), .D ( signal_11235 ), .Q ( signal_11236 ) ) ;
    buf_clk cell_5654 ( .C ( clk ), .D ( signal_11245 ), .Q ( signal_11246 ) ) ;
    buf_clk cell_5664 ( .C ( clk ), .D ( signal_11255 ), .Q ( signal_11256 ) ) ;
    buf_clk cell_5674 ( .C ( clk ), .D ( signal_11265 ), .Q ( signal_11266 ) ) ;
    buf_clk cell_5682 ( .C ( clk ), .D ( signal_11273 ), .Q ( signal_11274 ) ) ;
    buf_clk cell_5690 ( .C ( clk ), .D ( signal_11281 ), .Q ( signal_11282 ) ) ;
    buf_clk cell_5698 ( .C ( clk ), .D ( signal_11289 ), .Q ( signal_11290 ) ) ;
    buf_clk cell_5704 ( .C ( clk ), .D ( signal_11295 ), .Q ( signal_11296 ) ) ;
    buf_clk cell_5710 ( .C ( clk ), .D ( signal_11301 ), .Q ( signal_11302 ) ) ;
    buf_clk cell_5716 ( .C ( clk ), .D ( signal_11307 ), .Q ( signal_11308 ) ) ;
    buf_clk cell_5722 ( .C ( clk ), .D ( signal_11313 ), .Q ( signal_11314 ) ) ;
    buf_clk cell_5728 ( .C ( clk ), .D ( signal_11319 ), .Q ( signal_11320 ) ) ;
    buf_clk cell_5734 ( .C ( clk ), .D ( signal_11325 ), .Q ( signal_11326 ) ) ;
    buf_clk cell_5770 ( .C ( clk ), .D ( signal_11361 ), .Q ( signal_11362 ) ) ;
    buf_clk cell_5776 ( .C ( clk ), .D ( signal_11367 ), .Q ( signal_11368 ) ) ;
    buf_clk cell_5782 ( .C ( clk ), .D ( signal_11373 ), .Q ( signal_11374 ) ) ;
    buf_clk cell_5794 ( .C ( clk ), .D ( signal_11385 ), .Q ( signal_11386 ) ) ;
    buf_clk cell_5800 ( .C ( clk ), .D ( signal_11391 ), .Q ( signal_11392 ) ) ;
    buf_clk cell_5806 ( .C ( clk ), .D ( signal_11397 ), .Q ( signal_11398 ) ) ;
    buf_clk cell_5824 ( .C ( clk ), .D ( signal_11415 ), .Q ( signal_11416 ) ) ;
    buf_clk cell_5830 ( .C ( clk ), .D ( signal_11421 ), .Q ( signal_11422 ) ) ;
    buf_clk cell_5836 ( .C ( clk ), .D ( signal_11427 ), .Q ( signal_11428 ) ) ;
    buf_clk cell_5878 ( .C ( clk ), .D ( signal_11469 ), .Q ( signal_11470 ) ) ;
    buf_clk cell_5886 ( .C ( clk ), .D ( signal_11477 ), .Q ( signal_11478 ) ) ;
    buf_clk cell_5894 ( .C ( clk ), .D ( signal_11485 ), .Q ( signal_11486 ) ) ;
    buf_clk cell_5922 ( .C ( clk ), .D ( signal_11513 ), .Q ( signal_11514 ) ) ;
    buf_clk cell_5932 ( .C ( clk ), .D ( signal_11523 ), .Q ( signal_11524 ) ) ;
    buf_clk cell_5942 ( .C ( clk ), .D ( signal_11533 ), .Q ( signal_11534 ) ) ;
    buf_clk cell_5980 ( .C ( clk ), .D ( signal_11571 ), .Q ( signal_11572 ) ) ;
    buf_clk cell_5988 ( .C ( clk ), .D ( signal_11579 ), .Q ( signal_11580 ) ) ;
    buf_clk cell_5996 ( .C ( clk ), .D ( signal_11587 ), .Q ( signal_11588 ) ) ;
    buf_clk cell_6022 ( .C ( clk ), .D ( signal_11613 ), .Q ( signal_11614 ) ) ;
    buf_clk cell_6030 ( .C ( clk ), .D ( signal_11621 ), .Q ( signal_11622 ) ) ;
    buf_clk cell_6038 ( .C ( clk ), .D ( signal_11629 ), .Q ( signal_11630 ) ) ;
    buf_clk cell_6064 ( .C ( clk ), .D ( signal_11655 ), .Q ( signal_11656 ) ) ;
    buf_clk cell_6072 ( .C ( clk ), .D ( signal_11663 ), .Q ( signal_11664 ) ) ;
    buf_clk cell_6080 ( .C ( clk ), .D ( signal_11671 ), .Q ( signal_11672 ) ) ;
    buf_clk cell_6186 ( .C ( clk ), .D ( signal_11777 ), .Q ( signal_11778 ) ) ;
    buf_clk cell_6198 ( .C ( clk ), .D ( signal_11789 ), .Q ( signal_11790 ) ) ;
    buf_clk cell_6210 ( .C ( clk ), .D ( signal_11801 ), .Q ( signal_11802 ) ) ;
    buf_clk cell_6260 ( .C ( clk ), .D ( signal_11851 ), .Q ( signal_11852 ) ) ;
    buf_clk cell_6274 ( .C ( clk ), .D ( signal_11865 ), .Q ( signal_11866 ) ) ;
    buf_clk cell_6288 ( .C ( clk ), .D ( signal_11879 ), .Q ( signal_11880 ) ) ;
    buf_clk cell_6326 ( .C ( clk ), .D ( signal_11917 ), .Q ( signal_11918 ) ) ;
    buf_clk cell_6340 ( .C ( clk ), .D ( signal_11931 ), .Q ( signal_11932 ) ) ;
    buf_clk cell_6354 ( .C ( clk ), .D ( signal_11945 ), .Q ( signal_11946 ) ) ;
    buf_clk cell_6446 ( .C ( clk ), .D ( signal_12037 ), .Q ( signal_12038 ) ) ;
    buf_clk cell_6462 ( .C ( clk ), .D ( signal_12053 ), .Q ( signal_12054 ) ) ;
    buf_clk cell_6478 ( .C ( clk ), .D ( signal_12069 ), .Q ( signal_12070 ) ) ;
    buf_clk cell_6506 ( .C ( clk ), .D ( signal_12097 ), .Q ( signal_12098 ) ) ;
    buf_clk cell_6522 ( .C ( clk ), .D ( signal_12113 ), .Q ( signal_12114 ) ) ;
    buf_clk cell_6538 ( .C ( clk ), .D ( signal_12129 ), .Q ( signal_12130 ) ) ;
    buf_clk cell_6690 ( .C ( clk ), .D ( signal_12281 ), .Q ( signal_12282 ) ) ;
    buf_clk cell_6706 ( .C ( clk ), .D ( signal_12297 ), .Q ( signal_12298 ) ) ;
    buf_clk cell_6722 ( .C ( clk ), .D ( signal_12313 ), .Q ( signal_12314 ) ) ;
    buf_clk cell_6740 ( .C ( clk ), .D ( signal_12331 ), .Q ( signal_12332 ) ) ;
    buf_clk cell_6758 ( .C ( clk ), .D ( signal_12349 ), .Q ( signal_12350 ) ) ;
    buf_clk cell_6776 ( .C ( clk ), .D ( signal_12367 ), .Q ( signal_12368 ) ) ;
    buf_clk cell_6890 ( .C ( clk ), .D ( signal_12481 ), .Q ( signal_12482 ) ) ;
    buf_clk cell_6910 ( .C ( clk ), .D ( signal_12501 ), .Q ( signal_12502 ) ) ;
    buf_clk cell_6930 ( .C ( clk ), .D ( signal_12521 ), .Q ( signal_12522 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_5009 ( .C ( clk ), .D ( signal_10600 ), .Q ( signal_10601 ) ) ;
    buf_clk cell_5019 ( .C ( clk ), .D ( signal_10610 ), .Q ( signal_10611 ) ) ;
    buf_clk cell_5029 ( .C ( clk ), .D ( signal_10620 ), .Q ( signal_10621 ) ) ;
    buf_clk cell_5035 ( .C ( clk ), .D ( signal_10626 ), .Q ( signal_10627 ) ) ;
    buf_clk cell_5041 ( .C ( clk ), .D ( signal_10632 ), .Q ( signal_10633 ) ) ;
    buf_clk cell_5047 ( .C ( clk ), .D ( signal_10638 ), .Q ( signal_10639 ) ) ;
    buf_clk cell_5055 ( .C ( clk ), .D ( signal_10646 ), .Q ( signal_10647 ) ) ;
    buf_clk cell_5063 ( .C ( clk ), .D ( signal_10654 ), .Q ( signal_10655 ) ) ;
    buf_clk cell_5071 ( .C ( clk ), .D ( signal_10662 ), .Q ( signal_10663 ) ) ;
    buf_clk cell_5079 ( .C ( clk ), .D ( signal_10670 ), .Q ( signal_10671 ) ) ;
    buf_clk cell_5087 ( .C ( clk ), .D ( signal_10678 ), .Q ( signal_10679 ) ) ;
    buf_clk cell_5095 ( .C ( clk ), .D ( signal_10686 ), .Q ( signal_10687 ) ) ;
    buf_clk cell_5099 ( .C ( clk ), .D ( signal_10690 ), .Q ( signal_10691 ) ) ;
    buf_clk cell_5103 ( .C ( clk ), .D ( signal_10694 ), .Q ( signal_10695 ) ) ;
    buf_clk cell_5107 ( .C ( clk ), .D ( signal_10698 ), .Q ( signal_10699 ) ) ;
    buf_clk cell_5111 ( .C ( clk ), .D ( signal_10702 ), .Q ( signal_10703 ) ) ;
    buf_clk cell_5115 ( .C ( clk ), .D ( signal_10706 ), .Q ( signal_10707 ) ) ;
    buf_clk cell_5119 ( .C ( clk ), .D ( signal_10710 ), .Q ( signal_10711 ) ) ;
    buf_clk cell_5121 ( .C ( clk ), .D ( signal_10540 ), .Q ( signal_10713 ) ) ;
    buf_clk cell_5123 ( .C ( clk ), .D ( signal_10542 ), .Q ( signal_10715 ) ) ;
    buf_clk cell_5125 ( .C ( clk ), .D ( signal_10544 ), .Q ( signal_10717 ) ) ;
    buf_clk cell_5127 ( .C ( clk ), .D ( signal_2156 ), .Q ( signal_10719 ) ) ;
    buf_clk cell_5129 ( .C ( clk ), .D ( signal_4836 ), .Q ( signal_10721 ) ) ;
    buf_clk cell_5131 ( .C ( clk ), .D ( signal_4837 ), .Q ( signal_10723 ) ) ;
    buf_clk cell_5135 ( .C ( clk ), .D ( signal_10726 ), .Q ( signal_10727 ) ) ;
    buf_clk cell_5139 ( .C ( clk ), .D ( signal_10730 ), .Q ( signal_10731 ) ) ;
    buf_clk cell_5143 ( .C ( clk ), .D ( signal_10734 ), .Q ( signal_10735 ) ) ;
    buf_clk cell_5153 ( .C ( clk ), .D ( signal_10744 ), .Q ( signal_10745 ) ) ;
    buf_clk cell_5163 ( .C ( clk ), .D ( signal_10754 ), .Q ( signal_10755 ) ) ;
    buf_clk cell_5173 ( .C ( clk ), .D ( signal_10764 ), .Q ( signal_10765 ) ) ;
    buf_clk cell_5179 ( .C ( clk ), .D ( signal_10770 ), .Q ( signal_10771 ) ) ;
    buf_clk cell_5185 ( .C ( clk ), .D ( signal_10776 ), .Q ( signal_10777 ) ) ;
    buf_clk cell_5191 ( .C ( clk ), .D ( signal_10782 ), .Q ( signal_10783 ) ) ;
    buf_clk cell_5193 ( .C ( clk ), .D ( signal_10290 ), .Q ( signal_10785 ) ) ;
    buf_clk cell_5195 ( .C ( clk ), .D ( signal_10294 ), .Q ( signal_10787 ) ) ;
    buf_clk cell_5197 ( .C ( clk ), .D ( signal_10298 ), .Q ( signal_10789 ) ) ;
    buf_clk cell_5205 ( .C ( clk ), .D ( signal_10796 ), .Q ( signal_10797 ) ) ;
    buf_clk cell_5213 ( .C ( clk ), .D ( signal_10804 ), .Q ( signal_10805 ) ) ;
    buf_clk cell_5221 ( .C ( clk ), .D ( signal_10812 ), .Q ( signal_10813 ) ) ;
    buf_clk cell_5227 ( .C ( clk ), .D ( signal_10818 ), .Q ( signal_10819 ) ) ;
    buf_clk cell_5233 ( .C ( clk ), .D ( signal_10824 ), .Q ( signal_10825 ) ) ;
    buf_clk cell_5239 ( .C ( clk ), .D ( signal_10830 ), .Q ( signal_10831 ) ) ;
    buf_clk cell_5247 ( .C ( clk ), .D ( signal_10838 ), .Q ( signal_10839 ) ) ;
    buf_clk cell_5255 ( .C ( clk ), .D ( signal_10846 ), .Q ( signal_10847 ) ) ;
    buf_clk cell_5263 ( .C ( clk ), .D ( signal_10854 ), .Q ( signal_10855 ) ) ;
    buf_clk cell_5271 ( .C ( clk ), .D ( signal_10862 ), .Q ( signal_10863 ) ) ;
    buf_clk cell_5279 ( .C ( clk ), .D ( signal_10870 ), .Q ( signal_10871 ) ) ;
    buf_clk cell_5287 ( .C ( clk ), .D ( signal_10878 ), .Q ( signal_10879 ) ) ;
    buf_clk cell_5295 ( .C ( clk ), .D ( signal_10886 ), .Q ( signal_10887 ) ) ;
    buf_clk cell_5303 ( .C ( clk ), .D ( signal_10894 ), .Q ( signal_10895 ) ) ;
    buf_clk cell_5311 ( .C ( clk ), .D ( signal_10902 ), .Q ( signal_10903 ) ) ;
    buf_clk cell_5321 ( .C ( clk ), .D ( signal_10912 ), .Q ( signal_10913 ) ) ;
    buf_clk cell_5331 ( .C ( clk ), .D ( signal_10922 ), .Q ( signal_10923 ) ) ;
    buf_clk cell_5341 ( .C ( clk ), .D ( signal_10932 ), .Q ( signal_10933 ) ) ;
    buf_clk cell_5349 ( .C ( clk ), .D ( signal_10940 ), .Q ( signal_10941 ) ) ;
    buf_clk cell_5357 ( .C ( clk ), .D ( signal_10948 ), .Q ( signal_10949 ) ) ;
    buf_clk cell_5365 ( .C ( clk ), .D ( signal_10956 ), .Q ( signal_10957 ) ) ;
    buf_clk cell_5373 ( .C ( clk ), .D ( signal_10964 ), .Q ( signal_10965 ) ) ;
    buf_clk cell_5381 ( .C ( clk ), .D ( signal_10972 ), .Q ( signal_10973 ) ) ;
    buf_clk cell_5389 ( .C ( clk ), .D ( signal_10980 ), .Q ( signal_10981 ) ) ;
    buf_clk cell_5391 ( .C ( clk ), .D ( signal_10222 ), .Q ( signal_10983 ) ) ;
    buf_clk cell_5393 ( .C ( clk ), .D ( signal_10224 ), .Q ( signal_10985 ) ) ;
    buf_clk cell_5395 ( .C ( clk ), .D ( signal_10226 ), .Q ( signal_10987 ) ) ;
    buf_clk cell_5403 ( .C ( clk ), .D ( signal_10994 ), .Q ( signal_10995 ) ) ;
    buf_clk cell_5411 ( .C ( clk ), .D ( signal_11002 ), .Q ( signal_11003 ) ) ;
    buf_clk cell_5419 ( .C ( clk ), .D ( signal_11010 ), .Q ( signal_11011 ) ) ;
    buf_clk cell_5427 ( .C ( clk ), .D ( signal_11018 ), .Q ( signal_11019 ) ) ;
    buf_clk cell_5435 ( .C ( clk ), .D ( signal_11026 ), .Q ( signal_11027 ) ) ;
    buf_clk cell_5443 ( .C ( clk ), .D ( signal_11034 ), .Q ( signal_11035 ) ) ;
    buf_clk cell_5451 ( .C ( clk ), .D ( signal_11042 ), .Q ( signal_11043 ) ) ;
    buf_clk cell_5459 ( .C ( clk ), .D ( signal_11050 ), .Q ( signal_11051 ) ) ;
    buf_clk cell_5467 ( .C ( clk ), .D ( signal_11058 ), .Q ( signal_11059 ) ) ;
    buf_clk cell_5471 ( .C ( clk ), .D ( signal_11062 ), .Q ( signal_11063 ) ) ;
    buf_clk cell_5477 ( .C ( clk ), .D ( signal_11068 ), .Q ( signal_11069 ) ) ;
    buf_clk cell_5483 ( .C ( clk ), .D ( signal_11074 ), .Q ( signal_11075 ) ) ;
    buf_clk cell_5491 ( .C ( clk ), .D ( signal_11082 ), .Q ( signal_11083 ) ) ;
    buf_clk cell_5499 ( .C ( clk ), .D ( signal_11090 ), .Q ( signal_11091 ) ) ;
    buf_clk cell_5507 ( .C ( clk ), .D ( signal_11098 ), .Q ( signal_11099 ) ) ;
    buf_clk cell_5513 ( .C ( clk ), .D ( signal_11104 ), .Q ( signal_11105 ) ) ;
    buf_clk cell_5519 ( .C ( clk ), .D ( signal_11110 ), .Q ( signal_11111 ) ) ;
    buf_clk cell_5525 ( .C ( clk ), .D ( signal_11116 ), .Q ( signal_11117 ) ) ;
    buf_clk cell_5531 ( .C ( clk ), .D ( signal_11122 ), .Q ( signal_11123 ) ) ;
    buf_clk cell_5537 ( .C ( clk ), .D ( signal_11128 ), .Q ( signal_11129 ) ) ;
    buf_clk cell_5543 ( .C ( clk ), .D ( signal_11134 ), .Q ( signal_11135 ) ) ;
    buf_clk cell_5551 ( .C ( clk ), .D ( signal_11142 ), .Q ( signal_11143 ) ) ;
    buf_clk cell_5559 ( .C ( clk ), .D ( signal_11150 ), .Q ( signal_11151 ) ) ;
    buf_clk cell_5567 ( .C ( clk ), .D ( signal_11158 ), .Q ( signal_11159 ) ) ;
    buf_clk cell_5577 ( .C ( clk ), .D ( signal_11168 ), .Q ( signal_11169 ) ) ;
    buf_clk cell_5587 ( .C ( clk ), .D ( signal_11178 ), .Q ( signal_11179 ) ) ;
    buf_clk cell_5597 ( .C ( clk ), .D ( signal_11188 ), .Q ( signal_11189 ) ) ;
    buf_clk cell_5609 ( .C ( clk ), .D ( signal_11200 ), .Q ( signal_11201 ) ) ;
    buf_clk cell_5615 ( .C ( clk ), .D ( signal_11206 ), .Q ( signal_11207 ) ) ;
    buf_clk cell_5621 ( .C ( clk ), .D ( signal_11212 ), .Q ( signal_11213 ) ) ;
    buf_clk cell_5629 ( .C ( clk ), .D ( signal_11220 ), .Q ( signal_11221 ) ) ;
    buf_clk cell_5637 ( .C ( clk ), .D ( signal_11228 ), .Q ( signal_11229 ) ) ;
    buf_clk cell_5645 ( .C ( clk ), .D ( signal_11236 ), .Q ( signal_11237 ) ) ;
    buf_clk cell_5655 ( .C ( clk ), .D ( signal_11246 ), .Q ( signal_11247 ) ) ;
    buf_clk cell_5665 ( .C ( clk ), .D ( signal_11256 ), .Q ( signal_11257 ) ) ;
    buf_clk cell_5675 ( .C ( clk ), .D ( signal_11266 ), .Q ( signal_11267 ) ) ;
    buf_clk cell_5683 ( .C ( clk ), .D ( signal_11274 ), .Q ( signal_11275 ) ) ;
    buf_clk cell_5691 ( .C ( clk ), .D ( signal_11282 ), .Q ( signal_11283 ) ) ;
    buf_clk cell_5699 ( .C ( clk ), .D ( signal_11290 ), .Q ( signal_11291 ) ) ;
    buf_clk cell_5705 ( .C ( clk ), .D ( signal_11296 ), .Q ( signal_11297 ) ) ;
    buf_clk cell_5711 ( .C ( clk ), .D ( signal_11302 ), .Q ( signal_11303 ) ) ;
    buf_clk cell_5717 ( .C ( clk ), .D ( signal_11308 ), .Q ( signal_11309 ) ) ;
    buf_clk cell_5723 ( .C ( clk ), .D ( signal_11314 ), .Q ( signal_11315 ) ) ;
    buf_clk cell_5729 ( .C ( clk ), .D ( signal_11320 ), .Q ( signal_11321 ) ) ;
    buf_clk cell_5735 ( .C ( clk ), .D ( signal_11326 ), .Q ( signal_11327 ) ) ;
    buf_clk cell_5745 ( .C ( clk ), .D ( signal_10490 ), .Q ( signal_11337 ) ) ;
    buf_clk cell_5749 ( .C ( clk ), .D ( signal_10496 ), .Q ( signal_11341 ) ) ;
    buf_clk cell_5753 ( .C ( clk ), .D ( signal_10502 ), .Q ( signal_11345 ) ) ;
    buf_clk cell_5757 ( .C ( clk ), .D ( signal_2253 ), .Q ( signal_11349 ) ) ;
    buf_clk cell_5761 ( .C ( clk ), .D ( signal_5030 ), .Q ( signal_11353 ) ) ;
    buf_clk cell_5765 ( .C ( clk ), .D ( signal_5031 ), .Q ( signal_11357 ) ) ;
    buf_clk cell_5771 ( .C ( clk ), .D ( signal_11362 ), .Q ( signal_11363 ) ) ;
    buf_clk cell_5777 ( .C ( clk ), .D ( signal_11368 ), .Q ( signal_11369 ) ) ;
    buf_clk cell_5783 ( .C ( clk ), .D ( signal_11374 ), .Q ( signal_11375 ) ) ;
    buf_clk cell_5795 ( .C ( clk ), .D ( signal_11386 ), .Q ( signal_11387 ) ) ;
    buf_clk cell_5801 ( .C ( clk ), .D ( signal_11392 ), .Q ( signal_11393 ) ) ;
    buf_clk cell_5807 ( .C ( clk ), .D ( signal_11398 ), .Q ( signal_11399 ) ) ;
    buf_clk cell_5811 ( .C ( clk ), .D ( signal_2208 ), .Q ( signal_11403 ) ) ;
    buf_clk cell_5815 ( .C ( clk ), .D ( signal_4940 ), .Q ( signal_11407 ) ) ;
    buf_clk cell_5819 ( .C ( clk ), .D ( signal_4941 ), .Q ( signal_11411 ) ) ;
    buf_clk cell_5825 ( .C ( clk ), .D ( signal_11416 ), .Q ( signal_11417 ) ) ;
    buf_clk cell_5831 ( .C ( clk ), .D ( signal_11422 ), .Q ( signal_11423 ) ) ;
    buf_clk cell_5837 ( .C ( clk ), .D ( signal_11428 ), .Q ( signal_11429 ) ) ;
    buf_clk cell_5847 ( .C ( clk ), .D ( signal_2249 ), .Q ( signal_11439 ) ) ;
    buf_clk cell_5851 ( .C ( clk ), .D ( signal_5022 ), .Q ( signal_11443 ) ) ;
    buf_clk cell_5855 ( .C ( clk ), .D ( signal_5023 ), .Q ( signal_11447 ) ) ;
    buf_clk cell_5859 ( .C ( clk ), .D ( signal_2161 ), .Q ( signal_11451 ) ) ;
    buf_clk cell_5865 ( .C ( clk ), .D ( signal_4846 ), .Q ( signal_11457 ) ) ;
    buf_clk cell_5871 ( .C ( clk ), .D ( signal_4847 ), .Q ( signal_11463 ) ) ;
    buf_clk cell_5879 ( .C ( clk ), .D ( signal_11470 ), .Q ( signal_11471 ) ) ;
    buf_clk cell_5887 ( .C ( clk ), .D ( signal_11478 ), .Q ( signal_11479 ) ) ;
    buf_clk cell_5895 ( .C ( clk ), .D ( signal_11486 ), .Q ( signal_11487 ) ) ;
    buf_clk cell_5901 ( .C ( clk ), .D ( signal_2199 ), .Q ( signal_11493 ) ) ;
    buf_clk cell_5907 ( .C ( clk ), .D ( signal_4922 ), .Q ( signal_11499 ) ) ;
    buf_clk cell_5913 ( .C ( clk ), .D ( signal_4923 ), .Q ( signal_11505 ) ) ;
    buf_clk cell_5923 ( .C ( clk ), .D ( signal_11514 ), .Q ( signal_11515 ) ) ;
    buf_clk cell_5933 ( .C ( clk ), .D ( signal_11524 ), .Q ( signal_11525 ) ) ;
    buf_clk cell_5943 ( .C ( clk ), .D ( signal_11534 ), .Q ( signal_11535 ) ) ;
    buf_clk cell_5949 ( .C ( clk ), .D ( signal_2255 ), .Q ( signal_11541 ) ) ;
    buf_clk cell_5955 ( .C ( clk ), .D ( signal_5034 ), .Q ( signal_11547 ) ) ;
    buf_clk cell_5961 ( .C ( clk ), .D ( signal_5035 ), .Q ( signal_11553 ) ) ;
    buf_clk cell_5981 ( .C ( clk ), .D ( signal_11572 ), .Q ( signal_11573 ) ) ;
    buf_clk cell_5989 ( .C ( clk ), .D ( signal_11580 ), .Q ( signal_11581 ) ) ;
    buf_clk cell_5997 ( .C ( clk ), .D ( signal_11588 ), .Q ( signal_11589 ) ) ;
    buf_clk cell_6003 ( .C ( clk ), .D ( signal_2183 ), .Q ( signal_11595 ) ) ;
    buf_clk cell_6009 ( .C ( clk ), .D ( signal_4890 ), .Q ( signal_11601 ) ) ;
    buf_clk cell_6015 ( .C ( clk ), .D ( signal_4891 ), .Q ( signal_11607 ) ) ;
    buf_clk cell_6023 ( .C ( clk ), .D ( signal_11614 ), .Q ( signal_11615 ) ) ;
    buf_clk cell_6031 ( .C ( clk ), .D ( signal_11622 ), .Q ( signal_11623 ) ) ;
    buf_clk cell_6039 ( .C ( clk ), .D ( signal_11630 ), .Q ( signal_11631 ) ) ;
    buf_clk cell_6045 ( .C ( clk ), .D ( signal_10534 ), .Q ( signal_11637 ) ) ;
    buf_clk cell_6051 ( .C ( clk ), .D ( signal_10536 ), .Q ( signal_11643 ) ) ;
    buf_clk cell_6057 ( .C ( clk ), .D ( signal_10538 ), .Q ( signal_11649 ) ) ;
    buf_clk cell_6065 ( .C ( clk ), .D ( signal_11656 ), .Q ( signal_11657 ) ) ;
    buf_clk cell_6073 ( .C ( clk ), .D ( signal_11664 ), .Q ( signal_11665 ) ) ;
    buf_clk cell_6081 ( .C ( clk ), .D ( signal_11672 ), .Q ( signal_11673 ) ) ;
    buf_clk cell_6099 ( .C ( clk ), .D ( signal_2252 ), .Q ( signal_11691 ) ) ;
    buf_clk cell_6105 ( .C ( clk ), .D ( signal_5028 ), .Q ( signal_11697 ) ) ;
    buf_clk cell_6111 ( .C ( clk ), .D ( signal_5029 ), .Q ( signal_11703 ) ) ;
    buf_clk cell_6117 ( .C ( clk ), .D ( signal_2160 ), .Q ( signal_11709 ) ) ;
    buf_clk cell_6123 ( .C ( clk ), .D ( signal_4844 ), .Q ( signal_11715 ) ) ;
    buf_clk cell_6129 ( .C ( clk ), .D ( signal_4845 ), .Q ( signal_11721 ) ) ;
    buf_clk cell_6159 ( .C ( clk ), .D ( signal_2202 ), .Q ( signal_11751 ) ) ;
    buf_clk cell_6167 ( .C ( clk ), .D ( signal_4928 ), .Q ( signal_11759 ) ) ;
    buf_clk cell_6175 ( .C ( clk ), .D ( signal_4929 ), .Q ( signal_11767 ) ) ;
    buf_clk cell_6187 ( .C ( clk ), .D ( signal_11778 ), .Q ( signal_11779 ) ) ;
    buf_clk cell_6199 ( .C ( clk ), .D ( signal_11790 ), .Q ( signal_11791 ) ) ;
    buf_clk cell_6211 ( .C ( clk ), .D ( signal_11802 ), .Q ( signal_11803 ) ) ;
    buf_clk cell_6261 ( .C ( clk ), .D ( signal_11852 ), .Q ( signal_11853 ) ) ;
    buf_clk cell_6275 ( .C ( clk ), .D ( signal_11866 ), .Q ( signal_11867 ) ) ;
    buf_clk cell_6289 ( .C ( clk ), .D ( signal_11880 ), .Q ( signal_11881 ) ) ;
    buf_clk cell_6297 ( .C ( clk ), .D ( signal_2154 ), .Q ( signal_11889 ) ) ;
    buf_clk cell_6305 ( .C ( clk ), .D ( signal_4832 ), .Q ( signal_11897 ) ) ;
    buf_clk cell_6313 ( .C ( clk ), .D ( signal_4833 ), .Q ( signal_11905 ) ) ;
    buf_clk cell_6327 ( .C ( clk ), .D ( signal_11918 ), .Q ( signal_11919 ) ) ;
    buf_clk cell_6341 ( .C ( clk ), .D ( signal_11932 ), .Q ( signal_11933 ) ) ;
    buf_clk cell_6355 ( .C ( clk ), .D ( signal_11946 ), .Q ( signal_11947 ) ) ;
    buf_clk cell_6363 ( .C ( clk ), .D ( signal_2149 ), .Q ( signal_11955 ) ) ;
    buf_clk cell_6371 ( .C ( clk ), .D ( signal_4822 ), .Q ( signal_11963 ) ) ;
    buf_clk cell_6379 ( .C ( clk ), .D ( signal_4823 ), .Q ( signal_11971 ) ) ;
    buf_clk cell_6399 ( .C ( clk ), .D ( signal_2152 ), .Q ( signal_11991 ) ) ;
    buf_clk cell_6409 ( .C ( clk ), .D ( signal_4828 ), .Q ( signal_12001 ) ) ;
    buf_clk cell_6419 ( .C ( clk ), .D ( signal_4829 ), .Q ( signal_12011 ) ) ;
    buf_clk cell_6447 ( .C ( clk ), .D ( signal_12038 ), .Q ( signal_12039 ) ) ;
    buf_clk cell_6463 ( .C ( clk ), .D ( signal_12054 ), .Q ( signal_12055 ) ) ;
    buf_clk cell_6479 ( .C ( clk ), .D ( signal_12070 ), .Q ( signal_12071 ) ) ;
    buf_clk cell_6507 ( .C ( clk ), .D ( signal_12098 ), .Q ( signal_12099 ) ) ;
    buf_clk cell_6523 ( .C ( clk ), .D ( signal_12114 ), .Q ( signal_12115 ) ) ;
    buf_clk cell_6539 ( .C ( clk ), .D ( signal_12130 ), .Q ( signal_12131 ) ) ;
    buf_clk cell_6549 ( .C ( clk ), .D ( signal_2257 ), .Q ( signal_12141 ) ) ;
    buf_clk cell_6559 ( .C ( clk ), .D ( signal_5038 ), .Q ( signal_12151 ) ) ;
    buf_clk cell_6569 ( .C ( clk ), .D ( signal_5039 ), .Q ( signal_12161 ) ) ;
    buf_clk cell_6691 ( .C ( clk ), .D ( signal_12282 ), .Q ( signal_12283 ) ) ;
    buf_clk cell_6707 ( .C ( clk ), .D ( signal_12298 ), .Q ( signal_12299 ) ) ;
    buf_clk cell_6723 ( .C ( clk ), .D ( signal_12314 ), .Q ( signal_12315 ) ) ;
    buf_clk cell_6741 ( .C ( clk ), .D ( signal_12332 ), .Q ( signal_12333 ) ) ;
    buf_clk cell_6759 ( .C ( clk ), .D ( signal_12350 ), .Q ( signal_12351 ) ) ;
    buf_clk cell_6777 ( .C ( clk ), .D ( signal_12368 ), .Q ( signal_12369 ) ) ;
    buf_clk cell_6891 ( .C ( clk ), .D ( signal_12482 ), .Q ( signal_12483 ) ) ;
    buf_clk cell_6911 ( .C ( clk ), .D ( signal_12502 ), .Q ( signal_12503 ) ) ;
    buf_clk cell_6931 ( .C ( clk ), .D ( signal_12522 ), .Q ( signal_12523 ) ) ;

    /* cells in depth 14 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2116 ( .a ({signal_10112, signal_10104, signal_10096}), .b ({signal_4631, signal_4630, signal_2053}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187]}), .c ({signal_4787, signal_4786, signal_2131}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2118 ( .a ({signal_10124, signal_10120, signal_10116}), .b ({signal_4633, signal_4632, signal_2054}), .clk ( clk ), .r ({Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_4791, signal_4790, signal_2133}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2119 ( .a ({signal_10142, signal_10136, signal_10130}), .b ({signal_4635, signal_4634, signal_2055}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193]}), .c ({signal_4793, signal_4792, signal_2134}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2121 ( .a ({signal_10160, signal_10154, signal_10148}), .b ({signal_4639, signal_4638, signal_2057}), .clk ( clk ), .r ({Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({signal_4797, signal_4796, signal_2136}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2122 ( .a ({signal_10172, signal_10168, signal_10164}), .b ({signal_4643, signal_4642, signal_2059}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199]}), .c ({signal_4799, signal_4798, signal_2137}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2123 ( .a ({signal_10190, signal_10184, signal_10178}), .b ({signal_4645, signal_4644, signal_2060}), .clk ( clk ), .r ({Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({signal_4801, signal_4800, signal_2138}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2140 ( .a ({signal_4793, signal_4792, signal_2134}), .b ({signal_4835, signal_4834, signal_2155}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2162 ( .a ({signal_10202, signal_10198, signal_10194}), .b ({signal_4683, signal_4682, signal_2079}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205]}), .c ({signal_4879, signal_4878, signal_2177}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2170 ( .a ({signal_10214, signal_10210, signal_10206}), .b ({signal_4751, signal_4750, signal_2113}), .clk ( clk ), .r ({Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({signal_4895, signal_4894, signal_2185}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2172 ( .a ({signal_10220, signal_10218, signal_10216}), .b ({signal_4759, signal_4758, signal_2117}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211]}), .c ({signal_4899, signal_4898, signal_2187}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2173 ( .a ({signal_10226, signal_10224, signal_10222}), .b ({signal_4699, signal_4698, signal_2087}), .clk ( clk ), .r ({Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({signal_4901, signal_4900, signal_2188}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2174 ( .a ({signal_10244, signal_10238, signal_10232}), .b ({signal_4767, signal_4766, signal_2121}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217]}), .c ({signal_4903, signal_4902, signal_2189}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2175 ( .a ({signal_10262, signal_10256, signal_10250}), .b ({signal_4769, signal_4768, signal_2122}), .clk ( clk ), .r ({Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_4905, signal_4904, signal_2190}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2176 ( .a ({signal_10280, signal_10274, signal_10268}), .b ({signal_4771, signal_4770, signal_2123}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223]}), .c ({signal_4907, signal_4906, signal_2191}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2177 ( .a ({signal_4691, signal_4690, signal_2083}), .b ({signal_4637, signal_4636, signal_2056}), .clk ( clk ), .r ({Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({signal_4909, signal_4908, signal_2192}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2178 ( .a ({signal_10286, signal_10284, signal_10282}), .b ({signal_4701, signal_4700, signal_2088}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229]}), .c ({signal_4911, signal_4910, signal_2193}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2179 ( .a ({signal_10298, signal_10294, signal_10290}), .b ({signal_4781, signal_4780, signal_2128}), .clk ( clk ), .r ({Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({signal_4913, signal_4912, signal_2194}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2190 ( .a ({signal_4879, signal_4878, signal_2177}), .b ({signal_4935, signal_4934, signal_2205}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2195 ( .a ({signal_4901, signal_4900, signal_2188}), .b ({signal_4945, signal_4944, signal_2210}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2196 ( .a ({signal_4905, signal_4904, signal_2190}), .b ({signal_4947, signal_4946, signal_2211}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2197 ( .a ({signal_4907, signal_4906, signal_2191}), .b ({signal_4949, signal_4948, signal_2212}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2198 ( .a ({signal_4911, signal_4910, signal_2193}), .b ({signal_4951, signal_4950, signal_2213}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2200 ( .a ({signal_10316, signal_10310, signal_10304}), .b ({signal_4839, signal_4838, signal_2157}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235]}), .c ({signal_4955, signal_4954, signal_2215}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2207 ( .a ({signal_10322, signal_10320, signal_10318}), .b ({signal_4817, signal_4816, signal_2146}), .clk ( clk ), .r ({Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({signal_4969, signal_4968, signal_2222}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2208 ( .a ({signal_10340, signal_10334, signal_10328}), .b ({signal_4853, signal_4852, signal_2164}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241]}), .c ({signal_4971, signal_4970, signal_2223}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2209 ( .a ({signal_10346, signal_10344, signal_10342}), .b ({signal_4819, signal_4818, signal_2147}), .clk ( clk ), .r ({Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({signal_4973, signal_4972, signal_2224}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2210 ( .a ({signal_10370, signal_10362, signal_10354}), .b ({signal_4855, signal_4854, signal_2165}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247]}), .c ({signal_4975, signal_4974, signal_2225}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2211 ( .a ({signal_10382, signal_10378, signal_10374}), .b ({signal_4859, signal_4858, signal_2167}), .clk ( clk ), .r ({Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_4977, signal_4976, signal_2226}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2212 ( .a ({signal_4761, signal_4760, signal_2118}), .b ({signal_4861, signal_4860, signal_2168}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253]}), .c ({signal_4979, signal_4978, signal_2227}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2214 ( .a ({signal_10394, signal_10390, signal_10386}), .b ({signal_4863, signal_4862, signal_2169}), .clk ( clk ), .r ({Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({signal_4983, signal_4982, signal_2229}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2215 ( .a ({signal_4765, signal_4764, signal_2120}), .b ({signal_4865, signal_4864, signal_2170}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259]}), .c ({signal_4985, signal_4984, signal_2230}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2216 ( .a ({signal_10412, signal_10406, signal_10400}), .b ({signal_4867, signal_4866, signal_2171}), .clk ( clk ), .r ({Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({signal_4987, signal_4986, signal_2231}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2217 ( .a ({signal_10430, signal_10424, signal_10418}), .b ({signal_4871, signal_4870, signal_2173}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265]}), .c ({signal_4989, signal_4988, signal_2232}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2218 ( .a ({signal_10442, signal_10438, signal_10434}), .b ({signal_4875, signal_4874, signal_2175}), .clk ( clk ), .r ({Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({signal_4991, signal_4990, signal_2233}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2219 ( .a ({signal_10466, signal_10458, signal_10450}), .b ({signal_4877, signal_4876, signal_2176}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271]}), .c ({signal_4993, signal_4992, signal_2234}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2220 ( .a ({signal_10484, signal_10478, signal_10472}), .b ({signal_4881, signal_4880, signal_2178}), .clk ( clk ), .r ({Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({signal_4995, signal_4994, signal_2235}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2222 ( .a ({signal_4827, signal_4826, signal_2151}), .b ({signal_4779, signal_4778, signal_2127}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277]}), .c ({signal_4999, signal_4998, signal_2237}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2223 ( .a ({signal_4831, signal_4830, signal_2153}), .b ({signal_4889, signal_4888, signal_2182}), .clk ( clk ), .r ({Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_5001, signal_5000, signal_2238}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2224 ( .a ({signal_10502, signal_10496, signal_10490}), .b ({signal_4893, signal_4892, signal_2184}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283]}), .c ({signal_5003, signal_5002, signal_2239}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2239 ( .a ({signal_4971, signal_4970, signal_2223}), .b ({signal_5033, signal_5032, signal_2254}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2241 ( .a ({signal_4989, signal_4988, signal_2232}), .b ({signal_5037, signal_5036, signal_2256}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2243 ( .a ({signal_5003, signal_5002, signal_2239}), .b ({signal_5041, signal_5040, signal_2258}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2249 ( .a ({signal_4849, signal_4848, signal_2162}), .b ({signal_10508, signal_10506, signal_10504}), .clk ( clk ), .r ({Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({signal_5053, signal_5052, signal_2264}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2250 ( .a ({signal_4813, signal_4812, signal_2144}), .b ({signal_4931, signal_4930, signal_2203}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289]}), .c ({signal_5055, signal_5054, signal_2265}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2251 ( .a ({signal_10514, signal_10512, signal_10510}), .b ({signal_4933, signal_4932, signal_2204}), .clk ( clk ), .r ({Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({signal_5057, signal_5056, signal_2266}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2252 ( .a ({signal_10532, signal_10526, signal_10520}), .b ({signal_4937, signal_4936, signal_2206}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295]}), .c ({signal_5059, signal_5058, signal_2267}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2253 ( .a ({signal_10538, signal_10536, signal_10534}), .b ({signal_4939, signal_4938, signal_2207}), .clk ( clk ), .r ({Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({signal_5061, signal_5060, signal_2268}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2254 ( .a ({signal_10544, signal_10542, signal_10540}), .b ({signal_4943, signal_4942, signal_2209}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301]}), .c ({signal_5063, signal_5062, signal_2269}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2271 ( .a ({signal_5057, signal_5056, signal_2266}), .b ({signal_5097, signal_5096, signal_2286}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2272 ( .a ({signal_5059, signal_5058, signal_2267}), .b ({signal_5099, signal_5098, signal_2287}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2273 ( .a ({signal_5061, signal_5060, signal_2268}), .b ({signal_5101, signal_5100, signal_2288}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2274 ( .a ({signal_5063, signal_5062, signal_2269}), .b ({signal_5103, signal_5102, signal_2289}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2282 ( .a ({signal_5025, signal_5024, signal_2250}), .b ({signal_10562, signal_10556, signal_10550}), .clk ( clk ), .r ({Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({signal_5119, signal_5118, signal_2297}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2283 ( .a ({signal_10538, signal_10536, signal_10534}), .b ({signal_5021, signal_5020, signal_2248}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307]}), .c ({signal_5121, signal_5120, signal_2298}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2285 ( .a ({signal_10580, signal_10574, signal_10568}), .b ({signal_5051, signal_5050, signal_2263}), .clk ( clk ), .r ({Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_5125, signal_5124, signal_2300}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2286 ( .a ({signal_10592, signal_10588, signal_10584}), .b ({signal_5027, signal_5026, signal_2251}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313]}), .c ({signal_5127, signal_5126, signal_2301}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2297 ( .a ({signal_5121, signal_5120, signal_2298}), .b ({signal_5149, signal_5148, signal_2312}) ) ;
    buf_clk cell_5010 ( .C ( clk ), .D ( signal_10601 ), .Q ( signal_10602 ) ) ;
    buf_clk cell_5020 ( .C ( clk ), .D ( signal_10611 ), .Q ( signal_10612 ) ) ;
    buf_clk cell_5030 ( .C ( clk ), .D ( signal_10621 ), .Q ( signal_10622 ) ) ;
    buf_clk cell_5036 ( .C ( clk ), .D ( signal_10627 ), .Q ( signal_10628 ) ) ;
    buf_clk cell_5042 ( .C ( clk ), .D ( signal_10633 ), .Q ( signal_10634 ) ) ;
    buf_clk cell_5048 ( .C ( clk ), .D ( signal_10639 ), .Q ( signal_10640 ) ) ;
    buf_clk cell_5056 ( .C ( clk ), .D ( signal_10647 ), .Q ( signal_10648 ) ) ;
    buf_clk cell_5064 ( .C ( clk ), .D ( signal_10655 ), .Q ( signal_10656 ) ) ;
    buf_clk cell_5072 ( .C ( clk ), .D ( signal_10663 ), .Q ( signal_10664 ) ) ;
    buf_clk cell_5080 ( .C ( clk ), .D ( signal_10671 ), .Q ( signal_10672 ) ) ;
    buf_clk cell_5088 ( .C ( clk ), .D ( signal_10679 ), .Q ( signal_10680 ) ) ;
    buf_clk cell_5096 ( .C ( clk ), .D ( signal_10687 ), .Q ( signal_10688 ) ) ;
    buf_clk cell_5100 ( .C ( clk ), .D ( signal_10691 ), .Q ( signal_10692 ) ) ;
    buf_clk cell_5104 ( .C ( clk ), .D ( signal_10695 ), .Q ( signal_10696 ) ) ;
    buf_clk cell_5108 ( .C ( clk ), .D ( signal_10699 ), .Q ( signal_10700 ) ) ;
    buf_clk cell_5112 ( .C ( clk ), .D ( signal_10703 ), .Q ( signal_10704 ) ) ;
    buf_clk cell_5116 ( .C ( clk ), .D ( signal_10707 ), .Q ( signal_10708 ) ) ;
    buf_clk cell_5120 ( .C ( clk ), .D ( signal_10711 ), .Q ( signal_10712 ) ) ;
    buf_clk cell_5122 ( .C ( clk ), .D ( signal_10713 ), .Q ( signal_10714 ) ) ;
    buf_clk cell_5124 ( .C ( clk ), .D ( signal_10715 ), .Q ( signal_10716 ) ) ;
    buf_clk cell_5126 ( .C ( clk ), .D ( signal_10717 ), .Q ( signal_10718 ) ) ;
    buf_clk cell_5128 ( .C ( clk ), .D ( signal_10719 ), .Q ( signal_10720 ) ) ;
    buf_clk cell_5130 ( .C ( clk ), .D ( signal_10721 ), .Q ( signal_10722 ) ) ;
    buf_clk cell_5132 ( .C ( clk ), .D ( signal_10723 ), .Q ( signal_10724 ) ) ;
    buf_clk cell_5136 ( .C ( clk ), .D ( signal_10727 ), .Q ( signal_10728 ) ) ;
    buf_clk cell_5140 ( .C ( clk ), .D ( signal_10731 ), .Q ( signal_10732 ) ) ;
    buf_clk cell_5144 ( .C ( clk ), .D ( signal_10735 ), .Q ( signal_10736 ) ) ;
    buf_clk cell_5154 ( .C ( clk ), .D ( signal_10745 ), .Q ( signal_10746 ) ) ;
    buf_clk cell_5164 ( .C ( clk ), .D ( signal_10755 ), .Q ( signal_10756 ) ) ;
    buf_clk cell_5174 ( .C ( clk ), .D ( signal_10765 ), .Q ( signal_10766 ) ) ;
    buf_clk cell_5180 ( .C ( clk ), .D ( signal_10771 ), .Q ( signal_10772 ) ) ;
    buf_clk cell_5186 ( .C ( clk ), .D ( signal_10777 ), .Q ( signal_10778 ) ) ;
    buf_clk cell_5192 ( .C ( clk ), .D ( signal_10783 ), .Q ( signal_10784 ) ) ;
    buf_clk cell_5194 ( .C ( clk ), .D ( signal_10785 ), .Q ( signal_10786 ) ) ;
    buf_clk cell_5196 ( .C ( clk ), .D ( signal_10787 ), .Q ( signal_10788 ) ) ;
    buf_clk cell_5198 ( .C ( clk ), .D ( signal_10789 ), .Q ( signal_10790 ) ) ;
    buf_clk cell_5206 ( .C ( clk ), .D ( signal_10797 ), .Q ( signal_10798 ) ) ;
    buf_clk cell_5214 ( .C ( clk ), .D ( signal_10805 ), .Q ( signal_10806 ) ) ;
    buf_clk cell_5222 ( .C ( clk ), .D ( signal_10813 ), .Q ( signal_10814 ) ) ;
    buf_clk cell_5228 ( .C ( clk ), .D ( signal_10819 ), .Q ( signal_10820 ) ) ;
    buf_clk cell_5234 ( .C ( clk ), .D ( signal_10825 ), .Q ( signal_10826 ) ) ;
    buf_clk cell_5240 ( .C ( clk ), .D ( signal_10831 ), .Q ( signal_10832 ) ) ;
    buf_clk cell_5248 ( .C ( clk ), .D ( signal_10839 ), .Q ( signal_10840 ) ) ;
    buf_clk cell_5256 ( .C ( clk ), .D ( signal_10847 ), .Q ( signal_10848 ) ) ;
    buf_clk cell_5264 ( .C ( clk ), .D ( signal_10855 ), .Q ( signal_10856 ) ) ;
    buf_clk cell_5272 ( .C ( clk ), .D ( signal_10863 ), .Q ( signal_10864 ) ) ;
    buf_clk cell_5280 ( .C ( clk ), .D ( signal_10871 ), .Q ( signal_10872 ) ) ;
    buf_clk cell_5288 ( .C ( clk ), .D ( signal_10879 ), .Q ( signal_10880 ) ) ;
    buf_clk cell_5296 ( .C ( clk ), .D ( signal_10887 ), .Q ( signal_10888 ) ) ;
    buf_clk cell_5304 ( .C ( clk ), .D ( signal_10895 ), .Q ( signal_10896 ) ) ;
    buf_clk cell_5312 ( .C ( clk ), .D ( signal_10903 ), .Q ( signal_10904 ) ) ;
    buf_clk cell_5322 ( .C ( clk ), .D ( signal_10913 ), .Q ( signal_10914 ) ) ;
    buf_clk cell_5332 ( .C ( clk ), .D ( signal_10923 ), .Q ( signal_10924 ) ) ;
    buf_clk cell_5342 ( .C ( clk ), .D ( signal_10933 ), .Q ( signal_10934 ) ) ;
    buf_clk cell_5350 ( .C ( clk ), .D ( signal_10941 ), .Q ( signal_10942 ) ) ;
    buf_clk cell_5358 ( .C ( clk ), .D ( signal_10949 ), .Q ( signal_10950 ) ) ;
    buf_clk cell_5366 ( .C ( clk ), .D ( signal_10957 ), .Q ( signal_10958 ) ) ;
    buf_clk cell_5374 ( .C ( clk ), .D ( signal_10965 ), .Q ( signal_10966 ) ) ;
    buf_clk cell_5382 ( .C ( clk ), .D ( signal_10973 ), .Q ( signal_10974 ) ) ;
    buf_clk cell_5390 ( .C ( clk ), .D ( signal_10981 ), .Q ( signal_10982 ) ) ;
    buf_clk cell_5392 ( .C ( clk ), .D ( signal_10983 ), .Q ( signal_10984 ) ) ;
    buf_clk cell_5394 ( .C ( clk ), .D ( signal_10985 ), .Q ( signal_10986 ) ) ;
    buf_clk cell_5396 ( .C ( clk ), .D ( signal_10987 ), .Q ( signal_10988 ) ) ;
    buf_clk cell_5404 ( .C ( clk ), .D ( signal_10995 ), .Q ( signal_10996 ) ) ;
    buf_clk cell_5412 ( .C ( clk ), .D ( signal_11003 ), .Q ( signal_11004 ) ) ;
    buf_clk cell_5420 ( .C ( clk ), .D ( signal_11011 ), .Q ( signal_11012 ) ) ;
    buf_clk cell_5428 ( .C ( clk ), .D ( signal_11019 ), .Q ( signal_11020 ) ) ;
    buf_clk cell_5436 ( .C ( clk ), .D ( signal_11027 ), .Q ( signal_11028 ) ) ;
    buf_clk cell_5444 ( .C ( clk ), .D ( signal_11035 ), .Q ( signal_11036 ) ) ;
    buf_clk cell_5452 ( .C ( clk ), .D ( signal_11043 ), .Q ( signal_11044 ) ) ;
    buf_clk cell_5460 ( .C ( clk ), .D ( signal_11051 ), .Q ( signal_11052 ) ) ;
    buf_clk cell_5468 ( .C ( clk ), .D ( signal_11059 ), .Q ( signal_11060 ) ) ;
    buf_clk cell_5472 ( .C ( clk ), .D ( signal_11063 ), .Q ( signal_11064 ) ) ;
    buf_clk cell_5478 ( .C ( clk ), .D ( signal_11069 ), .Q ( signal_11070 ) ) ;
    buf_clk cell_5484 ( .C ( clk ), .D ( signal_11075 ), .Q ( signal_11076 ) ) ;
    buf_clk cell_5492 ( .C ( clk ), .D ( signal_11083 ), .Q ( signal_11084 ) ) ;
    buf_clk cell_5500 ( .C ( clk ), .D ( signal_11091 ), .Q ( signal_11092 ) ) ;
    buf_clk cell_5508 ( .C ( clk ), .D ( signal_11099 ), .Q ( signal_11100 ) ) ;
    buf_clk cell_5514 ( .C ( clk ), .D ( signal_11105 ), .Q ( signal_11106 ) ) ;
    buf_clk cell_5520 ( .C ( clk ), .D ( signal_11111 ), .Q ( signal_11112 ) ) ;
    buf_clk cell_5526 ( .C ( clk ), .D ( signal_11117 ), .Q ( signal_11118 ) ) ;
    buf_clk cell_5532 ( .C ( clk ), .D ( signal_11123 ), .Q ( signal_11124 ) ) ;
    buf_clk cell_5538 ( .C ( clk ), .D ( signal_11129 ), .Q ( signal_11130 ) ) ;
    buf_clk cell_5544 ( .C ( clk ), .D ( signal_11135 ), .Q ( signal_11136 ) ) ;
    buf_clk cell_5552 ( .C ( clk ), .D ( signal_11143 ), .Q ( signal_11144 ) ) ;
    buf_clk cell_5560 ( .C ( clk ), .D ( signal_11151 ), .Q ( signal_11152 ) ) ;
    buf_clk cell_5568 ( .C ( clk ), .D ( signal_11159 ), .Q ( signal_11160 ) ) ;
    buf_clk cell_5578 ( .C ( clk ), .D ( signal_11169 ), .Q ( signal_11170 ) ) ;
    buf_clk cell_5588 ( .C ( clk ), .D ( signal_11179 ), .Q ( signal_11180 ) ) ;
    buf_clk cell_5598 ( .C ( clk ), .D ( signal_11189 ), .Q ( signal_11190 ) ) ;
    buf_clk cell_5610 ( .C ( clk ), .D ( signal_11201 ), .Q ( signal_11202 ) ) ;
    buf_clk cell_5616 ( .C ( clk ), .D ( signal_11207 ), .Q ( signal_11208 ) ) ;
    buf_clk cell_5622 ( .C ( clk ), .D ( signal_11213 ), .Q ( signal_11214 ) ) ;
    buf_clk cell_5630 ( .C ( clk ), .D ( signal_11221 ), .Q ( signal_11222 ) ) ;
    buf_clk cell_5638 ( .C ( clk ), .D ( signal_11229 ), .Q ( signal_11230 ) ) ;
    buf_clk cell_5646 ( .C ( clk ), .D ( signal_11237 ), .Q ( signal_11238 ) ) ;
    buf_clk cell_5656 ( .C ( clk ), .D ( signal_11247 ), .Q ( signal_11248 ) ) ;
    buf_clk cell_5666 ( .C ( clk ), .D ( signal_11257 ), .Q ( signal_11258 ) ) ;
    buf_clk cell_5676 ( .C ( clk ), .D ( signal_11267 ), .Q ( signal_11268 ) ) ;
    buf_clk cell_5684 ( .C ( clk ), .D ( signal_11275 ), .Q ( signal_11276 ) ) ;
    buf_clk cell_5692 ( .C ( clk ), .D ( signal_11283 ), .Q ( signal_11284 ) ) ;
    buf_clk cell_5700 ( .C ( clk ), .D ( signal_11291 ), .Q ( signal_11292 ) ) ;
    buf_clk cell_5706 ( .C ( clk ), .D ( signal_11297 ), .Q ( signal_11298 ) ) ;
    buf_clk cell_5712 ( .C ( clk ), .D ( signal_11303 ), .Q ( signal_11304 ) ) ;
    buf_clk cell_5718 ( .C ( clk ), .D ( signal_11309 ), .Q ( signal_11310 ) ) ;
    buf_clk cell_5724 ( .C ( clk ), .D ( signal_11315 ), .Q ( signal_11316 ) ) ;
    buf_clk cell_5730 ( .C ( clk ), .D ( signal_11321 ), .Q ( signal_11322 ) ) ;
    buf_clk cell_5736 ( .C ( clk ), .D ( signal_11327 ), .Q ( signal_11328 ) ) ;
    buf_clk cell_5746 ( .C ( clk ), .D ( signal_11337 ), .Q ( signal_11338 ) ) ;
    buf_clk cell_5750 ( .C ( clk ), .D ( signal_11341 ), .Q ( signal_11342 ) ) ;
    buf_clk cell_5754 ( .C ( clk ), .D ( signal_11345 ), .Q ( signal_11346 ) ) ;
    buf_clk cell_5758 ( .C ( clk ), .D ( signal_11349 ), .Q ( signal_11350 ) ) ;
    buf_clk cell_5762 ( .C ( clk ), .D ( signal_11353 ), .Q ( signal_11354 ) ) ;
    buf_clk cell_5766 ( .C ( clk ), .D ( signal_11357 ), .Q ( signal_11358 ) ) ;
    buf_clk cell_5772 ( .C ( clk ), .D ( signal_11363 ), .Q ( signal_11364 ) ) ;
    buf_clk cell_5778 ( .C ( clk ), .D ( signal_11369 ), .Q ( signal_11370 ) ) ;
    buf_clk cell_5784 ( .C ( clk ), .D ( signal_11375 ), .Q ( signal_11376 ) ) ;
    buf_clk cell_5796 ( .C ( clk ), .D ( signal_11387 ), .Q ( signal_11388 ) ) ;
    buf_clk cell_5802 ( .C ( clk ), .D ( signal_11393 ), .Q ( signal_11394 ) ) ;
    buf_clk cell_5808 ( .C ( clk ), .D ( signal_11399 ), .Q ( signal_11400 ) ) ;
    buf_clk cell_5812 ( .C ( clk ), .D ( signal_11403 ), .Q ( signal_11404 ) ) ;
    buf_clk cell_5816 ( .C ( clk ), .D ( signal_11407 ), .Q ( signal_11408 ) ) ;
    buf_clk cell_5820 ( .C ( clk ), .D ( signal_11411 ), .Q ( signal_11412 ) ) ;
    buf_clk cell_5826 ( .C ( clk ), .D ( signal_11417 ), .Q ( signal_11418 ) ) ;
    buf_clk cell_5832 ( .C ( clk ), .D ( signal_11423 ), .Q ( signal_11424 ) ) ;
    buf_clk cell_5838 ( .C ( clk ), .D ( signal_11429 ), .Q ( signal_11430 ) ) ;
    buf_clk cell_5848 ( .C ( clk ), .D ( signal_11439 ), .Q ( signal_11440 ) ) ;
    buf_clk cell_5852 ( .C ( clk ), .D ( signal_11443 ), .Q ( signal_11444 ) ) ;
    buf_clk cell_5856 ( .C ( clk ), .D ( signal_11447 ), .Q ( signal_11448 ) ) ;
    buf_clk cell_5860 ( .C ( clk ), .D ( signal_11451 ), .Q ( signal_11452 ) ) ;
    buf_clk cell_5866 ( .C ( clk ), .D ( signal_11457 ), .Q ( signal_11458 ) ) ;
    buf_clk cell_5872 ( .C ( clk ), .D ( signal_11463 ), .Q ( signal_11464 ) ) ;
    buf_clk cell_5880 ( .C ( clk ), .D ( signal_11471 ), .Q ( signal_11472 ) ) ;
    buf_clk cell_5888 ( .C ( clk ), .D ( signal_11479 ), .Q ( signal_11480 ) ) ;
    buf_clk cell_5896 ( .C ( clk ), .D ( signal_11487 ), .Q ( signal_11488 ) ) ;
    buf_clk cell_5902 ( .C ( clk ), .D ( signal_11493 ), .Q ( signal_11494 ) ) ;
    buf_clk cell_5908 ( .C ( clk ), .D ( signal_11499 ), .Q ( signal_11500 ) ) ;
    buf_clk cell_5914 ( .C ( clk ), .D ( signal_11505 ), .Q ( signal_11506 ) ) ;
    buf_clk cell_5924 ( .C ( clk ), .D ( signal_11515 ), .Q ( signal_11516 ) ) ;
    buf_clk cell_5934 ( .C ( clk ), .D ( signal_11525 ), .Q ( signal_11526 ) ) ;
    buf_clk cell_5944 ( .C ( clk ), .D ( signal_11535 ), .Q ( signal_11536 ) ) ;
    buf_clk cell_5950 ( .C ( clk ), .D ( signal_11541 ), .Q ( signal_11542 ) ) ;
    buf_clk cell_5956 ( .C ( clk ), .D ( signal_11547 ), .Q ( signal_11548 ) ) ;
    buf_clk cell_5962 ( .C ( clk ), .D ( signal_11553 ), .Q ( signal_11554 ) ) ;
    buf_clk cell_5982 ( .C ( clk ), .D ( signal_11573 ), .Q ( signal_11574 ) ) ;
    buf_clk cell_5990 ( .C ( clk ), .D ( signal_11581 ), .Q ( signal_11582 ) ) ;
    buf_clk cell_5998 ( .C ( clk ), .D ( signal_11589 ), .Q ( signal_11590 ) ) ;
    buf_clk cell_6004 ( .C ( clk ), .D ( signal_11595 ), .Q ( signal_11596 ) ) ;
    buf_clk cell_6010 ( .C ( clk ), .D ( signal_11601 ), .Q ( signal_11602 ) ) ;
    buf_clk cell_6016 ( .C ( clk ), .D ( signal_11607 ), .Q ( signal_11608 ) ) ;
    buf_clk cell_6024 ( .C ( clk ), .D ( signal_11615 ), .Q ( signal_11616 ) ) ;
    buf_clk cell_6032 ( .C ( clk ), .D ( signal_11623 ), .Q ( signal_11624 ) ) ;
    buf_clk cell_6040 ( .C ( clk ), .D ( signal_11631 ), .Q ( signal_11632 ) ) ;
    buf_clk cell_6046 ( .C ( clk ), .D ( signal_11637 ), .Q ( signal_11638 ) ) ;
    buf_clk cell_6052 ( .C ( clk ), .D ( signal_11643 ), .Q ( signal_11644 ) ) ;
    buf_clk cell_6058 ( .C ( clk ), .D ( signal_11649 ), .Q ( signal_11650 ) ) ;
    buf_clk cell_6066 ( .C ( clk ), .D ( signal_11657 ), .Q ( signal_11658 ) ) ;
    buf_clk cell_6074 ( .C ( clk ), .D ( signal_11665 ), .Q ( signal_11666 ) ) ;
    buf_clk cell_6082 ( .C ( clk ), .D ( signal_11673 ), .Q ( signal_11674 ) ) ;
    buf_clk cell_6100 ( .C ( clk ), .D ( signal_11691 ), .Q ( signal_11692 ) ) ;
    buf_clk cell_6106 ( .C ( clk ), .D ( signal_11697 ), .Q ( signal_11698 ) ) ;
    buf_clk cell_6112 ( .C ( clk ), .D ( signal_11703 ), .Q ( signal_11704 ) ) ;
    buf_clk cell_6118 ( .C ( clk ), .D ( signal_11709 ), .Q ( signal_11710 ) ) ;
    buf_clk cell_6124 ( .C ( clk ), .D ( signal_11715 ), .Q ( signal_11716 ) ) ;
    buf_clk cell_6130 ( .C ( clk ), .D ( signal_11721 ), .Q ( signal_11722 ) ) ;
    buf_clk cell_6160 ( .C ( clk ), .D ( signal_11751 ), .Q ( signal_11752 ) ) ;
    buf_clk cell_6168 ( .C ( clk ), .D ( signal_11759 ), .Q ( signal_11760 ) ) ;
    buf_clk cell_6176 ( .C ( clk ), .D ( signal_11767 ), .Q ( signal_11768 ) ) ;
    buf_clk cell_6188 ( .C ( clk ), .D ( signal_11779 ), .Q ( signal_11780 ) ) ;
    buf_clk cell_6200 ( .C ( clk ), .D ( signal_11791 ), .Q ( signal_11792 ) ) ;
    buf_clk cell_6212 ( .C ( clk ), .D ( signal_11803 ), .Q ( signal_11804 ) ) ;
    buf_clk cell_6262 ( .C ( clk ), .D ( signal_11853 ), .Q ( signal_11854 ) ) ;
    buf_clk cell_6276 ( .C ( clk ), .D ( signal_11867 ), .Q ( signal_11868 ) ) ;
    buf_clk cell_6290 ( .C ( clk ), .D ( signal_11881 ), .Q ( signal_11882 ) ) ;
    buf_clk cell_6298 ( .C ( clk ), .D ( signal_11889 ), .Q ( signal_11890 ) ) ;
    buf_clk cell_6306 ( .C ( clk ), .D ( signal_11897 ), .Q ( signal_11898 ) ) ;
    buf_clk cell_6314 ( .C ( clk ), .D ( signal_11905 ), .Q ( signal_11906 ) ) ;
    buf_clk cell_6328 ( .C ( clk ), .D ( signal_11919 ), .Q ( signal_11920 ) ) ;
    buf_clk cell_6342 ( .C ( clk ), .D ( signal_11933 ), .Q ( signal_11934 ) ) ;
    buf_clk cell_6356 ( .C ( clk ), .D ( signal_11947 ), .Q ( signal_11948 ) ) ;
    buf_clk cell_6364 ( .C ( clk ), .D ( signal_11955 ), .Q ( signal_11956 ) ) ;
    buf_clk cell_6372 ( .C ( clk ), .D ( signal_11963 ), .Q ( signal_11964 ) ) ;
    buf_clk cell_6380 ( .C ( clk ), .D ( signal_11971 ), .Q ( signal_11972 ) ) ;
    buf_clk cell_6400 ( .C ( clk ), .D ( signal_11991 ), .Q ( signal_11992 ) ) ;
    buf_clk cell_6410 ( .C ( clk ), .D ( signal_12001 ), .Q ( signal_12002 ) ) ;
    buf_clk cell_6420 ( .C ( clk ), .D ( signal_12011 ), .Q ( signal_12012 ) ) ;
    buf_clk cell_6448 ( .C ( clk ), .D ( signal_12039 ), .Q ( signal_12040 ) ) ;
    buf_clk cell_6464 ( .C ( clk ), .D ( signal_12055 ), .Q ( signal_12056 ) ) ;
    buf_clk cell_6480 ( .C ( clk ), .D ( signal_12071 ), .Q ( signal_12072 ) ) ;
    buf_clk cell_6508 ( .C ( clk ), .D ( signal_12099 ), .Q ( signal_12100 ) ) ;
    buf_clk cell_6524 ( .C ( clk ), .D ( signal_12115 ), .Q ( signal_12116 ) ) ;
    buf_clk cell_6540 ( .C ( clk ), .D ( signal_12131 ), .Q ( signal_12132 ) ) ;
    buf_clk cell_6550 ( .C ( clk ), .D ( signal_12141 ), .Q ( signal_12142 ) ) ;
    buf_clk cell_6560 ( .C ( clk ), .D ( signal_12151 ), .Q ( signal_12152 ) ) ;
    buf_clk cell_6570 ( .C ( clk ), .D ( signal_12161 ), .Q ( signal_12162 ) ) ;
    buf_clk cell_6692 ( .C ( clk ), .D ( signal_12283 ), .Q ( signal_12284 ) ) ;
    buf_clk cell_6708 ( .C ( clk ), .D ( signal_12299 ), .Q ( signal_12300 ) ) ;
    buf_clk cell_6724 ( .C ( clk ), .D ( signal_12315 ), .Q ( signal_12316 ) ) ;
    buf_clk cell_6742 ( .C ( clk ), .D ( signal_12333 ), .Q ( signal_12334 ) ) ;
    buf_clk cell_6760 ( .C ( clk ), .D ( signal_12351 ), .Q ( signal_12352 ) ) ;
    buf_clk cell_6778 ( .C ( clk ), .D ( signal_12369 ), .Q ( signal_12370 ) ) ;
    buf_clk cell_6892 ( .C ( clk ), .D ( signal_12483 ), .Q ( signal_12484 ) ) ;
    buf_clk cell_6912 ( .C ( clk ), .D ( signal_12503 ), .Q ( signal_12504 ) ) ;
    buf_clk cell_6932 ( .C ( clk ), .D ( signal_12523 ), .Q ( signal_12524 ) ) ;

    /* cells in depth 15 */
    buf_clk cell_5473 ( .C ( clk ), .D ( signal_11064 ), .Q ( signal_11065 ) ) ;
    buf_clk cell_5479 ( .C ( clk ), .D ( signal_11070 ), .Q ( signal_11071 ) ) ;
    buf_clk cell_5485 ( .C ( clk ), .D ( signal_11076 ), .Q ( signal_11077 ) ) ;
    buf_clk cell_5493 ( .C ( clk ), .D ( signal_11084 ), .Q ( signal_11085 ) ) ;
    buf_clk cell_5501 ( .C ( clk ), .D ( signal_11092 ), .Q ( signal_11093 ) ) ;
    buf_clk cell_5509 ( .C ( clk ), .D ( signal_11100 ), .Q ( signal_11101 ) ) ;
    buf_clk cell_5515 ( .C ( clk ), .D ( signal_11106 ), .Q ( signal_11107 ) ) ;
    buf_clk cell_5521 ( .C ( clk ), .D ( signal_11112 ), .Q ( signal_11113 ) ) ;
    buf_clk cell_5527 ( .C ( clk ), .D ( signal_11118 ), .Q ( signal_11119 ) ) ;
    buf_clk cell_5533 ( .C ( clk ), .D ( signal_11124 ), .Q ( signal_11125 ) ) ;
    buf_clk cell_5539 ( .C ( clk ), .D ( signal_11130 ), .Q ( signal_11131 ) ) ;
    buf_clk cell_5545 ( .C ( clk ), .D ( signal_11136 ), .Q ( signal_11137 ) ) ;
    buf_clk cell_5553 ( .C ( clk ), .D ( signal_11144 ), .Q ( signal_11145 ) ) ;
    buf_clk cell_5561 ( .C ( clk ), .D ( signal_11152 ), .Q ( signal_11153 ) ) ;
    buf_clk cell_5569 ( .C ( clk ), .D ( signal_11160 ), .Q ( signal_11161 ) ) ;
    buf_clk cell_5579 ( .C ( clk ), .D ( signal_11170 ), .Q ( signal_11171 ) ) ;
    buf_clk cell_5589 ( .C ( clk ), .D ( signal_11180 ), .Q ( signal_11181 ) ) ;
    buf_clk cell_5599 ( .C ( clk ), .D ( signal_11190 ), .Q ( signal_11191 ) ) ;
    buf_clk cell_5601 ( .C ( clk ), .D ( signal_2258 ), .Q ( signal_11193 ) ) ;
    buf_clk cell_5603 ( .C ( clk ), .D ( signal_5040 ), .Q ( signal_11195 ) ) ;
    buf_clk cell_5605 ( .C ( clk ), .D ( signal_5041 ), .Q ( signal_11197 ) ) ;
    buf_clk cell_5611 ( .C ( clk ), .D ( signal_11202 ), .Q ( signal_11203 ) ) ;
    buf_clk cell_5617 ( .C ( clk ), .D ( signal_11208 ), .Q ( signal_11209 ) ) ;
    buf_clk cell_5623 ( .C ( clk ), .D ( signal_11214 ), .Q ( signal_11215 ) ) ;
    buf_clk cell_5631 ( .C ( clk ), .D ( signal_11222 ), .Q ( signal_11223 ) ) ;
    buf_clk cell_5639 ( .C ( clk ), .D ( signal_11230 ), .Q ( signal_11231 ) ) ;
    buf_clk cell_5647 ( .C ( clk ), .D ( signal_11238 ), .Q ( signal_11239 ) ) ;
    buf_clk cell_5657 ( .C ( clk ), .D ( signal_11248 ), .Q ( signal_11249 ) ) ;
    buf_clk cell_5667 ( .C ( clk ), .D ( signal_11258 ), .Q ( signal_11259 ) ) ;
    buf_clk cell_5677 ( .C ( clk ), .D ( signal_11268 ), .Q ( signal_11269 ) ) ;
    buf_clk cell_5685 ( .C ( clk ), .D ( signal_11276 ), .Q ( signal_11277 ) ) ;
    buf_clk cell_5693 ( .C ( clk ), .D ( signal_11284 ), .Q ( signal_11285 ) ) ;
    buf_clk cell_5701 ( .C ( clk ), .D ( signal_11292 ), .Q ( signal_11293 ) ) ;
    buf_clk cell_5707 ( .C ( clk ), .D ( signal_11298 ), .Q ( signal_11299 ) ) ;
    buf_clk cell_5713 ( .C ( clk ), .D ( signal_11304 ), .Q ( signal_11305 ) ) ;
    buf_clk cell_5719 ( .C ( clk ), .D ( signal_11310 ), .Q ( signal_11311 ) ) ;
    buf_clk cell_5725 ( .C ( clk ), .D ( signal_11316 ), .Q ( signal_11317 ) ) ;
    buf_clk cell_5731 ( .C ( clk ), .D ( signal_11322 ), .Q ( signal_11323 ) ) ;
    buf_clk cell_5737 ( .C ( clk ), .D ( signal_11328 ), .Q ( signal_11329 ) ) ;
    buf_clk cell_5739 ( .C ( clk ), .D ( signal_10714 ), .Q ( signal_11331 ) ) ;
    buf_clk cell_5741 ( .C ( clk ), .D ( signal_10716 ), .Q ( signal_11333 ) ) ;
    buf_clk cell_5743 ( .C ( clk ), .D ( signal_10718 ), .Q ( signal_11335 ) ) ;
    buf_clk cell_5747 ( .C ( clk ), .D ( signal_11338 ), .Q ( signal_11339 ) ) ;
    buf_clk cell_5751 ( .C ( clk ), .D ( signal_11342 ), .Q ( signal_11343 ) ) ;
    buf_clk cell_5755 ( .C ( clk ), .D ( signal_11346 ), .Q ( signal_11347 ) ) ;
    buf_clk cell_5759 ( .C ( clk ), .D ( signal_11350 ), .Q ( signal_11351 ) ) ;
    buf_clk cell_5763 ( .C ( clk ), .D ( signal_11354 ), .Q ( signal_11355 ) ) ;
    buf_clk cell_5767 ( .C ( clk ), .D ( signal_11358 ), .Q ( signal_11359 ) ) ;
    buf_clk cell_5773 ( .C ( clk ), .D ( signal_11364 ), .Q ( signal_11365 ) ) ;
    buf_clk cell_5779 ( .C ( clk ), .D ( signal_11370 ), .Q ( signal_11371 ) ) ;
    buf_clk cell_5785 ( .C ( clk ), .D ( signal_11376 ), .Q ( signal_11377 ) ) ;
    buf_clk cell_5787 ( .C ( clk ), .D ( signal_2287 ), .Q ( signal_11379 ) ) ;
    buf_clk cell_5789 ( .C ( clk ), .D ( signal_5098 ), .Q ( signal_11381 ) ) ;
    buf_clk cell_5791 ( .C ( clk ), .D ( signal_5099 ), .Q ( signal_11383 ) ) ;
    buf_clk cell_5797 ( .C ( clk ), .D ( signal_11388 ), .Q ( signal_11389 ) ) ;
    buf_clk cell_5803 ( .C ( clk ), .D ( signal_11394 ), .Q ( signal_11395 ) ) ;
    buf_clk cell_5809 ( .C ( clk ), .D ( signal_11400 ), .Q ( signal_11401 ) ) ;
    buf_clk cell_5813 ( .C ( clk ), .D ( signal_11404 ), .Q ( signal_11405 ) ) ;
    buf_clk cell_5817 ( .C ( clk ), .D ( signal_11408 ), .Q ( signal_11409 ) ) ;
    buf_clk cell_5821 ( .C ( clk ), .D ( signal_11412 ), .Q ( signal_11413 ) ) ;
    buf_clk cell_5827 ( .C ( clk ), .D ( signal_11418 ), .Q ( signal_11419 ) ) ;
    buf_clk cell_5833 ( .C ( clk ), .D ( signal_11424 ), .Q ( signal_11425 ) ) ;
    buf_clk cell_5839 ( .C ( clk ), .D ( signal_11430 ), .Q ( signal_11431 ) ) ;
    buf_clk cell_5841 ( .C ( clk ), .D ( signal_2312 ), .Q ( signal_11433 ) ) ;
    buf_clk cell_5843 ( .C ( clk ), .D ( signal_5148 ), .Q ( signal_11435 ) ) ;
    buf_clk cell_5845 ( .C ( clk ), .D ( signal_5149 ), .Q ( signal_11437 ) ) ;
    buf_clk cell_5849 ( .C ( clk ), .D ( signal_11440 ), .Q ( signal_11441 ) ) ;
    buf_clk cell_5853 ( .C ( clk ), .D ( signal_11444 ), .Q ( signal_11445 ) ) ;
    buf_clk cell_5857 ( .C ( clk ), .D ( signal_11448 ), .Q ( signal_11449 ) ) ;
    buf_clk cell_5861 ( .C ( clk ), .D ( signal_11452 ), .Q ( signal_11453 ) ) ;
    buf_clk cell_5867 ( .C ( clk ), .D ( signal_11458 ), .Q ( signal_11459 ) ) ;
    buf_clk cell_5873 ( .C ( clk ), .D ( signal_11464 ), .Q ( signal_11465 ) ) ;
    buf_clk cell_5881 ( .C ( clk ), .D ( signal_11472 ), .Q ( signal_11473 ) ) ;
    buf_clk cell_5889 ( .C ( clk ), .D ( signal_11480 ), .Q ( signal_11481 ) ) ;
    buf_clk cell_5897 ( .C ( clk ), .D ( signal_11488 ), .Q ( signal_11489 ) ) ;
    buf_clk cell_5903 ( .C ( clk ), .D ( signal_11494 ), .Q ( signal_11495 ) ) ;
    buf_clk cell_5909 ( .C ( clk ), .D ( signal_11500 ), .Q ( signal_11501 ) ) ;
    buf_clk cell_5915 ( .C ( clk ), .D ( signal_11506 ), .Q ( signal_11507 ) ) ;
    buf_clk cell_5925 ( .C ( clk ), .D ( signal_11516 ), .Q ( signal_11517 ) ) ;
    buf_clk cell_5935 ( .C ( clk ), .D ( signal_11526 ), .Q ( signal_11527 ) ) ;
    buf_clk cell_5945 ( .C ( clk ), .D ( signal_11536 ), .Q ( signal_11537 ) ) ;
    buf_clk cell_5951 ( .C ( clk ), .D ( signal_11542 ), .Q ( signal_11543 ) ) ;
    buf_clk cell_5957 ( .C ( clk ), .D ( signal_11548 ), .Q ( signal_11549 ) ) ;
    buf_clk cell_5963 ( .C ( clk ), .D ( signal_11554 ), .Q ( signal_11555 ) ) ;
    buf_clk cell_5967 ( .C ( clk ), .D ( signal_2288 ), .Q ( signal_11559 ) ) ;
    buf_clk cell_5971 ( .C ( clk ), .D ( signal_5100 ), .Q ( signal_11563 ) ) ;
    buf_clk cell_5975 ( .C ( clk ), .D ( signal_5101 ), .Q ( signal_11567 ) ) ;
    buf_clk cell_5983 ( .C ( clk ), .D ( signal_11574 ), .Q ( signal_11575 ) ) ;
    buf_clk cell_5991 ( .C ( clk ), .D ( signal_11582 ), .Q ( signal_11583 ) ) ;
    buf_clk cell_5999 ( .C ( clk ), .D ( signal_11590 ), .Q ( signal_11591 ) ) ;
    buf_clk cell_6005 ( .C ( clk ), .D ( signal_11596 ), .Q ( signal_11597 ) ) ;
    buf_clk cell_6011 ( .C ( clk ), .D ( signal_11602 ), .Q ( signal_11603 ) ) ;
    buf_clk cell_6017 ( .C ( clk ), .D ( signal_11608 ), .Q ( signal_11609 ) ) ;
    buf_clk cell_6025 ( .C ( clk ), .D ( signal_11616 ), .Q ( signal_11617 ) ) ;
    buf_clk cell_6033 ( .C ( clk ), .D ( signal_11624 ), .Q ( signal_11625 ) ) ;
    buf_clk cell_6041 ( .C ( clk ), .D ( signal_11632 ), .Q ( signal_11633 ) ) ;
    buf_clk cell_6047 ( .C ( clk ), .D ( signal_11638 ), .Q ( signal_11639 ) ) ;
    buf_clk cell_6053 ( .C ( clk ), .D ( signal_11644 ), .Q ( signal_11645 ) ) ;
    buf_clk cell_6059 ( .C ( clk ), .D ( signal_11650 ), .Q ( signal_11651 ) ) ;
    buf_clk cell_6067 ( .C ( clk ), .D ( signal_11658 ), .Q ( signal_11659 ) ) ;
    buf_clk cell_6075 ( .C ( clk ), .D ( signal_11666 ), .Q ( signal_11667 ) ) ;
    buf_clk cell_6083 ( .C ( clk ), .D ( signal_11674 ), .Q ( signal_11675 ) ) ;
    buf_clk cell_6087 ( .C ( clk ), .D ( signal_2213 ), .Q ( signal_11679 ) ) ;
    buf_clk cell_6091 ( .C ( clk ), .D ( signal_4950 ), .Q ( signal_11683 ) ) ;
    buf_clk cell_6095 ( .C ( clk ), .D ( signal_4951 ), .Q ( signal_11687 ) ) ;
    buf_clk cell_6101 ( .C ( clk ), .D ( signal_11692 ), .Q ( signal_11693 ) ) ;
    buf_clk cell_6107 ( .C ( clk ), .D ( signal_11698 ), .Q ( signal_11699 ) ) ;
    buf_clk cell_6113 ( .C ( clk ), .D ( signal_11704 ), .Q ( signal_11705 ) ) ;
    buf_clk cell_6119 ( .C ( clk ), .D ( signal_11710 ), .Q ( signal_11711 ) ) ;
    buf_clk cell_6125 ( .C ( clk ), .D ( signal_11716 ), .Q ( signal_11717 ) ) ;
    buf_clk cell_6131 ( .C ( clk ), .D ( signal_11722 ), .Q ( signal_11723 ) ) ;
    buf_clk cell_6135 ( .C ( clk ), .D ( signal_2189 ), .Q ( signal_11727 ) ) ;
    buf_clk cell_6139 ( .C ( clk ), .D ( signal_4902 ), .Q ( signal_11731 ) ) ;
    buf_clk cell_6143 ( .C ( clk ), .D ( signal_4903 ), .Q ( signal_11735 ) ) ;
    buf_clk cell_6147 ( .C ( clk ), .D ( signal_2138 ), .Q ( signal_11739 ) ) ;
    buf_clk cell_6151 ( .C ( clk ), .D ( signal_4800 ), .Q ( signal_11743 ) ) ;
    buf_clk cell_6155 ( .C ( clk ), .D ( signal_4801 ), .Q ( signal_11747 ) ) ;
    buf_clk cell_6161 ( .C ( clk ), .D ( signal_11752 ), .Q ( signal_11753 ) ) ;
    buf_clk cell_6169 ( .C ( clk ), .D ( signal_11760 ), .Q ( signal_11761 ) ) ;
    buf_clk cell_6177 ( .C ( clk ), .D ( signal_11768 ), .Q ( signal_11769 ) ) ;
    buf_clk cell_6189 ( .C ( clk ), .D ( signal_11780 ), .Q ( signal_11781 ) ) ;
    buf_clk cell_6201 ( .C ( clk ), .D ( signal_11792 ), .Q ( signal_11793 ) ) ;
    buf_clk cell_6213 ( .C ( clk ), .D ( signal_11804 ), .Q ( signal_11805 ) ) ;
    buf_clk cell_6219 ( .C ( clk ), .D ( signal_2238 ), .Q ( signal_11811 ) ) ;
    buf_clk cell_6225 ( .C ( clk ), .D ( signal_5000 ), .Q ( signal_11817 ) ) ;
    buf_clk cell_6231 ( .C ( clk ), .D ( signal_5001 ), .Q ( signal_11823 ) ) ;
    buf_clk cell_6237 ( .C ( clk ), .D ( signal_2210 ), .Q ( signal_11829 ) ) ;
    buf_clk cell_6243 ( .C ( clk ), .D ( signal_4944 ), .Q ( signal_11835 ) ) ;
    buf_clk cell_6249 ( .C ( clk ), .D ( signal_4945 ), .Q ( signal_11841 ) ) ;
    buf_clk cell_6263 ( .C ( clk ), .D ( signal_11854 ), .Q ( signal_11855 ) ) ;
    buf_clk cell_6277 ( .C ( clk ), .D ( signal_11868 ), .Q ( signal_11869 ) ) ;
    buf_clk cell_6291 ( .C ( clk ), .D ( signal_11882 ), .Q ( signal_11883 ) ) ;
    buf_clk cell_6299 ( .C ( clk ), .D ( signal_11890 ), .Q ( signal_11891 ) ) ;
    buf_clk cell_6307 ( .C ( clk ), .D ( signal_11898 ), .Q ( signal_11899 ) ) ;
    buf_clk cell_6315 ( .C ( clk ), .D ( signal_11906 ), .Q ( signal_11907 ) ) ;
    buf_clk cell_6329 ( .C ( clk ), .D ( signal_11920 ), .Q ( signal_11921 ) ) ;
    buf_clk cell_6343 ( .C ( clk ), .D ( signal_11934 ), .Q ( signal_11935 ) ) ;
    buf_clk cell_6357 ( .C ( clk ), .D ( signal_11948 ), .Q ( signal_11949 ) ) ;
    buf_clk cell_6365 ( .C ( clk ), .D ( signal_11956 ), .Q ( signal_11957 ) ) ;
    buf_clk cell_6373 ( .C ( clk ), .D ( signal_11964 ), .Q ( signal_11965 ) ) ;
    buf_clk cell_6381 ( .C ( clk ), .D ( signal_11972 ), .Q ( signal_11973 ) ) ;
    buf_clk cell_6401 ( .C ( clk ), .D ( signal_11992 ), .Q ( signal_11993 ) ) ;
    buf_clk cell_6411 ( .C ( clk ), .D ( signal_12002 ), .Q ( signal_12003 ) ) ;
    buf_clk cell_6421 ( .C ( clk ), .D ( signal_12012 ), .Q ( signal_12013 ) ) ;
    buf_clk cell_6449 ( .C ( clk ), .D ( signal_12040 ), .Q ( signal_12041 ) ) ;
    buf_clk cell_6465 ( .C ( clk ), .D ( signal_12056 ), .Q ( signal_12057 ) ) ;
    buf_clk cell_6481 ( .C ( clk ), .D ( signal_12072 ), .Q ( signal_12073 ) ) ;
    buf_clk cell_6509 ( .C ( clk ), .D ( signal_12100 ), .Q ( signal_12101 ) ) ;
    buf_clk cell_6525 ( .C ( clk ), .D ( signal_12116 ), .Q ( signal_12117 ) ) ;
    buf_clk cell_6541 ( .C ( clk ), .D ( signal_12132 ), .Q ( signal_12133 ) ) ;
    buf_clk cell_6551 ( .C ( clk ), .D ( signal_12142 ), .Q ( signal_12143 ) ) ;
    buf_clk cell_6561 ( .C ( clk ), .D ( signal_12152 ), .Q ( signal_12153 ) ) ;
    buf_clk cell_6571 ( .C ( clk ), .D ( signal_12162 ), .Q ( signal_12163 ) ) ;
    buf_clk cell_6609 ( .C ( clk ), .D ( signal_2289 ), .Q ( signal_12201 ) ) ;
    buf_clk cell_6619 ( .C ( clk ), .D ( signal_5102 ), .Q ( signal_12211 ) ) ;
    buf_clk cell_6629 ( .C ( clk ), .D ( signal_5103 ), .Q ( signal_12221 ) ) ;
    buf_clk cell_6657 ( .C ( clk ), .D ( signal_2265 ), .Q ( signal_12249 ) ) ;
    buf_clk cell_6667 ( .C ( clk ), .D ( signal_5054 ), .Q ( signal_12259 ) ) ;
    buf_clk cell_6677 ( .C ( clk ), .D ( signal_5055 ), .Q ( signal_12269 ) ) ;
    buf_clk cell_6693 ( .C ( clk ), .D ( signal_12284 ), .Q ( signal_12285 ) ) ;
    buf_clk cell_6709 ( .C ( clk ), .D ( signal_12300 ), .Q ( signal_12301 ) ) ;
    buf_clk cell_6725 ( .C ( clk ), .D ( signal_12316 ), .Q ( signal_12317 ) ) ;
    buf_clk cell_6743 ( .C ( clk ), .D ( signal_12334 ), .Q ( signal_12335 ) ) ;
    buf_clk cell_6761 ( .C ( clk ), .D ( signal_12352 ), .Q ( signal_12353 ) ) ;
    buf_clk cell_6779 ( .C ( clk ), .D ( signal_12370 ), .Q ( signal_12371 ) ) ;
    buf_clk cell_6893 ( .C ( clk ), .D ( signal_12484 ), .Q ( signal_12485 ) ) ;
    buf_clk cell_6913 ( .C ( clk ), .D ( signal_12504 ), .Q ( signal_12505 ) ) ;
    buf_clk cell_6933 ( .C ( clk ), .D ( signal_12524 ), .Q ( signal_12525 ) ) ;

    /* cells in depth 16 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2180 ( .a ({signal_10622, signal_10612, signal_10602}), .b ({signal_4787, signal_4786, signal_2131}), .clk ( clk ), .r ({Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({signal_4915, signal_4914, signal_2195}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2181 ( .a ({signal_10640, signal_10634, signal_10628}), .b ({signal_4791, signal_4790, signal_2133}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319]}), .c ({signal_4917, signal_4916, signal_2196}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2182 ( .a ({signal_10664, signal_10656, signal_10648}), .b ({signal_4797, signal_4796, signal_2136}), .clk ( clk ), .r ({Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({signal_4919, signal_4918, signal_2197}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2183 ( .a ({signal_10688, signal_10680, signal_10672}), .b ({signal_4799, signal_4798, signal_2137}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325]}), .c ({signal_4921, signal_4920, signal_2198}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2199 ( .a ({signal_4915, signal_4914, signal_2195}), .b ({signal_4953, signal_4952, signal_2214}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2225 ( .a ({signal_10700, signal_10696, signal_10692}), .b ({signal_4895, signal_4894, signal_2185}), .clk ( clk ), .r ({Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({signal_5005, signal_5004, signal_2240}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2226 ( .a ({signal_10712, signal_10708, signal_10704}), .b ({signal_4899, signal_4898, signal_2187}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331]}), .c ({signal_5007, signal_5006, signal_2241}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2227 ( .a ({signal_10718, signal_10716, signal_10714}), .b ({signal_4835, signal_4834, signal_2155}), .clk ( clk ), .r ({Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({signal_5009, signal_5008, signal_2242}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2228 ( .a ({signal_4909, signal_4908, signal_2192}), .b ({signal_10724, signal_10722, signal_10720}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337]}), .c ({signal_5011, signal_5010, signal_2243}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2229 ( .a ({signal_10736, signal_10732, signal_10728}), .b ({signal_4913, signal_4912, signal_2194}), .clk ( clk ), .r ({Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_5013, signal_5012, signal_2244}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2244 ( .a ({signal_5005, signal_5004, signal_2240}), .b ({signal_5043, signal_5042, signal_2259}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2245 ( .a ({signal_5009, signal_5008, signal_2242}), .b ({signal_5045, signal_5044, signal_2260}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2246 ( .a ({signal_5013, signal_5012, signal_2244}), .b ({signal_5047, signal_5046, signal_2261}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2247 ( .a ({signal_10766, signal_10756, signal_10746}), .b ({signal_4955, signal_4954, signal_2215}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343]}), .c ({signal_5049, signal_5048, signal_2262}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2255 ( .a ({signal_10784, signal_10778, signal_10772}), .b ({signal_4973, signal_4972, signal_2224}), .clk ( clk ), .r ({Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({signal_5065, signal_5064, signal_2270}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2256 ( .a ({signal_10790, signal_10788, signal_10786}), .b ({signal_4975, signal_4974, signal_2225}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349]}), .c ({signal_5067, signal_5066, signal_2271}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2257 ( .a ({signal_10814, signal_10806, signal_10798}), .b ({signal_4977, signal_4976, signal_2226}), .clk ( clk ), .r ({Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({signal_5069, signal_5068, signal_2272}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2258 ( .a ({signal_10832, signal_10826, signal_10820}), .b ({signal_4979, signal_4978, signal_2227}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355]}), .c ({signal_5071, signal_5070, signal_2273}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2259 ( .a ({signal_10856, signal_10848, signal_10840}), .b ({signal_4983, signal_4982, signal_2229}), .clk ( clk ), .r ({Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({signal_5073, signal_5072, signal_2274}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2260 ( .a ({signal_10880, signal_10872, signal_10864}), .b ({signal_4985, signal_4984, signal_2230}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361]}), .c ({signal_5075, signal_5074, signal_2275}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2261 ( .a ({signal_10904, signal_10896, signal_10888}), .b ({signal_4987, signal_4986, signal_2231}), .clk ( clk ), .r ({Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({signal_5077, signal_5076, signal_2276}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2262 ( .a ({signal_10700, signal_10696, signal_10692}), .b ({signal_4947, signal_4946, signal_2211}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367]}), .c ({signal_5079, signal_5078, signal_2277}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2263 ( .a ({signal_10934, signal_10924, signal_10914}), .b ({signal_4993, signal_4992, signal_2234}), .clk ( clk ), .r ({Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_5081, signal_5080, signal_2278}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2264 ( .a ({signal_4935, signal_4934, signal_2205}), .b ({signal_4995, signal_4994, signal_2235}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373]}), .c ({signal_5083, signal_5082, signal_2279}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2265 ( .a ({signal_10958, signal_10950, signal_10942}), .b ({signal_4949, signal_4948, signal_2212}), .clk ( clk ), .r ({Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({signal_5085, signal_5084, signal_2280}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2266 ( .a ({signal_10982, signal_10974, signal_10966}), .b ({signal_4999, signal_4998, signal_2237}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379]}), .c ({signal_5087, signal_5086, signal_2281}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2275 ( .a ({signal_5067, signal_5066, signal_2271}), .b ({signal_5105, signal_5104, signal_2290}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2276 ( .a ({signal_5069, signal_5068, signal_2272}), .b ({signal_5107, signal_5106, signal_2291}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2277 ( .a ({signal_5073, signal_5072, signal_2274}), .b ({signal_5109, signal_5108, signal_2292}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2278 ( .a ({signal_5077, signal_5076, signal_2276}), .b ({signal_5111, signal_5110, signal_2293}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2279 ( .a ({signal_5079, signal_5078, signal_2277}), .b ({signal_5113, signal_5112, signal_2294}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2280 ( .a ({signal_5085, signal_5084, signal_2280}), .b ({signal_5115, signal_5114, signal_2295}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2287 ( .a ({signal_5053, signal_5052, signal_2264}), .b ({signal_4969, signal_4968, signal_2222}), .clk ( clk ), .r ({Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({signal_5129, signal_5128, signal_2302}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2288 ( .a ({signal_10988, signal_10986, signal_10984}), .b ({signal_5033, signal_5032, signal_2254}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385]}), .c ({signal_5131, signal_5130, signal_2303}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2290 ( .a ({signal_10988, signal_10986, signal_10984}), .b ({signal_5037, signal_5036, signal_2256}), .clk ( clk ), .r ({Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({signal_5135, signal_5134, signal_2305}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2299 ( .a ({signal_5131, signal_5130, signal_2303}), .b ({signal_5153, signal_5152, signal_2314}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2301 ( .a ({signal_5135, signal_5134, signal_2305}), .b ({signal_5157, signal_5156, signal_2316}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2304 ( .a ({signal_11012, signal_11004, signal_10996}), .b ({signal_5119, signal_5118, signal_2297}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391]}), .c ({signal_5163, signal_5162, signal_2319}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2305 ( .a ({signal_11036, signal_11028, signal_11020}), .b ({signal_5125, signal_5124, signal_2300}), .clk ( clk ), .r ({Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({signal_5165, signal_5164, signal_2320}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2306 ( .a ({signal_11060, signal_11052, signal_11044}), .b ({signal_5127, signal_5126, signal_2301}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397]}), .c ({signal_5167, signal_5166, signal_2321}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2307 ( .a ({signal_5097, signal_5096, signal_2286}), .b ({signal_4991, signal_4990, signal_2233}), .clk ( clk ), .r ({Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_5169, signal_5168, signal_2322}) ) ;
    buf_clk cell_5474 ( .C ( clk ), .D ( signal_11065 ), .Q ( signal_11066 ) ) ;
    buf_clk cell_5480 ( .C ( clk ), .D ( signal_11071 ), .Q ( signal_11072 ) ) ;
    buf_clk cell_5486 ( .C ( clk ), .D ( signal_11077 ), .Q ( signal_11078 ) ) ;
    buf_clk cell_5494 ( .C ( clk ), .D ( signal_11085 ), .Q ( signal_11086 ) ) ;
    buf_clk cell_5502 ( .C ( clk ), .D ( signal_11093 ), .Q ( signal_11094 ) ) ;
    buf_clk cell_5510 ( .C ( clk ), .D ( signal_11101 ), .Q ( signal_11102 ) ) ;
    buf_clk cell_5516 ( .C ( clk ), .D ( signal_11107 ), .Q ( signal_11108 ) ) ;
    buf_clk cell_5522 ( .C ( clk ), .D ( signal_11113 ), .Q ( signal_11114 ) ) ;
    buf_clk cell_5528 ( .C ( clk ), .D ( signal_11119 ), .Q ( signal_11120 ) ) ;
    buf_clk cell_5534 ( .C ( clk ), .D ( signal_11125 ), .Q ( signal_11126 ) ) ;
    buf_clk cell_5540 ( .C ( clk ), .D ( signal_11131 ), .Q ( signal_11132 ) ) ;
    buf_clk cell_5546 ( .C ( clk ), .D ( signal_11137 ), .Q ( signal_11138 ) ) ;
    buf_clk cell_5554 ( .C ( clk ), .D ( signal_11145 ), .Q ( signal_11146 ) ) ;
    buf_clk cell_5562 ( .C ( clk ), .D ( signal_11153 ), .Q ( signal_11154 ) ) ;
    buf_clk cell_5570 ( .C ( clk ), .D ( signal_11161 ), .Q ( signal_11162 ) ) ;
    buf_clk cell_5580 ( .C ( clk ), .D ( signal_11171 ), .Q ( signal_11172 ) ) ;
    buf_clk cell_5590 ( .C ( clk ), .D ( signal_11181 ), .Q ( signal_11182 ) ) ;
    buf_clk cell_5600 ( .C ( clk ), .D ( signal_11191 ), .Q ( signal_11192 ) ) ;
    buf_clk cell_5602 ( .C ( clk ), .D ( signal_11193 ), .Q ( signal_11194 ) ) ;
    buf_clk cell_5604 ( .C ( clk ), .D ( signal_11195 ), .Q ( signal_11196 ) ) ;
    buf_clk cell_5606 ( .C ( clk ), .D ( signal_11197 ), .Q ( signal_11198 ) ) ;
    buf_clk cell_5612 ( .C ( clk ), .D ( signal_11203 ), .Q ( signal_11204 ) ) ;
    buf_clk cell_5618 ( .C ( clk ), .D ( signal_11209 ), .Q ( signal_11210 ) ) ;
    buf_clk cell_5624 ( .C ( clk ), .D ( signal_11215 ), .Q ( signal_11216 ) ) ;
    buf_clk cell_5632 ( .C ( clk ), .D ( signal_11223 ), .Q ( signal_11224 ) ) ;
    buf_clk cell_5640 ( .C ( clk ), .D ( signal_11231 ), .Q ( signal_11232 ) ) ;
    buf_clk cell_5648 ( .C ( clk ), .D ( signal_11239 ), .Q ( signal_11240 ) ) ;
    buf_clk cell_5658 ( .C ( clk ), .D ( signal_11249 ), .Q ( signal_11250 ) ) ;
    buf_clk cell_5668 ( .C ( clk ), .D ( signal_11259 ), .Q ( signal_11260 ) ) ;
    buf_clk cell_5678 ( .C ( clk ), .D ( signal_11269 ), .Q ( signal_11270 ) ) ;
    buf_clk cell_5686 ( .C ( clk ), .D ( signal_11277 ), .Q ( signal_11278 ) ) ;
    buf_clk cell_5694 ( .C ( clk ), .D ( signal_11285 ), .Q ( signal_11286 ) ) ;
    buf_clk cell_5702 ( .C ( clk ), .D ( signal_11293 ), .Q ( signal_11294 ) ) ;
    buf_clk cell_5708 ( .C ( clk ), .D ( signal_11299 ), .Q ( signal_11300 ) ) ;
    buf_clk cell_5714 ( .C ( clk ), .D ( signal_11305 ), .Q ( signal_11306 ) ) ;
    buf_clk cell_5720 ( .C ( clk ), .D ( signal_11311 ), .Q ( signal_11312 ) ) ;
    buf_clk cell_5726 ( .C ( clk ), .D ( signal_11317 ), .Q ( signal_11318 ) ) ;
    buf_clk cell_5732 ( .C ( clk ), .D ( signal_11323 ), .Q ( signal_11324 ) ) ;
    buf_clk cell_5738 ( .C ( clk ), .D ( signal_11329 ), .Q ( signal_11330 ) ) ;
    buf_clk cell_5740 ( .C ( clk ), .D ( signal_11331 ), .Q ( signal_11332 ) ) ;
    buf_clk cell_5742 ( .C ( clk ), .D ( signal_11333 ), .Q ( signal_11334 ) ) ;
    buf_clk cell_5744 ( .C ( clk ), .D ( signal_11335 ), .Q ( signal_11336 ) ) ;
    buf_clk cell_5748 ( .C ( clk ), .D ( signal_11339 ), .Q ( signal_11340 ) ) ;
    buf_clk cell_5752 ( .C ( clk ), .D ( signal_11343 ), .Q ( signal_11344 ) ) ;
    buf_clk cell_5756 ( .C ( clk ), .D ( signal_11347 ), .Q ( signal_11348 ) ) ;
    buf_clk cell_5760 ( .C ( clk ), .D ( signal_11351 ), .Q ( signal_11352 ) ) ;
    buf_clk cell_5764 ( .C ( clk ), .D ( signal_11355 ), .Q ( signal_11356 ) ) ;
    buf_clk cell_5768 ( .C ( clk ), .D ( signal_11359 ), .Q ( signal_11360 ) ) ;
    buf_clk cell_5774 ( .C ( clk ), .D ( signal_11365 ), .Q ( signal_11366 ) ) ;
    buf_clk cell_5780 ( .C ( clk ), .D ( signal_11371 ), .Q ( signal_11372 ) ) ;
    buf_clk cell_5786 ( .C ( clk ), .D ( signal_11377 ), .Q ( signal_11378 ) ) ;
    buf_clk cell_5788 ( .C ( clk ), .D ( signal_11379 ), .Q ( signal_11380 ) ) ;
    buf_clk cell_5790 ( .C ( clk ), .D ( signal_11381 ), .Q ( signal_11382 ) ) ;
    buf_clk cell_5792 ( .C ( clk ), .D ( signal_11383 ), .Q ( signal_11384 ) ) ;
    buf_clk cell_5798 ( .C ( clk ), .D ( signal_11389 ), .Q ( signal_11390 ) ) ;
    buf_clk cell_5804 ( .C ( clk ), .D ( signal_11395 ), .Q ( signal_11396 ) ) ;
    buf_clk cell_5810 ( .C ( clk ), .D ( signal_11401 ), .Q ( signal_11402 ) ) ;
    buf_clk cell_5814 ( .C ( clk ), .D ( signal_11405 ), .Q ( signal_11406 ) ) ;
    buf_clk cell_5818 ( .C ( clk ), .D ( signal_11409 ), .Q ( signal_11410 ) ) ;
    buf_clk cell_5822 ( .C ( clk ), .D ( signal_11413 ), .Q ( signal_11414 ) ) ;
    buf_clk cell_5828 ( .C ( clk ), .D ( signal_11419 ), .Q ( signal_11420 ) ) ;
    buf_clk cell_5834 ( .C ( clk ), .D ( signal_11425 ), .Q ( signal_11426 ) ) ;
    buf_clk cell_5840 ( .C ( clk ), .D ( signal_11431 ), .Q ( signal_11432 ) ) ;
    buf_clk cell_5842 ( .C ( clk ), .D ( signal_11433 ), .Q ( signal_11434 ) ) ;
    buf_clk cell_5844 ( .C ( clk ), .D ( signal_11435 ), .Q ( signal_11436 ) ) ;
    buf_clk cell_5846 ( .C ( clk ), .D ( signal_11437 ), .Q ( signal_11438 ) ) ;
    buf_clk cell_5850 ( .C ( clk ), .D ( signal_11441 ), .Q ( signal_11442 ) ) ;
    buf_clk cell_5854 ( .C ( clk ), .D ( signal_11445 ), .Q ( signal_11446 ) ) ;
    buf_clk cell_5858 ( .C ( clk ), .D ( signal_11449 ), .Q ( signal_11450 ) ) ;
    buf_clk cell_5862 ( .C ( clk ), .D ( signal_11453 ), .Q ( signal_11454 ) ) ;
    buf_clk cell_5868 ( .C ( clk ), .D ( signal_11459 ), .Q ( signal_11460 ) ) ;
    buf_clk cell_5874 ( .C ( clk ), .D ( signal_11465 ), .Q ( signal_11466 ) ) ;
    buf_clk cell_5882 ( .C ( clk ), .D ( signal_11473 ), .Q ( signal_11474 ) ) ;
    buf_clk cell_5890 ( .C ( clk ), .D ( signal_11481 ), .Q ( signal_11482 ) ) ;
    buf_clk cell_5898 ( .C ( clk ), .D ( signal_11489 ), .Q ( signal_11490 ) ) ;
    buf_clk cell_5904 ( .C ( clk ), .D ( signal_11495 ), .Q ( signal_11496 ) ) ;
    buf_clk cell_5910 ( .C ( clk ), .D ( signal_11501 ), .Q ( signal_11502 ) ) ;
    buf_clk cell_5916 ( .C ( clk ), .D ( signal_11507 ), .Q ( signal_11508 ) ) ;
    buf_clk cell_5926 ( .C ( clk ), .D ( signal_11517 ), .Q ( signal_11518 ) ) ;
    buf_clk cell_5936 ( .C ( clk ), .D ( signal_11527 ), .Q ( signal_11528 ) ) ;
    buf_clk cell_5946 ( .C ( clk ), .D ( signal_11537 ), .Q ( signal_11538 ) ) ;
    buf_clk cell_5952 ( .C ( clk ), .D ( signal_11543 ), .Q ( signal_11544 ) ) ;
    buf_clk cell_5958 ( .C ( clk ), .D ( signal_11549 ), .Q ( signal_11550 ) ) ;
    buf_clk cell_5964 ( .C ( clk ), .D ( signal_11555 ), .Q ( signal_11556 ) ) ;
    buf_clk cell_5968 ( .C ( clk ), .D ( signal_11559 ), .Q ( signal_11560 ) ) ;
    buf_clk cell_5972 ( .C ( clk ), .D ( signal_11563 ), .Q ( signal_11564 ) ) ;
    buf_clk cell_5976 ( .C ( clk ), .D ( signal_11567 ), .Q ( signal_11568 ) ) ;
    buf_clk cell_5984 ( .C ( clk ), .D ( signal_11575 ), .Q ( signal_11576 ) ) ;
    buf_clk cell_5992 ( .C ( clk ), .D ( signal_11583 ), .Q ( signal_11584 ) ) ;
    buf_clk cell_6000 ( .C ( clk ), .D ( signal_11591 ), .Q ( signal_11592 ) ) ;
    buf_clk cell_6006 ( .C ( clk ), .D ( signal_11597 ), .Q ( signal_11598 ) ) ;
    buf_clk cell_6012 ( .C ( clk ), .D ( signal_11603 ), .Q ( signal_11604 ) ) ;
    buf_clk cell_6018 ( .C ( clk ), .D ( signal_11609 ), .Q ( signal_11610 ) ) ;
    buf_clk cell_6026 ( .C ( clk ), .D ( signal_11617 ), .Q ( signal_11618 ) ) ;
    buf_clk cell_6034 ( .C ( clk ), .D ( signal_11625 ), .Q ( signal_11626 ) ) ;
    buf_clk cell_6042 ( .C ( clk ), .D ( signal_11633 ), .Q ( signal_11634 ) ) ;
    buf_clk cell_6048 ( .C ( clk ), .D ( signal_11639 ), .Q ( signal_11640 ) ) ;
    buf_clk cell_6054 ( .C ( clk ), .D ( signal_11645 ), .Q ( signal_11646 ) ) ;
    buf_clk cell_6060 ( .C ( clk ), .D ( signal_11651 ), .Q ( signal_11652 ) ) ;
    buf_clk cell_6068 ( .C ( clk ), .D ( signal_11659 ), .Q ( signal_11660 ) ) ;
    buf_clk cell_6076 ( .C ( clk ), .D ( signal_11667 ), .Q ( signal_11668 ) ) ;
    buf_clk cell_6084 ( .C ( clk ), .D ( signal_11675 ), .Q ( signal_11676 ) ) ;
    buf_clk cell_6088 ( .C ( clk ), .D ( signal_11679 ), .Q ( signal_11680 ) ) ;
    buf_clk cell_6092 ( .C ( clk ), .D ( signal_11683 ), .Q ( signal_11684 ) ) ;
    buf_clk cell_6096 ( .C ( clk ), .D ( signal_11687 ), .Q ( signal_11688 ) ) ;
    buf_clk cell_6102 ( .C ( clk ), .D ( signal_11693 ), .Q ( signal_11694 ) ) ;
    buf_clk cell_6108 ( .C ( clk ), .D ( signal_11699 ), .Q ( signal_11700 ) ) ;
    buf_clk cell_6114 ( .C ( clk ), .D ( signal_11705 ), .Q ( signal_11706 ) ) ;
    buf_clk cell_6120 ( .C ( clk ), .D ( signal_11711 ), .Q ( signal_11712 ) ) ;
    buf_clk cell_6126 ( .C ( clk ), .D ( signal_11717 ), .Q ( signal_11718 ) ) ;
    buf_clk cell_6132 ( .C ( clk ), .D ( signal_11723 ), .Q ( signal_11724 ) ) ;
    buf_clk cell_6136 ( .C ( clk ), .D ( signal_11727 ), .Q ( signal_11728 ) ) ;
    buf_clk cell_6140 ( .C ( clk ), .D ( signal_11731 ), .Q ( signal_11732 ) ) ;
    buf_clk cell_6144 ( .C ( clk ), .D ( signal_11735 ), .Q ( signal_11736 ) ) ;
    buf_clk cell_6148 ( .C ( clk ), .D ( signal_11739 ), .Q ( signal_11740 ) ) ;
    buf_clk cell_6152 ( .C ( clk ), .D ( signal_11743 ), .Q ( signal_11744 ) ) ;
    buf_clk cell_6156 ( .C ( clk ), .D ( signal_11747 ), .Q ( signal_11748 ) ) ;
    buf_clk cell_6162 ( .C ( clk ), .D ( signal_11753 ), .Q ( signal_11754 ) ) ;
    buf_clk cell_6170 ( .C ( clk ), .D ( signal_11761 ), .Q ( signal_11762 ) ) ;
    buf_clk cell_6178 ( .C ( clk ), .D ( signal_11769 ), .Q ( signal_11770 ) ) ;
    buf_clk cell_6190 ( .C ( clk ), .D ( signal_11781 ), .Q ( signal_11782 ) ) ;
    buf_clk cell_6202 ( .C ( clk ), .D ( signal_11793 ), .Q ( signal_11794 ) ) ;
    buf_clk cell_6214 ( .C ( clk ), .D ( signal_11805 ), .Q ( signal_11806 ) ) ;
    buf_clk cell_6220 ( .C ( clk ), .D ( signal_11811 ), .Q ( signal_11812 ) ) ;
    buf_clk cell_6226 ( .C ( clk ), .D ( signal_11817 ), .Q ( signal_11818 ) ) ;
    buf_clk cell_6232 ( .C ( clk ), .D ( signal_11823 ), .Q ( signal_11824 ) ) ;
    buf_clk cell_6238 ( .C ( clk ), .D ( signal_11829 ), .Q ( signal_11830 ) ) ;
    buf_clk cell_6244 ( .C ( clk ), .D ( signal_11835 ), .Q ( signal_11836 ) ) ;
    buf_clk cell_6250 ( .C ( clk ), .D ( signal_11841 ), .Q ( signal_11842 ) ) ;
    buf_clk cell_6264 ( .C ( clk ), .D ( signal_11855 ), .Q ( signal_11856 ) ) ;
    buf_clk cell_6278 ( .C ( clk ), .D ( signal_11869 ), .Q ( signal_11870 ) ) ;
    buf_clk cell_6292 ( .C ( clk ), .D ( signal_11883 ), .Q ( signal_11884 ) ) ;
    buf_clk cell_6300 ( .C ( clk ), .D ( signal_11891 ), .Q ( signal_11892 ) ) ;
    buf_clk cell_6308 ( .C ( clk ), .D ( signal_11899 ), .Q ( signal_11900 ) ) ;
    buf_clk cell_6316 ( .C ( clk ), .D ( signal_11907 ), .Q ( signal_11908 ) ) ;
    buf_clk cell_6330 ( .C ( clk ), .D ( signal_11921 ), .Q ( signal_11922 ) ) ;
    buf_clk cell_6344 ( .C ( clk ), .D ( signal_11935 ), .Q ( signal_11936 ) ) ;
    buf_clk cell_6358 ( .C ( clk ), .D ( signal_11949 ), .Q ( signal_11950 ) ) ;
    buf_clk cell_6366 ( .C ( clk ), .D ( signal_11957 ), .Q ( signal_11958 ) ) ;
    buf_clk cell_6374 ( .C ( clk ), .D ( signal_11965 ), .Q ( signal_11966 ) ) ;
    buf_clk cell_6382 ( .C ( clk ), .D ( signal_11973 ), .Q ( signal_11974 ) ) ;
    buf_clk cell_6402 ( .C ( clk ), .D ( signal_11993 ), .Q ( signal_11994 ) ) ;
    buf_clk cell_6412 ( .C ( clk ), .D ( signal_12003 ), .Q ( signal_12004 ) ) ;
    buf_clk cell_6422 ( .C ( clk ), .D ( signal_12013 ), .Q ( signal_12014 ) ) ;
    buf_clk cell_6450 ( .C ( clk ), .D ( signal_12041 ), .Q ( signal_12042 ) ) ;
    buf_clk cell_6466 ( .C ( clk ), .D ( signal_12057 ), .Q ( signal_12058 ) ) ;
    buf_clk cell_6482 ( .C ( clk ), .D ( signal_12073 ), .Q ( signal_12074 ) ) ;
    buf_clk cell_6510 ( .C ( clk ), .D ( signal_12101 ), .Q ( signal_12102 ) ) ;
    buf_clk cell_6526 ( .C ( clk ), .D ( signal_12117 ), .Q ( signal_12118 ) ) ;
    buf_clk cell_6542 ( .C ( clk ), .D ( signal_12133 ), .Q ( signal_12134 ) ) ;
    buf_clk cell_6552 ( .C ( clk ), .D ( signal_12143 ), .Q ( signal_12144 ) ) ;
    buf_clk cell_6562 ( .C ( clk ), .D ( signal_12153 ), .Q ( signal_12154 ) ) ;
    buf_clk cell_6572 ( .C ( clk ), .D ( signal_12163 ), .Q ( signal_12164 ) ) ;
    buf_clk cell_6610 ( .C ( clk ), .D ( signal_12201 ), .Q ( signal_12202 ) ) ;
    buf_clk cell_6620 ( .C ( clk ), .D ( signal_12211 ), .Q ( signal_12212 ) ) ;
    buf_clk cell_6630 ( .C ( clk ), .D ( signal_12221 ), .Q ( signal_12222 ) ) ;
    buf_clk cell_6658 ( .C ( clk ), .D ( signal_12249 ), .Q ( signal_12250 ) ) ;
    buf_clk cell_6668 ( .C ( clk ), .D ( signal_12259 ), .Q ( signal_12260 ) ) ;
    buf_clk cell_6678 ( .C ( clk ), .D ( signal_12269 ), .Q ( signal_12270 ) ) ;
    buf_clk cell_6694 ( .C ( clk ), .D ( signal_12285 ), .Q ( signal_12286 ) ) ;
    buf_clk cell_6710 ( .C ( clk ), .D ( signal_12301 ), .Q ( signal_12302 ) ) ;
    buf_clk cell_6726 ( .C ( clk ), .D ( signal_12317 ), .Q ( signal_12318 ) ) ;
    buf_clk cell_6744 ( .C ( clk ), .D ( signal_12335 ), .Q ( signal_12336 ) ) ;
    buf_clk cell_6762 ( .C ( clk ), .D ( signal_12353 ), .Q ( signal_12354 ) ) ;
    buf_clk cell_6780 ( .C ( clk ), .D ( signal_12371 ), .Q ( signal_12372 ) ) ;
    buf_clk cell_6894 ( .C ( clk ), .D ( signal_12485 ), .Q ( signal_12486 ) ) ;
    buf_clk cell_6914 ( .C ( clk ), .D ( signal_12505 ), .Q ( signal_12506 ) ) ;
    buf_clk cell_6934 ( .C ( clk ), .D ( signal_12525 ), .Q ( signal_12526 ) ) ;

    /* cells in depth 17 */
    buf_clk cell_5863 ( .C ( clk ), .D ( signal_11454 ), .Q ( signal_11455 ) ) ;
    buf_clk cell_5869 ( .C ( clk ), .D ( signal_11460 ), .Q ( signal_11461 ) ) ;
    buf_clk cell_5875 ( .C ( clk ), .D ( signal_11466 ), .Q ( signal_11467 ) ) ;
    buf_clk cell_5883 ( .C ( clk ), .D ( signal_11474 ), .Q ( signal_11475 ) ) ;
    buf_clk cell_5891 ( .C ( clk ), .D ( signal_11482 ), .Q ( signal_11483 ) ) ;
    buf_clk cell_5899 ( .C ( clk ), .D ( signal_11490 ), .Q ( signal_11491 ) ) ;
    buf_clk cell_5905 ( .C ( clk ), .D ( signal_11496 ), .Q ( signal_11497 ) ) ;
    buf_clk cell_5911 ( .C ( clk ), .D ( signal_11502 ), .Q ( signal_11503 ) ) ;
    buf_clk cell_5917 ( .C ( clk ), .D ( signal_11508 ), .Q ( signal_11509 ) ) ;
    buf_clk cell_5927 ( .C ( clk ), .D ( signal_11518 ), .Q ( signal_11519 ) ) ;
    buf_clk cell_5937 ( .C ( clk ), .D ( signal_11528 ), .Q ( signal_11529 ) ) ;
    buf_clk cell_5947 ( .C ( clk ), .D ( signal_11538 ), .Q ( signal_11539 ) ) ;
    buf_clk cell_5953 ( .C ( clk ), .D ( signal_11544 ), .Q ( signal_11545 ) ) ;
    buf_clk cell_5959 ( .C ( clk ), .D ( signal_11550 ), .Q ( signal_11551 ) ) ;
    buf_clk cell_5965 ( .C ( clk ), .D ( signal_11556 ), .Q ( signal_11557 ) ) ;
    buf_clk cell_5969 ( .C ( clk ), .D ( signal_11560 ), .Q ( signal_11561 ) ) ;
    buf_clk cell_5973 ( .C ( clk ), .D ( signal_11564 ), .Q ( signal_11565 ) ) ;
    buf_clk cell_5977 ( .C ( clk ), .D ( signal_11568 ), .Q ( signal_11569 ) ) ;
    buf_clk cell_5985 ( .C ( clk ), .D ( signal_11576 ), .Q ( signal_11577 ) ) ;
    buf_clk cell_5993 ( .C ( clk ), .D ( signal_11584 ), .Q ( signal_11585 ) ) ;
    buf_clk cell_6001 ( .C ( clk ), .D ( signal_11592 ), .Q ( signal_11593 ) ) ;
    buf_clk cell_6007 ( .C ( clk ), .D ( signal_11598 ), .Q ( signal_11599 ) ) ;
    buf_clk cell_6013 ( .C ( clk ), .D ( signal_11604 ), .Q ( signal_11605 ) ) ;
    buf_clk cell_6019 ( .C ( clk ), .D ( signal_11610 ), .Q ( signal_11611 ) ) ;
    buf_clk cell_6027 ( .C ( clk ), .D ( signal_11618 ), .Q ( signal_11619 ) ) ;
    buf_clk cell_6035 ( .C ( clk ), .D ( signal_11626 ), .Q ( signal_11627 ) ) ;
    buf_clk cell_6043 ( .C ( clk ), .D ( signal_11634 ), .Q ( signal_11635 ) ) ;
    buf_clk cell_6049 ( .C ( clk ), .D ( signal_11640 ), .Q ( signal_11641 ) ) ;
    buf_clk cell_6055 ( .C ( clk ), .D ( signal_11646 ), .Q ( signal_11647 ) ) ;
    buf_clk cell_6061 ( .C ( clk ), .D ( signal_11652 ), .Q ( signal_11653 ) ) ;
    buf_clk cell_6069 ( .C ( clk ), .D ( signal_11660 ), .Q ( signal_11661 ) ) ;
    buf_clk cell_6077 ( .C ( clk ), .D ( signal_11668 ), .Q ( signal_11669 ) ) ;
    buf_clk cell_6085 ( .C ( clk ), .D ( signal_11676 ), .Q ( signal_11677 ) ) ;
    buf_clk cell_6089 ( .C ( clk ), .D ( signal_11680 ), .Q ( signal_11681 ) ) ;
    buf_clk cell_6093 ( .C ( clk ), .D ( signal_11684 ), .Q ( signal_11685 ) ) ;
    buf_clk cell_6097 ( .C ( clk ), .D ( signal_11688 ), .Q ( signal_11689 ) ) ;
    buf_clk cell_6103 ( .C ( clk ), .D ( signal_11694 ), .Q ( signal_11695 ) ) ;
    buf_clk cell_6109 ( .C ( clk ), .D ( signal_11700 ), .Q ( signal_11701 ) ) ;
    buf_clk cell_6115 ( .C ( clk ), .D ( signal_11706 ), .Q ( signal_11707 ) ) ;
    buf_clk cell_6121 ( .C ( clk ), .D ( signal_11712 ), .Q ( signal_11713 ) ) ;
    buf_clk cell_6127 ( .C ( clk ), .D ( signal_11718 ), .Q ( signal_11719 ) ) ;
    buf_clk cell_6133 ( .C ( clk ), .D ( signal_11724 ), .Q ( signal_11725 ) ) ;
    buf_clk cell_6137 ( .C ( clk ), .D ( signal_11728 ), .Q ( signal_11729 ) ) ;
    buf_clk cell_6141 ( .C ( clk ), .D ( signal_11732 ), .Q ( signal_11733 ) ) ;
    buf_clk cell_6145 ( .C ( clk ), .D ( signal_11736 ), .Q ( signal_11737 ) ) ;
    buf_clk cell_6149 ( .C ( clk ), .D ( signal_11740 ), .Q ( signal_11741 ) ) ;
    buf_clk cell_6153 ( .C ( clk ), .D ( signal_11744 ), .Q ( signal_11745 ) ) ;
    buf_clk cell_6157 ( .C ( clk ), .D ( signal_11748 ), .Q ( signal_11749 ) ) ;
    buf_clk cell_6163 ( .C ( clk ), .D ( signal_11754 ), .Q ( signal_11755 ) ) ;
    buf_clk cell_6171 ( .C ( clk ), .D ( signal_11762 ), .Q ( signal_11763 ) ) ;
    buf_clk cell_6179 ( .C ( clk ), .D ( signal_11770 ), .Q ( signal_11771 ) ) ;
    buf_clk cell_6191 ( .C ( clk ), .D ( signal_11782 ), .Q ( signal_11783 ) ) ;
    buf_clk cell_6203 ( .C ( clk ), .D ( signal_11794 ), .Q ( signal_11795 ) ) ;
    buf_clk cell_6215 ( .C ( clk ), .D ( signal_11806 ), .Q ( signal_11807 ) ) ;
    buf_clk cell_6221 ( .C ( clk ), .D ( signal_11812 ), .Q ( signal_11813 ) ) ;
    buf_clk cell_6227 ( .C ( clk ), .D ( signal_11818 ), .Q ( signal_11819 ) ) ;
    buf_clk cell_6233 ( .C ( clk ), .D ( signal_11824 ), .Q ( signal_11825 ) ) ;
    buf_clk cell_6239 ( .C ( clk ), .D ( signal_11830 ), .Q ( signal_11831 ) ) ;
    buf_clk cell_6245 ( .C ( clk ), .D ( signal_11836 ), .Q ( signal_11837 ) ) ;
    buf_clk cell_6251 ( .C ( clk ), .D ( signal_11842 ), .Q ( signal_11843 ) ) ;
    buf_clk cell_6265 ( .C ( clk ), .D ( signal_11856 ), .Q ( signal_11857 ) ) ;
    buf_clk cell_6279 ( .C ( clk ), .D ( signal_11870 ), .Q ( signal_11871 ) ) ;
    buf_clk cell_6293 ( .C ( clk ), .D ( signal_11884 ), .Q ( signal_11885 ) ) ;
    buf_clk cell_6301 ( .C ( clk ), .D ( signal_11892 ), .Q ( signal_11893 ) ) ;
    buf_clk cell_6309 ( .C ( clk ), .D ( signal_11900 ), .Q ( signal_11901 ) ) ;
    buf_clk cell_6317 ( .C ( clk ), .D ( signal_11908 ), .Q ( signal_11909 ) ) ;
    buf_clk cell_6331 ( .C ( clk ), .D ( signal_11922 ), .Q ( signal_11923 ) ) ;
    buf_clk cell_6345 ( .C ( clk ), .D ( signal_11936 ), .Q ( signal_11937 ) ) ;
    buf_clk cell_6359 ( .C ( clk ), .D ( signal_11950 ), .Q ( signal_11951 ) ) ;
    buf_clk cell_6367 ( .C ( clk ), .D ( signal_11958 ), .Q ( signal_11959 ) ) ;
    buf_clk cell_6375 ( .C ( clk ), .D ( signal_11966 ), .Q ( signal_11967 ) ) ;
    buf_clk cell_6383 ( .C ( clk ), .D ( signal_11974 ), .Q ( signal_11975 ) ) ;
    buf_clk cell_6403 ( .C ( clk ), .D ( signal_11994 ), .Q ( signal_11995 ) ) ;
    buf_clk cell_6413 ( .C ( clk ), .D ( signal_12004 ), .Q ( signal_12005 ) ) ;
    buf_clk cell_6423 ( .C ( clk ), .D ( signal_12014 ), .Q ( signal_12015 ) ) ;
    buf_clk cell_6451 ( .C ( clk ), .D ( signal_12042 ), .Q ( signal_12043 ) ) ;
    buf_clk cell_6467 ( .C ( clk ), .D ( signal_12058 ), .Q ( signal_12059 ) ) ;
    buf_clk cell_6483 ( .C ( clk ), .D ( signal_12074 ), .Q ( signal_12075 ) ) ;
    buf_clk cell_6511 ( .C ( clk ), .D ( signal_12102 ), .Q ( signal_12103 ) ) ;
    buf_clk cell_6527 ( .C ( clk ), .D ( signal_12118 ), .Q ( signal_12119 ) ) ;
    buf_clk cell_6543 ( .C ( clk ), .D ( signal_12134 ), .Q ( signal_12135 ) ) ;
    buf_clk cell_6553 ( .C ( clk ), .D ( signal_12144 ), .Q ( signal_12145 ) ) ;
    buf_clk cell_6563 ( .C ( clk ), .D ( signal_12154 ), .Q ( signal_12155 ) ) ;
    buf_clk cell_6573 ( .C ( clk ), .D ( signal_12164 ), .Q ( signal_12165 ) ) ;
    buf_clk cell_6611 ( .C ( clk ), .D ( signal_12202 ), .Q ( signal_12203 ) ) ;
    buf_clk cell_6621 ( .C ( clk ), .D ( signal_12212 ), .Q ( signal_12213 ) ) ;
    buf_clk cell_6631 ( .C ( clk ), .D ( signal_12222 ), .Q ( signal_12223 ) ) ;
    buf_clk cell_6659 ( .C ( clk ), .D ( signal_12250 ), .Q ( signal_12251 ) ) ;
    buf_clk cell_6669 ( .C ( clk ), .D ( signal_12260 ), .Q ( signal_12261 ) ) ;
    buf_clk cell_6679 ( .C ( clk ), .D ( signal_12270 ), .Q ( signal_12271 ) ) ;
    buf_clk cell_6695 ( .C ( clk ), .D ( signal_12286 ), .Q ( signal_12287 ) ) ;
    buf_clk cell_6711 ( .C ( clk ), .D ( signal_12302 ), .Q ( signal_12303 ) ) ;
    buf_clk cell_6727 ( .C ( clk ), .D ( signal_12318 ), .Q ( signal_12319 ) ) ;
    buf_clk cell_6745 ( .C ( clk ), .D ( signal_12336 ), .Q ( signal_12337 ) ) ;
    buf_clk cell_6763 ( .C ( clk ), .D ( signal_12354 ), .Q ( signal_12355 ) ) ;
    buf_clk cell_6781 ( .C ( clk ), .D ( signal_12372 ), .Q ( signal_12373 ) ) ;
    buf_clk cell_6801 ( .C ( clk ), .D ( signal_2281 ), .Q ( signal_12393 ) ) ;
    buf_clk cell_6809 ( .C ( clk ), .D ( signal_5086 ), .Q ( signal_12401 ) ) ;
    buf_clk cell_6817 ( .C ( clk ), .D ( signal_5087 ), .Q ( signal_12409 ) ) ;
    buf_clk cell_6895 ( .C ( clk ), .D ( signal_12486 ), .Q ( signal_12487 ) ) ;
    buf_clk cell_6915 ( .C ( clk ), .D ( signal_12506 ), .Q ( signal_12507 ) ) ;
    buf_clk cell_6935 ( .C ( clk ), .D ( signal_12526 ), .Q ( signal_12527 ) ) ;
    buf_clk cell_6969 ( .C ( clk ), .D ( signal_2260 ), .Q ( signal_12561 ) ) ;
    buf_clk cell_6981 ( .C ( clk ), .D ( signal_5044 ), .Q ( signal_12573 ) ) ;
    buf_clk cell_6993 ( .C ( clk ), .D ( signal_5045 ), .Q ( signal_12585 ) ) ;
    buf_clk cell_7005 ( .C ( clk ), .D ( signal_2322 ), .Q ( signal_12597 ) ) ;
    buf_clk cell_7019 ( .C ( clk ), .D ( signal_5168 ), .Q ( signal_12611 ) ) ;
    buf_clk cell_7033 ( .C ( clk ), .D ( signal_5169 ), .Q ( signal_12625 ) ) ;

    /* cells in depth 18 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2230 ( .a ({signal_11078, signal_11072, signal_11066}), .b ({signal_4917, signal_4916, signal_2196}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403]}), .c ({signal_5015, signal_5014, signal_2245}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2231 ( .a ({signal_11102, signal_11094, signal_11086}), .b ({signal_4919, signal_4918, signal_2197}), .clk ( clk ), .r ({Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({signal_5017, signal_5016, signal_2246}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2232 ( .a ({signal_11120, signal_11114, signal_11108}), .b ({signal_4921, signal_4920, signal_2198}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409]}), .c ({signal_5019, signal_5018, signal_2247}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2267 ( .a ({signal_11138, signal_11132, signal_11126}), .b ({signal_5007, signal_5006, signal_2241}), .clk ( clk ), .r ({Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({signal_5089, signal_5088, signal_2282}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2268 ( .a ({signal_11162, signal_11154, signal_11146}), .b ({signal_4953, signal_4952, signal_2214}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415]}), .c ({signal_5091, signal_5090, signal_2283}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2281 ( .a ({signal_5091, signal_5090, signal_2283}), .b ({signal_5117, signal_5116, signal_2296}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2284 ( .a ({signal_11192, signal_11182, signal_11172}), .b ({signal_5049, signal_5048, signal_2262}), .clk ( clk ), .r ({Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({signal_5123, signal_5122, signal_2299}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2289 ( .a ({signal_11198, signal_11196, signal_11194}), .b ({signal_5043, signal_5042, signal_2259}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421]}), .c ({signal_5133, signal_5132, signal_2304}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2291 ( .a ({signal_11216, signal_11210, signal_11204}), .b ({signal_5065, signal_5064, signal_2270}), .clk ( clk ), .r ({Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({signal_5137, signal_5136, signal_2306}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2292 ( .a ({signal_11240, signal_11232, signal_11224}), .b ({signal_5071, signal_5070, signal_2273}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427]}), .c ({signal_5139, signal_5138, signal_2307}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2293 ( .a ({signal_11270, signal_11260, signal_11250}), .b ({signal_5075, signal_5074, signal_2275}), .clk ( clk ), .r ({Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_5141, signal_5140, signal_2308}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2294 ( .a ({signal_11294, signal_11286, signal_11278}), .b ({signal_5081, signal_5080, signal_2278}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433]}), .c ({signal_5143, signal_5142, signal_2309}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2295 ( .a ({signal_11312, signal_11306, signal_11300}), .b ({signal_5047, signal_5046, signal_2261}), .clk ( clk ), .r ({Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({signal_5145, signal_5144, signal_2310}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2298 ( .a ({signal_5123, signal_5122, signal_2299}), .b ({signal_5151, signal_5150, signal_2313}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2300 ( .a ({signal_5133, signal_5132, signal_2304}), .b ({signal_5155, signal_5154, signal_2315}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2302 ( .a ({signal_5143, signal_5142, signal_2309}), .b ({signal_5159, signal_5158, signal_2317}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2303 ( .a ({signal_5145, signal_5144, signal_2310}), .b ({signal_5161, signal_5160, signal_2318}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2308 ( .a ({signal_11330, signal_11324, signal_11318}), .b ({signal_5105, signal_5104, signal_2290}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439]}), .c ({signal_5171, signal_5170, signal_2323}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2309 ( .a ({signal_11336, signal_11334, signal_11332}), .b ({signal_5107, signal_5106, signal_2291}), .clk ( clk ), .r ({Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({signal_5173, signal_5172, signal_2324}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2310 ( .a ({signal_11336, signal_11334, signal_11332}), .b ({signal_5109, signal_5108, signal_2292}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445]}), .c ({signal_5175, signal_5174, signal_2325}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2311 ( .a ({signal_11348, signal_11344, signal_11340}), .b ({signal_5111, signal_5110, signal_2293}), .clk ( clk ), .r ({Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({signal_5177, signal_5176, signal_2326}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2312 ( .a ({signal_11360, signal_11356, signal_11352}), .b ({signal_5113, signal_5112, signal_2294}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451]}), .c ({signal_5179, signal_5178, signal_2327}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2313 ( .a ({signal_5129, signal_5128, signal_2302}), .b ({signal_5083, signal_5082, signal_2279}), .clk ( clk ), .r ({Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({signal_5181, signal_5180, signal_2328}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2314 ( .a ({signal_11378, signal_11372, signal_11366}), .b ({signal_5115, signal_5114, signal_2295}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457]}), .c ({signal_5183, signal_5182, signal_2329}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2315 ( .a ({signal_11384, signal_11382, signal_11380}), .b ({signal_5011, signal_5010, signal_2243}), .clk ( clk ), .r ({Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_5185, signal_5184, signal_2330}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2320 ( .a ({signal_5171, signal_5170, signal_2323}), .b ({signal_5195, signal_5194, signal_2335}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2321 ( .a ({signal_5173, signal_5172, signal_2324}), .b ({signal_5197, signal_5196, signal_2336}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2322 ( .a ({signal_5175, signal_5174, signal_2325}), .b ({signal_5199, signal_5198, signal_2337}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2323 ( .a ({signal_5177, signal_5176, signal_2326}), .b ({signal_5201, signal_5200, signal_2338}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2324 ( .a ({signal_11402, signal_11396, signal_11390}), .b ({signal_5163, signal_5162, signal_2319}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463]}), .c ({signal_5203, signal_5202, signal_2339}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2326 ( .a ({signal_11414, signal_11410, signal_11406}), .b ({signal_5153, signal_5152, signal_2314}), .clk ( clk ), .r ({Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({signal_5207, signal_5206, signal_2341}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2328 ( .a ({signal_11432, signal_11426, signal_11420}), .b ({signal_5165, signal_5164, signal_2320}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469]}), .c ({signal_5211, signal_5210, signal_2343}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2329 ( .a ({signal_11438, signal_11436, signal_11434}), .b ({signal_5167, signal_5166, signal_2321}), .clk ( clk ), .r ({Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({signal_5213, signal_5212, signal_2344}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2330 ( .a ({signal_11450, signal_11446, signal_11442}), .b ({signal_5157, signal_5156, signal_2316}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475]}), .c ({signal_5215, signal_5214, signal_2345}) ) ;
    buf_clk cell_5864 ( .C ( clk ), .D ( signal_11455 ), .Q ( signal_11456 ) ) ;
    buf_clk cell_5870 ( .C ( clk ), .D ( signal_11461 ), .Q ( signal_11462 ) ) ;
    buf_clk cell_5876 ( .C ( clk ), .D ( signal_11467 ), .Q ( signal_11468 ) ) ;
    buf_clk cell_5884 ( .C ( clk ), .D ( signal_11475 ), .Q ( signal_11476 ) ) ;
    buf_clk cell_5892 ( .C ( clk ), .D ( signal_11483 ), .Q ( signal_11484 ) ) ;
    buf_clk cell_5900 ( .C ( clk ), .D ( signal_11491 ), .Q ( signal_11492 ) ) ;
    buf_clk cell_5906 ( .C ( clk ), .D ( signal_11497 ), .Q ( signal_11498 ) ) ;
    buf_clk cell_5912 ( .C ( clk ), .D ( signal_11503 ), .Q ( signal_11504 ) ) ;
    buf_clk cell_5918 ( .C ( clk ), .D ( signal_11509 ), .Q ( signal_11510 ) ) ;
    buf_clk cell_5928 ( .C ( clk ), .D ( signal_11519 ), .Q ( signal_11520 ) ) ;
    buf_clk cell_5938 ( .C ( clk ), .D ( signal_11529 ), .Q ( signal_11530 ) ) ;
    buf_clk cell_5948 ( .C ( clk ), .D ( signal_11539 ), .Q ( signal_11540 ) ) ;
    buf_clk cell_5954 ( .C ( clk ), .D ( signal_11545 ), .Q ( signal_11546 ) ) ;
    buf_clk cell_5960 ( .C ( clk ), .D ( signal_11551 ), .Q ( signal_11552 ) ) ;
    buf_clk cell_5966 ( .C ( clk ), .D ( signal_11557 ), .Q ( signal_11558 ) ) ;
    buf_clk cell_5970 ( .C ( clk ), .D ( signal_11561 ), .Q ( signal_11562 ) ) ;
    buf_clk cell_5974 ( .C ( clk ), .D ( signal_11565 ), .Q ( signal_11566 ) ) ;
    buf_clk cell_5978 ( .C ( clk ), .D ( signal_11569 ), .Q ( signal_11570 ) ) ;
    buf_clk cell_5986 ( .C ( clk ), .D ( signal_11577 ), .Q ( signal_11578 ) ) ;
    buf_clk cell_5994 ( .C ( clk ), .D ( signal_11585 ), .Q ( signal_11586 ) ) ;
    buf_clk cell_6002 ( .C ( clk ), .D ( signal_11593 ), .Q ( signal_11594 ) ) ;
    buf_clk cell_6008 ( .C ( clk ), .D ( signal_11599 ), .Q ( signal_11600 ) ) ;
    buf_clk cell_6014 ( .C ( clk ), .D ( signal_11605 ), .Q ( signal_11606 ) ) ;
    buf_clk cell_6020 ( .C ( clk ), .D ( signal_11611 ), .Q ( signal_11612 ) ) ;
    buf_clk cell_6028 ( .C ( clk ), .D ( signal_11619 ), .Q ( signal_11620 ) ) ;
    buf_clk cell_6036 ( .C ( clk ), .D ( signal_11627 ), .Q ( signal_11628 ) ) ;
    buf_clk cell_6044 ( .C ( clk ), .D ( signal_11635 ), .Q ( signal_11636 ) ) ;
    buf_clk cell_6050 ( .C ( clk ), .D ( signal_11641 ), .Q ( signal_11642 ) ) ;
    buf_clk cell_6056 ( .C ( clk ), .D ( signal_11647 ), .Q ( signal_11648 ) ) ;
    buf_clk cell_6062 ( .C ( clk ), .D ( signal_11653 ), .Q ( signal_11654 ) ) ;
    buf_clk cell_6070 ( .C ( clk ), .D ( signal_11661 ), .Q ( signal_11662 ) ) ;
    buf_clk cell_6078 ( .C ( clk ), .D ( signal_11669 ), .Q ( signal_11670 ) ) ;
    buf_clk cell_6086 ( .C ( clk ), .D ( signal_11677 ), .Q ( signal_11678 ) ) ;
    buf_clk cell_6090 ( .C ( clk ), .D ( signal_11681 ), .Q ( signal_11682 ) ) ;
    buf_clk cell_6094 ( .C ( clk ), .D ( signal_11685 ), .Q ( signal_11686 ) ) ;
    buf_clk cell_6098 ( .C ( clk ), .D ( signal_11689 ), .Q ( signal_11690 ) ) ;
    buf_clk cell_6104 ( .C ( clk ), .D ( signal_11695 ), .Q ( signal_11696 ) ) ;
    buf_clk cell_6110 ( .C ( clk ), .D ( signal_11701 ), .Q ( signal_11702 ) ) ;
    buf_clk cell_6116 ( .C ( clk ), .D ( signal_11707 ), .Q ( signal_11708 ) ) ;
    buf_clk cell_6122 ( .C ( clk ), .D ( signal_11713 ), .Q ( signal_11714 ) ) ;
    buf_clk cell_6128 ( .C ( clk ), .D ( signal_11719 ), .Q ( signal_11720 ) ) ;
    buf_clk cell_6134 ( .C ( clk ), .D ( signal_11725 ), .Q ( signal_11726 ) ) ;
    buf_clk cell_6138 ( .C ( clk ), .D ( signal_11729 ), .Q ( signal_11730 ) ) ;
    buf_clk cell_6142 ( .C ( clk ), .D ( signal_11733 ), .Q ( signal_11734 ) ) ;
    buf_clk cell_6146 ( .C ( clk ), .D ( signal_11737 ), .Q ( signal_11738 ) ) ;
    buf_clk cell_6150 ( .C ( clk ), .D ( signal_11741 ), .Q ( signal_11742 ) ) ;
    buf_clk cell_6154 ( .C ( clk ), .D ( signal_11745 ), .Q ( signal_11746 ) ) ;
    buf_clk cell_6158 ( .C ( clk ), .D ( signal_11749 ), .Q ( signal_11750 ) ) ;
    buf_clk cell_6164 ( .C ( clk ), .D ( signal_11755 ), .Q ( signal_11756 ) ) ;
    buf_clk cell_6172 ( .C ( clk ), .D ( signal_11763 ), .Q ( signal_11764 ) ) ;
    buf_clk cell_6180 ( .C ( clk ), .D ( signal_11771 ), .Q ( signal_11772 ) ) ;
    buf_clk cell_6192 ( .C ( clk ), .D ( signal_11783 ), .Q ( signal_11784 ) ) ;
    buf_clk cell_6204 ( .C ( clk ), .D ( signal_11795 ), .Q ( signal_11796 ) ) ;
    buf_clk cell_6216 ( .C ( clk ), .D ( signal_11807 ), .Q ( signal_11808 ) ) ;
    buf_clk cell_6222 ( .C ( clk ), .D ( signal_11813 ), .Q ( signal_11814 ) ) ;
    buf_clk cell_6228 ( .C ( clk ), .D ( signal_11819 ), .Q ( signal_11820 ) ) ;
    buf_clk cell_6234 ( .C ( clk ), .D ( signal_11825 ), .Q ( signal_11826 ) ) ;
    buf_clk cell_6240 ( .C ( clk ), .D ( signal_11831 ), .Q ( signal_11832 ) ) ;
    buf_clk cell_6246 ( .C ( clk ), .D ( signal_11837 ), .Q ( signal_11838 ) ) ;
    buf_clk cell_6252 ( .C ( clk ), .D ( signal_11843 ), .Q ( signal_11844 ) ) ;
    buf_clk cell_6266 ( .C ( clk ), .D ( signal_11857 ), .Q ( signal_11858 ) ) ;
    buf_clk cell_6280 ( .C ( clk ), .D ( signal_11871 ), .Q ( signal_11872 ) ) ;
    buf_clk cell_6294 ( .C ( clk ), .D ( signal_11885 ), .Q ( signal_11886 ) ) ;
    buf_clk cell_6302 ( .C ( clk ), .D ( signal_11893 ), .Q ( signal_11894 ) ) ;
    buf_clk cell_6310 ( .C ( clk ), .D ( signal_11901 ), .Q ( signal_11902 ) ) ;
    buf_clk cell_6318 ( .C ( clk ), .D ( signal_11909 ), .Q ( signal_11910 ) ) ;
    buf_clk cell_6332 ( .C ( clk ), .D ( signal_11923 ), .Q ( signal_11924 ) ) ;
    buf_clk cell_6346 ( .C ( clk ), .D ( signal_11937 ), .Q ( signal_11938 ) ) ;
    buf_clk cell_6360 ( .C ( clk ), .D ( signal_11951 ), .Q ( signal_11952 ) ) ;
    buf_clk cell_6368 ( .C ( clk ), .D ( signal_11959 ), .Q ( signal_11960 ) ) ;
    buf_clk cell_6376 ( .C ( clk ), .D ( signal_11967 ), .Q ( signal_11968 ) ) ;
    buf_clk cell_6384 ( .C ( clk ), .D ( signal_11975 ), .Q ( signal_11976 ) ) ;
    buf_clk cell_6404 ( .C ( clk ), .D ( signal_11995 ), .Q ( signal_11996 ) ) ;
    buf_clk cell_6414 ( .C ( clk ), .D ( signal_12005 ), .Q ( signal_12006 ) ) ;
    buf_clk cell_6424 ( .C ( clk ), .D ( signal_12015 ), .Q ( signal_12016 ) ) ;
    buf_clk cell_6452 ( .C ( clk ), .D ( signal_12043 ), .Q ( signal_12044 ) ) ;
    buf_clk cell_6468 ( .C ( clk ), .D ( signal_12059 ), .Q ( signal_12060 ) ) ;
    buf_clk cell_6484 ( .C ( clk ), .D ( signal_12075 ), .Q ( signal_12076 ) ) ;
    buf_clk cell_6512 ( .C ( clk ), .D ( signal_12103 ), .Q ( signal_12104 ) ) ;
    buf_clk cell_6528 ( .C ( clk ), .D ( signal_12119 ), .Q ( signal_12120 ) ) ;
    buf_clk cell_6544 ( .C ( clk ), .D ( signal_12135 ), .Q ( signal_12136 ) ) ;
    buf_clk cell_6554 ( .C ( clk ), .D ( signal_12145 ), .Q ( signal_12146 ) ) ;
    buf_clk cell_6564 ( .C ( clk ), .D ( signal_12155 ), .Q ( signal_12156 ) ) ;
    buf_clk cell_6574 ( .C ( clk ), .D ( signal_12165 ), .Q ( signal_12166 ) ) ;
    buf_clk cell_6612 ( .C ( clk ), .D ( signal_12203 ), .Q ( signal_12204 ) ) ;
    buf_clk cell_6622 ( .C ( clk ), .D ( signal_12213 ), .Q ( signal_12214 ) ) ;
    buf_clk cell_6632 ( .C ( clk ), .D ( signal_12223 ), .Q ( signal_12224 ) ) ;
    buf_clk cell_6660 ( .C ( clk ), .D ( signal_12251 ), .Q ( signal_12252 ) ) ;
    buf_clk cell_6670 ( .C ( clk ), .D ( signal_12261 ), .Q ( signal_12262 ) ) ;
    buf_clk cell_6680 ( .C ( clk ), .D ( signal_12271 ), .Q ( signal_12272 ) ) ;
    buf_clk cell_6696 ( .C ( clk ), .D ( signal_12287 ), .Q ( signal_12288 ) ) ;
    buf_clk cell_6712 ( .C ( clk ), .D ( signal_12303 ), .Q ( signal_12304 ) ) ;
    buf_clk cell_6728 ( .C ( clk ), .D ( signal_12319 ), .Q ( signal_12320 ) ) ;
    buf_clk cell_6746 ( .C ( clk ), .D ( signal_12337 ), .Q ( signal_12338 ) ) ;
    buf_clk cell_6764 ( .C ( clk ), .D ( signal_12355 ), .Q ( signal_12356 ) ) ;
    buf_clk cell_6782 ( .C ( clk ), .D ( signal_12373 ), .Q ( signal_12374 ) ) ;
    buf_clk cell_6802 ( .C ( clk ), .D ( signal_12393 ), .Q ( signal_12394 ) ) ;
    buf_clk cell_6810 ( .C ( clk ), .D ( signal_12401 ), .Q ( signal_12402 ) ) ;
    buf_clk cell_6818 ( .C ( clk ), .D ( signal_12409 ), .Q ( signal_12410 ) ) ;
    buf_clk cell_6896 ( .C ( clk ), .D ( signal_12487 ), .Q ( signal_12488 ) ) ;
    buf_clk cell_6916 ( .C ( clk ), .D ( signal_12507 ), .Q ( signal_12508 ) ) ;
    buf_clk cell_6936 ( .C ( clk ), .D ( signal_12527 ), .Q ( signal_12528 ) ) ;
    buf_clk cell_6970 ( .C ( clk ), .D ( signal_12561 ), .Q ( signal_12562 ) ) ;
    buf_clk cell_6982 ( .C ( clk ), .D ( signal_12573 ), .Q ( signal_12574 ) ) ;
    buf_clk cell_6994 ( .C ( clk ), .D ( signal_12585 ), .Q ( signal_12586 ) ) ;
    buf_clk cell_7006 ( .C ( clk ), .D ( signal_12597 ), .Q ( signal_12598 ) ) ;
    buf_clk cell_7020 ( .C ( clk ), .D ( signal_12611 ), .Q ( signal_12612 ) ) ;
    buf_clk cell_7034 ( .C ( clk ), .D ( signal_12625 ), .Q ( signal_12626 ) ) ;

    /* cells in depth 19 */
    buf_clk cell_6165 ( .C ( clk ), .D ( signal_11756 ), .Q ( signal_11757 ) ) ;
    buf_clk cell_6173 ( .C ( clk ), .D ( signal_11764 ), .Q ( signal_11765 ) ) ;
    buf_clk cell_6181 ( .C ( clk ), .D ( signal_11772 ), .Q ( signal_11773 ) ) ;
    buf_clk cell_6193 ( .C ( clk ), .D ( signal_11784 ), .Q ( signal_11785 ) ) ;
    buf_clk cell_6205 ( .C ( clk ), .D ( signal_11796 ), .Q ( signal_11797 ) ) ;
    buf_clk cell_6217 ( .C ( clk ), .D ( signal_11808 ), .Q ( signal_11809 ) ) ;
    buf_clk cell_6223 ( .C ( clk ), .D ( signal_11814 ), .Q ( signal_11815 ) ) ;
    buf_clk cell_6229 ( .C ( clk ), .D ( signal_11820 ), .Q ( signal_11821 ) ) ;
    buf_clk cell_6235 ( .C ( clk ), .D ( signal_11826 ), .Q ( signal_11827 ) ) ;
    buf_clk cell_6241 ( .C ( clk ), .D ( signal_11832 ), .Q ( signal_11833 ) ) ;
    buf_clk cell_6247 ( .C ( clk ), .D ( signal_11838 ), .Q ( signal_11839 ) ) ;
    buf_clk cell_6253 ( .C ( clk ), .D ( signal_11844 ), .Q ( signal_11845 ) ) ;
    buf_clk cell_6267 ( .C ( clk ), .D ( signal_11858 ), .Q ( signal_11859 ) ) ;
    buf_clk cell_6281 ( .C ( clk ), .D ( signal_11872 ), .Q ( signal_11873 ) ) ;
    buf_clk cell_6295 ( .C ( clk ), .D ( signal_11886 ), .Q ( signal_11887 ) ) ;
    buf_clk cell_6303 ( .C ( clk ), .D ( signal_11894 ), .Q ( signal_11895 ) ) ;
    buf_clk cell_6311 ( .C ( clk ), .D ( signal_11902 ), .Q ( signal_11903 ) ) ;
    buf_clk cell_6319 ( .C ( clk ), .D ( signal_11910 ), .Q ( signal_11911 ) ) ;
    buf_clk cell_6333 ( .C ( clk ), .D ( signal_11924 ), .Q ( signal_11925 ) ) ;
    buf_clk cell_6347 ( .C ( clk ), .D ( signal_11938 ), .Q ( signal_11939 ) ) ;
    buf_clk cell_6361 ( .C ( clk ), .D ( signal_11952 ), .Q ( signal_11953 ) ) ;
    buf_clk cell_6369 ( .C ( clk ), .D ( signal_11960 ), .Q ( signal_11961 ) ) ;
    buf_clk cell_6377 ( .C ( clk ), .D ( signal_11968 ), .Q ( signal_11969 ) ) ;
    buf_clk cell_6385 ( .C ( clk ), .D ( signal_11976 ), .Q ( signal_11977 ) ) ;
    buf_clk cell_6387 ( .C ( clk ), .D ( signal_2335 ), .Q ( signal_11979 ) ) ;
    buf_clk cell_6391 ( .C ( clk ), .D ( signal_5194 ), .Q ( signal_11983 ) ) ;
    buf_clk cell_6395 ( .C ( clk ), .D ( signal_5195 ), .Q ( signal_11987 ) ) ;
    buf_clk cell_6405 ( .C ( clk ), .D ( signal_11996 ), .Q ( signal_11997 ) ) ;
    buf_clk cell_6415 ( .C ( clk ), .D ( signal_12006 ), .Q ( signal_12007 ) ) ;
    buf_clk cell_6425 ( .C ( clk ), .D ( signal_12016 ), .Q ( signal_12017 ) ) ;
    buf_clk cell_6453 ( .C ( clk ), .D ( signal_12044 ), .Q ( signal_12045 ) ) ;
    buf_clk cell_6469 ( .C ( clk ), .D ( signal_12060 ), .Q ( signal_12061 ) ) ;
    buf_clk cell_6485 ( .C ( clk ), .D ( signal_12076 ), .Q ( signal_12077 ) ) ;
    buf_clk cell_6489 ( .C ( clk ), .D ( signal_2308 ), .Q ( signal_12081 ) ) ;
    buf_clk cell_6493 ( .C ( clk ), .D ( signal_5140 ), .Q ( signal_12085 ) ) ;
    buf_clk cell_6497 ( .C ( clk ), .D ( signal_5141 ), .Q ( signal_12089 ) ) ;
    buf_clk cell_6513 ( .C ( clk ), .D ( signal_12104 ), .Q ( signal_12105 ) ) ;
    buf_clk cell_6529 ( .C ( clk ), .D ( signal_12120 ), .Q ( signal_12121 ) ) ;
    buf_clk cell_6545 ( .C ( clk ), .D ( signal_12136 ), .Q ( signal_12137 ) ) ;
    buf_clk cell_6555 ( .C ( clk ), .D ( signal_12146 ), .Q ( signal_12147 ) ) ;
    buf_clk cell_6565 ( .C ( clk ), .D ( signal_12156 ), .Q ( signal_12157 ) ) ;
    buf_clk cell_6575 ( .C ( clk ), .D ( signal_12166 ), .Q ( signal_12167 ) ) ;
    buf_clk cell_6579 ( .C ( clk ), .D ( signal_2318 ), .Q ( signal_12171 ) ) ;
    buf_clk cell_6583 ( .C ( clk ), .D ( signal_5160 ), .Q ( signal_12175 ) ) ;
    buf_clk cell_6587 ( .C ( clk ), .D ( signal_5161 ), .Q ( signal_12179 ) ) ;
    buf_clk cell_6591 ( .C ( clk ), .D ( signal_2336 ), .Q ( signal_12183 ) ) ;
    buf_clk cell_6597 ( .C ( clk ), .D ( signal_5196 ), .Q ( signal_12189 ) ) ;
    buf_clk cell_6603 ( .C ( clk ), .D ( signal_5197 ), .Q ( signal_12195 ) ) ;
    buf_clk cell_6613 ( .C ( clk ), .D ( signal_12204 ), .Q ( signal_12205 ) ) ;
    buf_clk cell_6623 ( .C ( clk ), .D ( signal_12214 ), .Q ( signal_12215 ) ) ;
    buf_clk cell_6633 ( .C ( clk ), .D ( signal_12224 ), .Q ( signal_12225 ) ) ;
    buf_clk cell_6639 ( .C ( clk ), .D ( signal_2343 ), .Q ( signal_12231 ) ) ;
    buf_clk cell_6645 ( .C ( clk ), .D ( signal_5210 ), .Q ( signal_12237 ) ) ;
    buf_clk cell_6651 ( .C ( clk ), .D ( signal_5211 ), .Q ( signal_12243 ) ) ;
    buf_clk cell_6661 ( .C ( clk ), .D ( signal_12252 ), .Q ( signal_12253 ) ) ;
    buf_clk cell_6671 ( .C ( clk ), .D ( signal_12262 ), .Q ( signal_12263 ) ) ;
    buf_clk cell_6681 ( .C ( clk ), .D ( signal_12272 ), .Q ( signal_12273 ) ) ;
    buf_clk cell_6697 ( .C ( clk ), .D ( signal_12288 ), .Q ( signal_12289 ) ) ;
    buf_clk cell_6713 ( .C ( clk ), .D ( signal_12304 ), .Q ( signal_12305 ) ) ;
    buf_clk cell_6729 ( .C ( clk ), .D ( signal_12320 ), .Q ( signal_12321 ) ) ;
    buf_clk cell_6747 ( .C ( clk ), .D ( signal_12338 ), .Q ( signal_12339 ) ) ;
    buf_clk cell_6765 ( .C ( clk ), .D ( signal_12356 ), .Q ( signal_12357 ) ) ;
    buf_clk cell_6783 ( .C ( clk ), .D ( signal_12374 ), .Q ( signal_12375 ) ) ;
    buf_clk cell_6803 ( .C ( clk ), .D ( signal_12394 ), .Q ( signal_12395 ) ) ;
    buf_clk cell_6811 ( .C ( clk ), .D ( signal_12402 ), .Q ( signal_12403 ) ) ;
    buf_clk cell_6819 ( .C ( clk ), .D ( signal_12410 ), .Q ( signal_12411 ) ) ;
    buf_clk cell_6825 ( .C ( clk ), .D ( signal_2306 ), .Q ( signal_12417 ) ) ;
    buf_clk cell_6833 ( .C ( clk ), .D ( signal_5136 ), .Q ( signal_12425 ) ) ;
    buf_clk cell_6841 ( .C ( clk ), .D ( signal_5137 ), .Q ( signal_12433 ) ) ;
    buf_clk cell_6897 ( .C ( clk ), .D ( signal_12488 ), .Q ( signal_12489 ) ) ;
    buf_clk cell_6917 ( .C ( clk ), .D ( signal_12508 ), .Q ( signal_12509 ) ) ;
    buf_clk cell_6937 ( .C ( clk ), .D ( signal_12528 ), .Q ( signal_12529 ) ) ;
    buf_clk cell_6971 ( .C ( clk ), .D ( signal_12562 ), .Q ( signal_12563 ) ) ;
    buf_clk cell_6983 ( .C ( clk ), .D ( signal_12574 ), .Q ( signal_12575 ) ) ;
    buf_clk cell_6995 ( .C ( clk ), .D ( signal_12586 ), .Q ( signal_12587 ) ) ;
    buf_clk cell_7007 ( .C ( clk ), .D ( signal_12598 ), .Q ( signal_12599 ) ) ;
    buf_clk cell_7021 ( .C ( clk ), .D ( signal_12612 ), .Q ( signal_12613 ) ) ;
    buf_clk cell_7035 ( .C ( clk ), .D ( signal_12626 ), .Q ( signal_12627 ) ) ;
    buf_clk cell_7047 ( .C ( clk ), .D ( signal_2328 ), .Q ( signal_12639 ) ) ;
    buf_clk cell_7061 ( .C ( clk ), .D ( signal_5180 ), .Q ( signal_12653 ) ) ;
    buf_clk cell_7075 ( .C ( clk ), .D ( signal_5181 ), .Q ( signal_12667 ) ) ;

    /* cells in depth 20 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2269 ( .a ({signal_11468, signal_11462, signal_11456}), .b ({signal_5015, signal_5014, signal_2245}), .clk ( clk ), .r ({Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({signal_5093, signal_5092, signal_2284}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2270 ( .a ({signal_11492, signal_11484, signal_11476}), .b ({signal_5019, signal_5018, signal_2247}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481]}), .c ({signal_5095, signal_5094, signal_2285}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2296 ( .a ({signal_11510, signal_11504, signal_11498}), .b ({signal_5089, signal_5088, signal_2282}), .clk ( clk ), .r ({Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({signal_5147, signal_5146, signal_2311}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2316 ( .a ({signal_11540, signal_11530, signal_11520}), .b ({signal_5139, signal_5138, signal_2307}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487]}), .c ({signal_5187, signal_5186, signal_2331}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2317 ( .a ({signal_11558, signal_11552, signal_11546}), .b ({signal_5117, signal_5116, signal_2296}), .clk ( clk ), .r ({Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_5189, signal_5188, signal_2332}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2318 ( .a ({signal_11570, signal_11566, signal_11562}), .b ({signal_5017, signal_5016, signal_2246}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493]}), .c ({signal_5191, signal_5190, signal_2333}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2325 ( .a ({signal_11594, signal_11586, signal_11578}), .b ({signal_5151, signal_5150, signal_2313}), .clk ( clk ), .r ({Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({signal_5205, signal_5204, signal_2340}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2327 ( .a ({signal_11612, signal_11606, signal_11600}), .b ({signal_5155, signal_5154, signal_2315}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499]}), .c ({signal_5209, signal_5208, signal_2342}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2331 ( .a ({signal_11636, signal_11628, signal_11620}), .b ({signal_5179, signal_5178, signal_2327}), .clk ( clk ), .r ({Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({signal_5217, signal_5216, signal_2346}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2332 ( .a ({signal_11654, signal_11648, signal_11642}), .b ({signal_5159, signal_5158, signal_2317}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505]}), .c ({signal_5219, signal_5218, signal_2347}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2333 ( .a ({signal_11678, signal_11670, signal_11662}), .b ({signal_5183, signal_5182, signal_2329}), .clk ( clk ), .r ({Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({signal_5221, signal_5220, signal_2348}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2335 ( .a ({signal_5205, signal_5204, signal_2340}), .b ({signal_5225, signal_5224, signal_2350}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2336 ( .a ({signal_5219, signal_5218, signal_2347}), .b ({signal_5227, signal_5226, signal_2351}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2337 ( .a ({signal_11690, signal_11686, signal_11682}), .b ({signal_5207, signal_5206, signal_2341}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511]}), .c ({signal_5229, signal_5228, signal_2352}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2339 ( .a ({signal_11708, signal_11702, signal_11696}), .b ({signal_5213, signal_5212, signal_2344}), .clk ( clk ), .r ({Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({signal_5233, signal_5232, signal_2354}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2340 ( .a ({signal_11726, signal_11720, signal_11714}), .b ({signal_5199, signal_5198, signal_2337}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517]}), .c ({signal_5235, signal_5234, signal_2355}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2341 ( .a ({signal_11738, signal_11734, signal_11730}), .b ({signal_5201, signal_5200, signal_2338}), .clk ( clk ), .r ({Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_5237, signal_5236, signal_2356}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2342 ( .a ({signal_11750, signal_11746, signal_11742}), .b ({signal_5215, signal_5214, signal_2345}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523]}), .c ({signal_5239, signal_5238, signal_2357}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2343 ( .a ({signal_5203, signal_5202, signal_2339}), .b ({signal_5185, signal_5184, signal_2330}), .clk ( clk ), .r ({Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({signal_5241, signal_5240, signal_2358}) ) ;
    buf_clk cell_6166 ( .C ( clk ), .D ( signal_11757 ), .Q ( signal_11758 ) ) ;
    buf_clk cell_6174 ( .C ( clk ), .D ( signal_11765 ), .Q ( signal_11766 ) ) ;
    buf_clk cell_6182 ( .C ( clk ), .D ( signal_11773 ), .Q ( signal_11774 ) ) ;
    buf_clk cell_6194 ( .C ( clk ), .D ( signal_11785 ), .Q ( signal_11786 ) ) ;
    buf_clk cell_6206 ( .C ( clk ), .D ( signal_11797 ), .Q ( signal_11798 ) ) ;
    buf_clk cell_6218 ( .C ( clk ), .D ( signal_11809 ), .Q ( signal_11810 ) ) ;
    buf_clk cell_6224 ( .C ( clk ), .D ( signal_11815 ), .Q ( signal_11816 ) ) ;
    buf_clk cell_6230 ( .C ( clk ), .D ( signal_11821 ), .Q ( signal_11822 ) ) ;
    buf_clk cell_6236 ( .C ( clk ), .D ( signal_11827 ), .Q ( signal_11828 ) ) ;
    buf_clk cell_6242 ( .C ( clk ), .D ( signal_11833 ), .Q ( signal_11834 ) ) ;
    buf_clk cell_6248 ( .C ( clk ), .D ( signal_11839 ), .Q ( signal_11840 ) ) ;
    buf_clk cell_6254 ( .C ( clk ), .D ( signal_11845 ), .Q ( signal_11846 ) ) ;
    buf_clk cell_6268 ( .C ( clk ), .D ( signal_11859 ), .Q ( signal_11860 ) ) ;
    buf_clk cell_6282 ( .C ( clk ), .D ( signal_11873 ), .Q ( signal_11874 ) ) ;
    buf_clk cell_6296 ( .C ( clk ), .D ( signal_11887 ), .Q ( signal_11888 ) ) ;
    buf_clk cell_6304 ( .C ( clk ), .D ( signal_11895 ), .Q ( signal_11896 ) ) ;
    buf_clk cell_6312 ( .C ( clk ), .D ( signal_11903 ), .Q ( signal_11904 ) ) ;
    buf_clk cell_6320 ( .C ( clk ), .D ( signal_11911 ), .Q ( signal_11912 ) ) ;
    buf_clk cell_6334 ( .C ( clk ), .D ( signal_11925 ), .Q ( signal_11926 ) ) ;
    buf_clk cell_6348 ( .C ( clk ), .D ( signal_11939 ), .Q ( signal_11940 ) ) ;
    buf_clk cell_6362 ( .C ( clk ), .D ( signal_11953 ), .Q ( signal_11954 ) ) ;
    buf_clk cell_6370 ( .C ( clk ), .D ( signal_11961 ), .Q ( signal_11962 ) ) ;
    buf_clk cell_6378 ( .C ( clk ), .D ( signal_11969 ), .Q ( signal_11970 ) ) ;
    buf_clk cell_6386 ( .C ( clk ), .D ( signal_11977 ), .Q ( signal_11978 ) ) ;
    buf_clk cell_6388 ( .C ( clk ), .D ( signal_11979 ), .Q ( signal_11980 ) ) ;
    buf_clk cell_6392 ( .C ( clk ), .D ( signal_11983 ), .Q ( signal_11984 ) ) ;
    buf_clk cell_6396 ( .C ( clk ), .D ( signal_11987 ), .Q ( signal_11988 ) ) ;
    buf_clk cell_6406 ( .C ( clk ), .D ( signal_11997 ), .Q ( signal_11998 ) ) ;
    buf_clk cell_6416 ( .C ( clk ), .D ( signal_12007 ), .Q ( signal_12008 ) ) ;
    buf_clk cell_6426 ( .C ( clk ), .D ( signal_12017 ), .Q ( signal_12018 ) ) ;
    buf_clk cell_6454 ( .C ( clk ), .D ( signal_12045 ), .Q ( signal_12046 ) ) ;
    buf_clk cell_6470 ( .C ( clk ), .D ( signal_12061 ), .Q ( signal_12062 ) ) ;
    buf_clk cell_6486 ( .C ( clk ), .D ( signal_12077 ), .Q ( signal_12078 ) ) ;
    buf_clk cell_6490 ( .C ( clk ), .D ( signal_12081 ), .Q ( signal_12082 ) ) ;
    buf_clk cell_6494 ( .C ( clk ), .D ( signal_12085 ), .Q ( signal_12086 ) ) ;
    buf_clk cell_6498 ( .C ( clk ), .D ( signal_12089 ), .Q ( signal_12090 ) ) ;
    buf_clk cell_6514 ( .C ( clk ), .D ( signal_12105 ), .Q ( signal_12106 ) ) ;
    buf_clk cell_6530 ( .C ( clk ), .D ( signal_12121 ), .Q ( signal_12122 ) ) ;
    buf_clk cell_6546 ( .C ( clk ), .D ( signal_12137 ), .Q ( signal_12138 ) ) ;
    buf_clk cell_6556 ( .C ( clk ), .D ( signal_12147 ), .Q ( signal_12148 ) ) ;
    buf_clk cell_6566 ( .C ( clk ), .D ( signal_12157 ), .Q ( signal_12158 ) ) ;
    buf_clk cell_6576 ( .C ( clk ), .D ( signal_12167 ), .Q ( signal_12168 ) ) ;
    buf_clk cell_6580 ( .C ( clk ), .D ( signal_12171 ), .Q ( signal_12172 ) ) ;
    buf_clk cell_6584 ( .C ( clk ), .D ( signal_12175 ), .Q ( signal_12176 ) ) ;
    buf_clk cell_6588 ( .C ( clk ), .D ( signal_12179 ), .Q ( signal_12180 ) ) ;
    buf_clk cell_6592 ( .C ( clk ), .D ( signal_12183 ), .Q ( signal_12184 ) ) ;
    buf_clk cell_6598 ( .C ( clk ), .D ( signal_12189 ), .Q ( signal_12190 ) ) ;
    buf_clk cell_6604 ( .C ( clk ), .D ( signal_12195 ), .Q ( signal_12196 ) ) ;
    buf_clk cell_6614 ( .C ( clk ), .D ( signal_12205 ), .Q ( signal_12206 ) ) ;
    buf_clk cell_6624 ( .C ( clk ), .D ( signal_12215 ), .Q ( signal_12216 ) ) ;
    buf_clk cell_6634 ( .C ( clk ), .D ( signal_12225 ), .Q ( signal_12226 ) ) ;
    buf_clk cell_6640 ( .C ( clk ), .D ( signal_12231 ), .Q ( signal_12232 ) ) ;
    buf_clk cell_6646 ( .C ( clk ), .D ( signal_12237 ), .Q ( signal_12238 ) ) ;
    buf_clk cell_6652 ( .C ( clk ), .D ( signal_12243 ), .Q ( signal_12244 ) ) ;
    buf_clk cell_6662 ( .C ( clk ), .D ( signal_12253 ), .Q ( signal_12254 ) ) ;
    buf_clk cell_6672 ( .C ( clk ), .D ( signal_12263 ), .Q ( signal_12264 ) ) ;
    buf_clk cell_6682 ( .C ( clk ), .D ( signal_12273 ), .Q ( signal_12274 ) ) ;
    buf_clk cell_6698 ( .C ( clk ), .D ( signal_12289 ), .Q ( signal_12290 ) ) ;
    buf_clk cell_6714 ( .C ( clk ), .D ( signal_12305 ), .Q ( signal_12306 ) ) ;
    buf_clk cell_6730 ( .C ( clk ), .D ( signal_12321 ), .Q ( signal_12322 ) ) ;
    buf_clk cell_6748 ( .C ( clk ), .D ( signal_12339 ), .Q ( signal_12340 ) ) ;
    buf_clk cell_6766 ( .C ( clk ), .D ( signal_12357 ), .Q ( signal_12358 ) ) ;
    buf_clk cell_6784 ( .C ( clk ), .D ( signal_12375 ), .Q ( signal_12376 ) ) ;
    buf_clk cell_6804 ( .C ( clk ), .D ( signal_12395 ), .Q ( signal_12396 ) ) ;
    buf_clk cell_6812 ( .C ( clk ), .D ( signal_12403 ), .Q ( signal_12404 ) ) ;
    buf_clk cell_6820 ( .C ( clk ), .D ( signal_12411 ), .Q ( signal_12412 ) ) ;
    buf_clk cell_6826 ( .C ( clk ), .D ( signal_12417 ), .Q ( signal_12418 ) ) ;
    buf_clk cell_6834 ( .C ( clk ), .D ( signal_12425 ), .Q ( signal_12426 ) ) ;
    buf_clk cell_6842 ( .C ( clk ), .D ( signal_12433 ), .Q ( signal_12434 ) ) ;
    buf_clk cell_6898 ( .C ( clk ), .D ( signal_12489 ), .Q ( signal_12490 ) ) ;
    buf_clk cell_6918 ( .C ( clk ), .D ( signal_12509 ), .Q ( signal_12510 ) ) ;
    buf_clk cell_6938 ( .C ( clk ), .D ( signal_12529 ), .Q ( signal_12530 ) ) ;
    buf_clk cell_6972 ( .C ( clk ), .D ( signal_12563 ), .Q ( signal_12564 ) ) ;
    buf_clk cell_6984 ( .C ( clk ), .D ( signal_12575 ), .Q ( signal_12576 ) ) ;
    buf_clk cell_6996 ( .C ( clk ), .D ( signal_12587 ), .Q ( signal_12588 ) ) ;
    buf_clk cell_7008 ( .C ( clk ), .D ( signal_12599 ), .Q ( signal_12600 ) ) ;
    buf_clk cell_7022 ( .C ( clk ), .D ( signal_12613 ), .Q ( signal_12614 ) ) ;
    buf_clk cell_7036 ( .C ( clk ), .D ( signal_12627 ), .Q ( signal_12628 ) ) ;
    buf_clk cell_7048 ( .C ( clk ), .D ( signal_12639 ), .Q ( signal_12640 ) ) ;
    buf_clk cell_7062 ( .C ( clk ), .D ( signal_12653 ), .Q ( signal_12654 ) ) ;
    buf_clk cell_7076 ( .C ( clk ), .D ( signal_12667 ), .Q ( signal_12668 ) ) ;

    /* cells in depth 21 */
    buf_clk cell_6389 ( .C ( clk ), .D ( signal_11980 ), .Q ( signal_11981 ) ) ;
    buf_clk cell_6393 ( .C ( clk ), .D ( signal_11984 ), .Q ( signal_11985 ) ) ;
    buf_clk cell_6397 ( .C ( clk ), .D ( signal_11988 ), .Q ( signal_11989 ) ) ;
    buf_clk cell_6407 ( .C ( clk ), .D ( signal_11998 ), .Q ( signal_11999 ) ) ;
    buf_clk cell_6417 ( .C ( clk ), .D ( signal_12008 ), .Q ( signal_12009 ) ) ;
    buf_clk cell_6427 ( .C ( clk ), .D ( signal_12018 ), .Q ( signal_12019 ) ) ;
    buf_clk cell_6429 ( .C ( clk ), .D ( signal_2354 ), .Q ( signal_12021 ) ) ;
    buf_clk cell_6431 ( .C ( clk ), .D ( signal_5232 ), .Q ( signal_12023 ) ) ;
    buf_clk cell_6433 ( .C ( clk ), .D ( signal_5233 ), .Q ( signal_12025 ) ) ;
    buf_clk cell_6435 ( .C ( clk ), .D ( signal_2357 ), .Q ( signal_12027 ) ) ;
    buf_clk cell_6437 ( .C ( clk ), .D ( signal_5238 ), .Q ( signal_12029 ) ) ;
    buf_clk cell_6439 ( .C ( clk ), .D ( signal_5239 ), .Q ( signal_12031 ) ) ;
    buf_clk cell_6455 ( .C ( clk ), .D ( signal_12046 ), .Q ( signal_12047 ) ) ;
    buf_clk cell_6471 ( .C ( clk ), .D ( signal_12062 ), .Q ( signal_12063 ) ) ;
    buf_clk cell_6487 ( .C ( clk ), .D ( signal_12078 ), .Q ( signal_12079 ) ) ;
    buf_clk cell_6491 ( .C ( clk ), .D ( signal_12082 ), .Q ( signal_12083 ) ) ;
    buf_clk cell_6495 ( .C ( clk ), .D ( signal_12086 ), .Q ( signal_12087 ) ) ;
    buf_clk cell_6499 ( .C ( clk ), .D ( signal_12090 ), .Q ( signal_12091 ) ) ;
    buf_clk cell_6515 ( .C ( clk ), .D ( signal_12106 ), .Q ( signal_12107 ) ) ;
    buf_clk cell_6531 ( .C ( clk ), .D ( signal_12122 ), .Q ( signal_12123 ) ) ;
    buf_clk cell_6547 ( .C ( clk ), .D ( signal_12138 ), .Q ( signal_12139 ) ) ;
    buf_clk cell_6557 ( .C ( clk ), .D ( signal_12148 ), .Q ( signal_12149 ) ) ;
    buf_clk cell_6567 ( .C ( clk ), .D ( signal_12158 ), .Q ( signal_12159 ) ) ;
    buf_clk cell_6577 ( .C ( clk ), .D ( signal_12168 ), .Q ( signal_12169 ) ) ;
    buf_clk cell_6581 ( .C ( clk ), .D ( signal_12172 ), .Q ( signal_12173 ) ) ;
    buf_clk cell_6585 ( .C ( clk ), .D ( signal_12176 ), .Q ( signal_12177 ) ) ;
    buf_clk cell_6589 ( .C ( clk ), .D ( signal_12180 ), .Q ( signal_12181 ) ) ;
    buf_clk cell_6593 ( .C ( clk ), .D ( signal_12184 ), .Q ( signal_12185 ) ) ;
    buf_clk cell_6599 ( .C ( clk ), .D ( signal_12190 ), .Q ( signal_12191 ) ) ;
    buf_clk cell_6605 ( .C ( clk ), .D ( signal_12196 ), .Q ( signal_12197 ) ) ;
    buf_clk cell_6615 ( .C ( clk ), .D ( signal_12206 ), .Q ( signal_12207 ) ) ;
    buf_clk cell_6625 ( .C ( clk ), .D ( signal_12216 ), .Q ( signal_12217 ) ) ;
    buf_clk cell_6635 ( .C ( clk ), .D ( signal_12226 ), .Q ( signal_12227 ) ) ;
    buf_clk cell_6641 ( .C ( clk ), .D ( signal_12232 ), .Q ( signal_12233 ) ) ;
    buf_clk cell_6647 ( .C ( clk ), .D ( signal_12238 ), .Q ( signal_12239 ) ) ;
    buf_clk cell_6653 ( .C ( clk ), .D ( signal_12244 ), .Q ( signal_12245 ) ) ;
    buf_clk cell_6663 ( .C ( clk ), .D ( signal_12254 ), .Q ( signal_12255 ) ) ;
    buf_clk cell_6673 ( .C ( clk ), .D ( signal_12264 ), .Q ( signal_12265 ) ) ;
    buf_clk cell_6683 ( .C ( clk ), .D ( signal_12274 ), .Q ( signal_12275 ) ) ;
    buf_clk cell_6699 ( .C ( clk ), .D ( signal_12290 ), .Q ( signal_12291 ) ) ;
    buf_clk cell_6715 ( .C ( clk ), .D ( signal_12306 ), .Q ( signal_12307 ) ) ;
    buf_clk cell_6731 ( .C ( clk ), .D ( signal_12322 ), .Q ( signal_12323 ) ) ;
    buf_clk cell_6749 ( .C ( clk ), .D ( signal_12340 ), .Q ( signal_12341 ) ) ;
    buf_clk cell_6767 ( .C ( clk ), .D ( signal_12358 ), .Q ( signal_12359 ) ) ;
    buf_clk cell_6785 ( .C ( clk ), .D ( signal_12376 ), .Q ( signal_12377 ) ) ;
    buf_clk cell_6789 ( .C ( clk ), .D ( signal_2348 ), .Q ( signal_12381 ) ) ;
    buf_clk cell_6793 ( .C ( clk ), .D ( signal_5220 ), .Q ( signal_12385 ) ) ;
    buf_clk cell_6797 ( .C ( clk ), .D ( signal_5221 ), .Q ( signal_12389 ) ) ;
    buf_clk cell_6805 ( .C ( clk ), .D ( signal_12396 ), .Q ( signal_12397 ) ) ;
    buf_clk cell_6813 ( .C ( clk ), .D ( signal_12404 ), .Q ( signal_12405 ) ) ;
    buf_clk cell_6821 ( .C ( clk ), .D ( signal_12412 ), .Q ( signal_12413 ) ) ;
    buf_clk cell_6827 ( .C ( clk ), .D ( signal_12418 ), .Q ( signal_12419 ) ) ;
    buf_clk cell_6835 ( .C ( clk ), .D ( signal_12426 ), .Q ( signal_12427 ) ) ;
    buf_clk cell_6843 ( .C ( clk ), .D ( signal_12434 ), .Q ( signal_12435 ) ) ;
    buf_clk cell_6849 ( .C ( clk ), .D ( signal_2285 ), .Q ( signal_12441 ) ) ;
    buf_clk cell_6855 ( .C ( clk ), .D ( signal_5094 ), .Q ( signal_12447 ) ) ;
    buf_clk cell_6861 ( .C ( clk ), .D ( signal_5095 ), .Q ( signal_12453 ) ) ;
    buf_clk cell_6899 ( .C ( clk ), .D ( signal_12490 ), .Q ( signal_12491 ) ) ;
    buf_clk cell_6919 ( .C ( clk ), .D ( signal_12510 ), .Q ( signal_12511 ) ) ;
    buf_clk cell_6939 ( .C ( clk ), .D ( signal_12530 ), .Q ( signal_12531 ) ) ;
    buf_clk cell_6945 ( .C ( clk ), .D ( signal_2332 ), .Q ( signal_12537 ) ) ;
    buf_clk cell_6953 ( .C ( clk ), .D ( signal_5188 ), .Q ( signal_12545 ) ) ;
    buf_clk cell_6961 ( .C ( clk ), .D ( signal_5189 ), .Q ( signal_12553 ) ) ;
    buf_clk cell_6973 ( .C ( clk ), .D ( signal_12564 ), .Q ( signal_12565 ) ) ;
    buf_clk cell_6985 ( .C ( clk ), .D ( signal_12576 ), .Q ( signal_12577 ) ) ;
    buf_clk cell_6997 ( .C ( clk ), .D ( signal_12588 ), .Q ( signal_12589 ) ) ;
    buf_clk cell_7009 ( .C ( clk ), .D ( signal_12600 ), .Q ( signal_12601 ) ) ;
    buf_clk cell_7023 ( .C ( clk ), .D ( signal_12614 ), .Q ( signal_12615 ) ) ;
    buf_clk cell_7037 ( .C ( clk ), .D ( signal_12628 ), .Q ( signal_12629 ) ) ;
    buf_clk cell_7049 ( .C ( clk ), .D ( signal_12640 ), .Q ( signal_12641 ) ) ;
    buf_clk cell_7063 ( .C ( clk ), .D ( signal_12654 ), .Q ( signal_12655 ) ) ;
    buf_clk cell_7077 ( .C ( clk ), .D ( signal_12668 ), .Q ( signal_12669 ) ) ;

    /* cells in depth 22 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2319 ( .a ({signal_11774, signal_11766, signal_11758}), .b ({signal_5147, signal_5146, signal_2311}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529]}), .c ({signal_5193, signal_5192, signal_2334}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2334 ( .a ({signal_11810, signal_11798, signal_11786}), .b ({signal_5187, signal_5186, signal_2331}), .clk ( clk ), .r ({Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({signal_5223, signal_5222, signal_2349}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2338 ( .a ({signal_11828, signal_11822, signal_11816}), .b ({signal_5209, signal_5208, signal_2342}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535]}), .c ({signal_5231, signal_5230, signal_2353}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2344 ( .a ({signal_5217, signal_5216, signal_2346}), .b ({signal_5093, signal_5092, signal_2284}), .clk ( clk ), .r ({Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({signal_5243, signal_5242, signal_2359}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2346 ( .a ({signal_11846, signal_11840, signal_11834}), .b ({signal_5225, signal_5224, signal_2350}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541]}), .c ({signal_5247, signal_5246, signal_2361}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2348 ( .a ({signal_11888, signal_11874, signal_11860}), .b ({signal_5235, signal_5234, signal_2355}), .clk ( clk ), .r ({Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({signal_5251, signal_5250, signal_2363}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2349 ( .a ({signal_11912, signal_11904, signal_11896}), .b ({signal_5237, signal_5236, signal_2356}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547]}), .c ({signal_5253, signal_5252, signal_2364}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2350 ( .a ({signal_11954, signal_11940, signal_11926}), .b ({signal_5227, signal_5226, signal_2351}), .clk ( clk ), .r ({Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_5255, signal_5254, signal_2365}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2351 ( .a ({signal_11978, signal_11970, signal_11962}), .b ({signal_5241, signal_5240, signal_2358}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553]}), .c ({signal_5257, signal_5256, signal_2366}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2352 ( .a ({signal_5229, signal_5228, signal_2352}), .b ({signal_5191, signal_5190, signal_2333}), .clk ( clk ), .r ({Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({signal_5259, signal_5258, signal_2367}) ) ;
    buf_clk cell_6390 ( .C ( clk ), .D ( signal_11981 ), .Q ( signal_11982 ) ) ;
    buf_clk cell_6394 ( .C ( clk ), .D ( signal_11985 ), .Q ( signal_11986 ) ) ;
    buf_clk cell_6398 ( .C ( clk ), .D ( signal_11989 ), .Q ( signal_11990 ) ) ;
    buf_clk cell_6408 ( .C ( clk ), .D ( signal_11999 ), .Q ( signal_12000 ) ) ;
    buf_clk cell_6418 ( .C ( clk ), .D ( signal_12009 ), .Q ( signal_12010 ) ) ;
    buf_clk cell_6428 ( .C ( clk ), .D ( signal_12019 ), .Q ( signal_12020 ) ) ;
    buf_clk cell_6430 ( .C ( clk ), .D ( signal_12021 ), .Q ( signal_12022 ) ) ;
    buf_clk cell_6432 ( .C ( clk ), .D ( signal_12023 ), .Q ( signal_12024 ) ) ;
    buf_clk cell_6434 ( .C ( clk ), .D ( signal_12025 ), .Q ( signal_12026 ) ) ;
    buf_clk cell_6436 ( .C ( clk ), .D ( signal_12027 ), .Q ( signal_12028 ) ) ;
    buf_clk cell_6438 ( .C ( clk ), .D ( signal_12029 ), .Q ( signal_12030 ) ) ;
    buf_clk cell_6440 ( .C ( clk ), .D ( signal_12031 ), .Q ( signal_12032 ) ) ;
    buf_clk cell_6456 ( .C ( clk ), .D ( signal_12047 ), .Q ( signal_12048 ) ) ;
    buf_clk cell_6472 ( .C ( clk ), .D ( signal_12063 ), .Q ( signal_12064 ) ) ;
    buf_clk cell_6488 ( .C ( clk ), .D ( signal_12079 ), .Q ( signal_12080 ) ) ;
    buf_clk cell_6492 ( .C ( clk ), .D ( signal_12083 ), .Q ( signal_12084 ) ) ;
    buf_clk cell_6496 ( .C ( clk ), .D ( signal_12087 ), .Q ( signal_12088 ) ) ;
    buf_clk cell_6500 ( .C ( clk ), .D ( signal_12091 ), .Q ( signal_12092 ) ) ;
    buf_clk cell_6516 ( .C ( clk ), .D ( signal_12107 ), .Q ( signal_12108 ) ) ;
    buf_clk cell_6532 ( .C ( clk ), .D ( signal_12123 ), .Q ( signal_12124 ) ) ;
    buf_clk cell_6548 ( .C ( clk ), .D ( signal_12139 ), .Q ( signal_12140 ) ) ;
    buf_clk cell_6558 ( .C ( clk ), .D ( signal_12149 ), .Q ( signal_12150 ) ) ;
    buf_clk cell_6568 ( .C ( clk ), .D ( signal_12159 ), .Q ( signal_12160 ) ) ;
    buf_clk cell_6578 ( .C ( clk ), .D ( signal_12169 ), .Q ( signal_12170 ) ) ;
    buf_clk cell_6582 ( .C ( clk ), .D ( signal_12173 ), .Q ( signal_12174 ) ) ;
    buf_clk cell_6586 ( .C ( clk ), .D ( signal_12177 ), .Q ( signal_12178 ) ) ;
    buf_clk cell_6590 ( .C ( clk ), .D ( signal_12181 ), .Q ( signal_12182 ) ) ;
    buf_clk cell_6594 ( .C ( clk ), .D ( signal_12185 ), .Q ( signal_12186 ) ) ;
    buf_clk cell_6600 ( .C ( clk ), .D ( signal_12191 ), .Q ( signal_12192 ) ) ;
    buf_clk cell_6606 ( .C ( clk ), .D ( signal_12197 ), .Q ( signal_12198 ) ) ;
    buf_clk cell_6616 ( .C ( clk ), .D ( signal_12207 ), .Q ( signal_12208 ) ) ;
    buf_clk cell_6626 ( .C ( clk ), .D ( signal_12217 ), .Q ( signal_12218 ) ) ;
    buf_clk cell_6636 ( .C ( clk ), .D ( signal_12227 ), .Q ( signal_12228 ) ) ;
    buf_clk cell_6642 ( .C ( clk ), .D ( signal_12233 ), .Q ( signal_12234 ) ) ;
    buf_clk cell_6648 ( .C ( clk ), .D ( signal_12239 ), .Q ( signal_12240 ) ) ;
    buf_clk cell_6654 ( .C ( clk ), .D ( signal_12245 ), .Q ( signal_12246 ) ) ;
    buf_clk cell_6664 ( .C ( clk ), .D ( signal_12255 ), .Q ( signal_12256 ) ) ;
    buf_clk cell_6674 ( .C ( clk ), .D ( signal_12265 ), .Q ( signal_12266 ) ) ;
    buf_clk cell_6684 ( .C ( clk ), .D ( signal_12275 ), .Q ( signal_12276 ) ) ;
    buf_clk cell_6700 ( .C ( clk ), .D ( signal_12291 ), .Q ( signal_12292 ) ) ;
    buf_clk cell_6716 ( .C ( clk ), .D ( signal_12307 ), .Q ( signal_12308 ) ) ;
    buf_clk cell_6732 ( .C ( clk ), .D ( signal_12323 ), .Q ( signal_12324 ) ) ;
    buf_clk cell_6750 ( .C ( clk ), .D ( signal_12341 ), .Q ( signal_12342 ) ) ;
    buf_clk cell_6768 ( .C ( clk ), .D ( signal_12359 ), .Q ( signal_12360 ) ) ;
    buf_clk cell_6786 ( .C ( clk ), .D ( signal_12377 ), .Q ( signal_12378 ) ) ;
    buf_clk cell_6790 ( .C ( clk ), .D ( signal_12381 ), .Q ( signal_12382 ) ) ;
    buf_clk cell_6794 ( .C ( clk ), .D ( signal_12385 ), .Q ( signal_12386 ) ) ;
    buf_clk cell_6798 ( .C ( clk ), .D ( signal_12389 ), .Q ( signal_12390 ) ) ;
    buf_clk cell_6806 ( .C ( clk ), .D ( signal_12397 ), .Q ( signal_12398 ) ) ;
    buf_clk cell_6814 ( .C ( clk ), .D ( signal_12405 ), .Q ( signal_12406 ) ) ;
    buf_clk cell_6822 ( .C ( clk ), .D ( signal_12413 ), .Q ( signal_12414 ) ) ;
    buf_clk cell_6828 ( .C ( clk ), .D ( signal_12419 ), .Q ( signal_12420 ) ) ;
    buf_clk cell_6836 ( .C ( clk ), .D ( signal_12427 ), .Q ( signal_12428 ) ) ;
    buf_clk cell_6844 ( .C ( clk ), .D ( signal_12435 ), .Q ( signal_12436 ) ) ;
    buf_clk cell_6850 ( .C ( clk ), .D ( signal_12441 ), .Q ( signal_12442 ) ) ;
    buf_clk cell_6856 ( .C ( clk ), .D ( signal_12447 ), .Q ( signal_12448 ) ) ;
    buf_clk cell_6862 ( .C ( clk ), .D ( signal_12453 ), .Q ( signal_12454 ) ) ;
    buf_clk cell_6900 ( .C ( clk ), .D ( signal_12491 ), .Q ( signal_12492 ) ) ;
    buf_clk cell_6920 ( .C ( clk ), .D ( signal_12511 ), .Q ( signal_12512 ) ) ;
    buf_clk cell_6940 ( .C ( clk ), .D ( signal_12531 ), .Q ( signal_12532 ) ) ;
    buf_clk cell_6946 ( .C ( clk ), .D ( signal_12537 ), .Q ( signal_12538 ) ) ;
    buf_clk cell_6954 ( .C ( clk ), .D ( signal_12545 ), .Q ( signal_12546 ) ) ;
    buf_clk cell_6962 ( .C ( clk ), .D ( signal_12553 ), .Q ( signal_12554 ) ) ;
    buf_clk cell_6974 ( .C ( clk ), .D ( signal_12565 ), .Q ( signal_12566 ) ) ;
    buf_clk cell_6986 ( .C ( clk ), .D ( signal_12577 ), .Q ( signal_12578 ) ) ;
    buf_clk cell_6998 ( .C ( clk ), .D ( signal_12589 ), .Q ( signal_12590 ) ) ;
    buf_clk cell_7010 ( .C ( clk ), .D ( signal_12601 ), .Q ( signal_12602 ) ) ;
    buf_clk cell_7024 ( .C ( clk ), .D ( signal_12615 ), .Q ( signal_12616 ) ) ;
    buf_clk cell_7038 ( .C ( clk ), .D ( signal_12629 ), .Q ( signal_12630 ) ) ;
    buf_clk cell_7050 ( .C ( clk ), .D ( signal_12641 ), .Q ( signal_12642 ) ) ;
    buf_clk cell_7064 ( .C ( clk ), .D ( signal_12655 ), .Q ( signal_12656 ) ) ;
    buf_clk cell_7078 ( .C ( clk ), .D ( signal_12669 ), .Q ( signal_12670 ) ) ;

    /* cells in depth 23 */
    buf_clk cell_6595 ( .C ( clk ), .D ( signal_12186 ), .Q ( signal_12187 ) ) ;
    buf_clk cell_6601 ( .C ( clk ), .D ( signal_12192 ), .Q ( signal_12193 ) ) ;
    buf_clk cell_6607 ( .C ( clk ), .D ( signal_12198 ), .Q ( signal_12199 ) ) ;
    buf_clk cell_6617 ( .C ( clk ), .D ( signal_12208 ), .Q ( signal_12209 ) ) ;
    buf_clk cell_6627 ( .C ( clk ), .D ( signal_12218 ), .Q ( signal_12219 ) ) ;
    buf_clk cell_6637 ( .C ( clk ), .D ( signal_12228 ), .Q ( signal_12229 ) ) ;
    buf_clk cell_6643 ( .C ( clk ), .D ( signal_12234 ), .Q ( signal_12235 ) ) ;
    buf_clk cell_6649 ( .C ( clk ), .D ( signal_12240 ), .Q ( signal_12241 ) ) ;
    buf_clk cell_6655 ( .C ( clk ), .D ( signal_12246 ), .Q ( signal_12247 ) ) ;
    buf_clk cell_6665 ( .C ( clk ), .D ( signal_12256 ), .Q ( signal_12257 ) ) ;
    buf_clk cell_6675 ( .C ( clk ), .D ( signal_12266 ), .Q ( signal_12267 ) ) ;
    buf_clk cell_6685 ( .C ( clk ), .D ( signal_12276 ), .Q ( signal_12277 ) ) ;
    buf_clk cell_6701 ( .C ( clk ), .D ( signal_12292 ), .Q ( signal_12293 ) ) ;
    buf_clk cell_6717 ( .C ( clk ), .D ( signal_12308 ), .Q ( signal_12309 ) ) ;
    buf_clk cell_6733 ( .C ( clk ), .D ( signal_12324 ), .Q ( signal_12325 ) ) ;
    buf_clk cell_6751 ( .C ( clk ), .D ( signal_12342 ), .Q ( signal_12343 ) ) ;
    buf_clk cell_6769 ( .C ( clk ), .D ( signal_12360 ), .Q ( signal_12361 ) ) ;
    buf_clk cell_6787 ( .C ( clk ), .D ( signal_12378 ), .Q ( signal_12379 ) ) ;
    buf_clk cell_6791 ( .C ( clk ), .D ( signal_12382 ), .Q ( signal_12383 ) ) ;
    buf_clk cell_6795 ( .C ( clk ), .D ( signal_12386 ), .Q ( signal_12387 ) ) ;
    buf_clk cell_6799 ( .C ( clk ), .D ( signal_12390 ), .Q ( signal_12391 ) ) ;
    buf_clk cell_6807 ( .C ( clk ), .D ( signal_12398 ), .Q ( signal_12399 ) ) ;
    buf_clk cell_6815 ( .C ( clk ), .D ( signal_12406 ), .Q ( signal_12407 ) ) ;
    buf_clk cell_6823 ( .C ( clk ), .D ( signal_12414 ), .Q ( signal_12415 ) ) ;
    buf_clk cell_6829 ( .C ( clk ), .D ( signal_12420 ), .Q ( signal_12421 ) ) ;
    buf_clk cell_6837 ( .C ( clk ), .D ( signal_12428 ), .Q ( signal_12429 ) ) ;
    buf_clk cell_6845 ( .C ( clk ), .D ( signal_12436 ), .Q ( signal_12437 ) ) ;
    buf_clk cell_6851 ( .C ( clk ), .D ( signal_12442 ), .Q ( signal_12443 ) ) ;
    buf_clk cell_6857 ( .C ( clk ), .D ( signal_12448 ), .Q ( signal_12449 ) ) ;
    buf_clk cell_6863 ( .C ( clk ), .D ( signal_12454 ), .Q ( signal_12455 ) ) ;
    buf_clk cell_6867 ( .C ( clk ), .D ( signal_2361 ), .Q ( signal_12459 ) ) ;
    buf_clk cell_6871 ( .C ( clk ), .D ( signal_5246 ), .Q ( signal_12463 ) ) ;
    buf_clk cell_6875 ( .C ( clk ), .D ( signal_5247 ), .Q ( signal_12467 ) ) ;
    buf_clk cell_6901 ( .C ( clk ), .D ( signal_12492 ), .Q ( signal_12493 ) ) ;
    buf_clk cell_6921 ( .C ( clk ), .D ( signal_12512 ), .Q ( signal_12513 ) ) ;
    buf_clk cell_6941 ( .C ( clk ), .D ( signal_12532 ), .Q ( signal_12533 ) ) ;
    buf_clk cell_6947 ( .C ( clk ), .D ( signal_12538 ), .Q ( signal_12539 ) ) ;
    buf_clk cell_6955 ( .C ( clk ), .D ( signal_12546 ), .Q ( signal_12547 ) ) ;
    buf_clk cell_6963 ( .C ( clk ), .D ( signal_12554 ), .Q ( signal_12555 ) ) ;
    buf_clk cell_6975 ( .C ( clk ), .D ( signal_12566 ), .Q ( signal_12567 ) ) ;
    buf_clk cell_6987 ( .C ( clk ), .D ( signal_12578 ), .Q ( signal_12579 ) ) ;
    buf_clk cell_6999 ( .C ( clk ), .D ( signal_12590 ), .Q ( signal_12591 ) ) ;
    buf_clk cell_7011 ( .C ( clk ), .D ( signal_12602 ), .Q ( signal_12603 ) ) ;
    buf_clk cell_7025 ( .C ( clk ), .D ( signal_12616 ), .Q ( signal_12617 ) ) ;
    buf_clk cell_7039 ( .C ( clk ), .D ( signal_12630 ), .Q ( signal_12631 ) ) ;
    buf_clk cell_7051 ( .C ( clk ), .D ( signal_12642 ), .Q ( signal_12643 ) ) ;
    buf_clk cell_7065 ( .C ( clk ), .D ( signal_12656 ), .Q ( signal_12657 ) ) ;
    buf_clk cell_7079 ( .C ( clk ), .D ( signal_12670 ), .Q ( signal_12671 ) ) ;

    /* cells in depth 24 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2345 ( .a ({signal_11990, signal_11986, signal_11982}), .b ({signal_5193, signal_5192, signal_2334}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559]}), .c ({signal_5245, signal_5244, signal_2360}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2347 ( .a ({signal_12020, signal_12010, signal_12000}), .b ({signal_5231, signal_5230, signal_2353}), .clk ( clk ), .r ({Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({signal_5249, signal_5248, signal_2362}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2353 ( .a ({signal_12026, signal_12024, signal_12022}), .b ({signal_5223, signal_5222, signal_2349}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565]}), .c ({signal_5261, signal_5260, signal_2368}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2354 ( .a ({signal_12032, signal_12030, signal_12028}), .b ({signal_5243, signal_5242, signal_2359}), .clk ( clk ), .r ({Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({signal_5263, signal_5262, signal_2369}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2357 ( .a ({signal_12080, signal_12064, signal_12048}), .b ({signal_5251, signal_5250, signal_2363}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571]}), .c ({signal_5269, signal_5268, signal_2372}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2358 ( .a ({signal_12092, signal_12088, signal_12084}), .b ({signal_5253, signal_5252, signal_2364}), .clk ( clk ), .r ({Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({signal_5271, signal_5270, signal_2373}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2359 ( .a ({signal_12140, signal_12124, signal_12108}), .b ({signal_5255, signal_5254, signal_2365}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577]}), .c ({signal_5273, signal_5272, signal_2374}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2360 ( .a ({signal_12170, signal_12160, signal_12150}), .b ({signal_5257, signal_5256, signal_2366}), .clk ( clk ), .r ({Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_5275, signal_5274, signal_2375}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2361 ( .a ({signal_12182, signal_12178, signal_12174}), .b ({signal_5259, signal_5258, signal_2367}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583]}), .c ({signal_5277, signal_5276, signal_2376}) ) ;
    buf_clk cell_6596 ( .C ( clk ), .D ( signal_12187 ), .Q ( signal_12188 ) ) ;
    buf_clk cell_6602 ( .C ( clk ), .D ( signal_12193 ), .Q ( signal_12194 ) ) ;
    buf_clk cell_6608 ( .C ( clk ), .D ( signal_12199 ), .Q ( signal_12200 ) ) ;
    buf_clk cell_6618 ( .C ( clk ), .D ( signal_12209 ), .Q ( signal_12210 ) ) ;
    buf_clk cell_6628 ( .C ( clk ), .D ( signal_12219 ), .Q ( signal_12220 ) ) ;
    buf_clk cell_6638 ( .C ( clk ), .D ( signal_12229 ), .Q ( signal_12230 ) ) ;
    buf_clk cell_6644 ( .C ( clk ), .D ( signal_12235 ), .Q ( signal_12236 ) ) ;
    buf_clk cell_6650 ( .C ( clk ), .D ( signal_12241 ), .Q ( signal_12242 ) ) ;
    buf_clk cell_6656 ( .C ( clk ), .D ( signal_12247 ), .Q ( signal_12248 ) ) ;
    buf_clk cell_6666 ( .C ( clk ), .D ( signal_12257 ), .Q ( signal_12258 ) ) ;
    buf_clk cell_6676 ( .C ( clk ), .D ( signal_12267 ), .Q ( signal_12268 ) ) ;
    buf_clk cell_6686 ( .C ( clk ), .D ( signal_12277 ), .Q ( signal_12278 ) ) ;
    buf_clk cell_6702 ( .C ( clk ), .D ( signal_12293 ), .Q ( signal_12294 ) ) ;
    buf_clk cell_6718 ( .C ( clk ), .D ( signal_12309 ), .Q ( signal_12310 ) ) ;
    buf_clk cell_6734 ( .C ( clk ), .D ( signal_12325 ), .Q ( signal_12326 ) ) ;
    buf_clk cell_6752 ( .C ( clk ), .D ( signal_12343 ), .Q ( signal_12344 ) ) ;
    buf_clk cell_6770 ( .C ( clk ), .D ( signal_12361 ), .Q ( signal_12362 ) ) ;
    buf_clk cell_6788 ( .C ( clk ), .D ( signal_12379 ), .Q ( signal_12380 ) ) ;
    buf_clk cell_6792 ( .C ( clk ), .D ( signal_12383 ), .Q ( signal_12384 ) ) ;
    buf_clk cell_6796 ( .C ( clk ), .D ( signal_12387 ), .Q ( signal_12388 ) ) ;
    buf_clk cell_6800 ( .C ( clk ), .D ( signal_12391 ), .Q ( signal_12392 ) ) ;
    buf_clk cell_6808 ( .C ( clk ), .D ( signal_12399 ), .Q ( signal_12400 ) ) ;
    buf_clk cell_6816 ( .C ( clk ), .D ( signal_12407 ), .Q ( signal_12408 ) ) ;
    buf_clk cell_6824 ( .C ( clk ), .D ( signal_12415 ), .Q ( signal_12416 ) ) ;
    buf_clk cell_6830 ( .C ( clk ), .D ( signal_12421 ), .Q ( signal_12422 ) ) ;
    buf_clk cell_6838 ( .C ( clk ), .D ( signal_12429 ), .Q ( signal_12430 ) ) ;
    buf_clk cell_6846 ( .C ( clk ), .D ( signal_12437 ), .Q ( signal_12438 ) ) ;
    buf_clk cell_6852 ( .C ( clk ), .D ( signal_12443 ), .Q ( signal_12444 ) ) ;
    buf_clk cell_6858 ( .C ( clk ), .D ( signal_12449 ), .Q ( signal_12450 ) ) ;
    buf_clk cell_6864 ( .C ( clk ), .D ( signal_12455 ), .Q ( signal_12456 ) ) ;
    buf_clk cell_6868 ( .C ( clk ), .D ( signal_12459 ), .Q ( signal_12460 ) ) ;
    buf_clk cell_6872 ( .C ( clk ), .D ( signal_12463 ), .Q ( signal_12464 ) ) ;
    buf_clk cell_6876 ( .C ( clk ), .D ( signal_12467 ), .Q ( signal_12468 ) ) ;
    buf_clk cell_6902 ( .C ( clk ), .D ( signal_12493 ), .Q ( signal_12494 ) ) ;
    buf_clk cell_6922 ( .C ( clk ), .D ( signal_12513 ), .Q ( signal_12514 ) ) ;
    buf_clk cell_6942 ( .C ( clk ), .D ( signal_12533 ), .Q ( signal_12534 ) ) ;
    buf_clk cell_6948 ( .C ( clk ), .D ( signal_12539 ), .Q ( signal_12540 ) ) ;
    buf_clk cell_6956 ( .C ( clk ), .D ( signal_12547 ), .Q ( signal_12548 ) ) ;
    buf_clk cell_6964 ( .C ( clk ), .D ( signal_12555 ), .Q ( signal_12556 ) ) ;
    buf_clk cell_6976 ( .C ( clk ), .D ( signal_12567 ), .Q ( signal_12568 ) ) ;
    buf_clk cell_6988 ( .C ( clk ), .D ( signal_12579 ), .Q ( signal_12580 ) ) ;
    buf_clk cell_7000 ( .C ( clk ), .D ( signal_12591 ), .Q ( signal_12592 ) ) ;
    buf_clk cell_7012 ( .C ( clk ), .D ( signal_12603 ), .Q ( signal_12604 ) ) ;
    buf_clk cell_7026 ( .C ( clk ), .D ( signal_12617 ), .Q ( signal_12618 ) ) ;
    buf_clk cell_7040 ( .C ( clk ), .D ( signal_12631 ), .Q ( signal_12632 ) ) ;
    buf_clk cell_7052 ( .C ( clk ), .D ( signal_12643 ), .Q ( signal_12644 ) ) ;
    buf_clk cell_7066 ( .C ( clk ), .D ( signal_12657 ), .Q ( signal_12658 ) ) ;
    buf_clk cell_7080 ( .C ( clk ), .D ( signal_12671 ), .Q ( signal_12672 ) ) ;

    /* cells in depth 25 */
    buf_clk cell_6831 ( .C ( clk ), .D ( signal_12422 ), .Q ( signal_12423 ) ) ;
    buf_clk cell_6839 ( .C ( clk ), .D ( signal_12430 ), .Q ( signal_12431 ) ) ;
    buf_clk cell_6847 ( .C ( clk ), .D ( signal_12438 ), .Q ( signal_12439 ) ) ;
    buf_clk cell_6853 ( .C ( clk ), .D ( signal_12444 ), .Q ( signal_12445 ) ) ;
    buf_clk cell_6859 ( .C ( clk ), .D ( signal_12450 ), .Q ( signal_12451 ) ) ;
    buf_clk cell_6865 ( .C ( clk ), .D ( signal_12456 ), .Q ( signal_12457 ) ) ;
    buf_clk cell_6869 ( .C ( clk ), .D ( signal_12460 ), .Q ( signal_12461 ) ) ;
    buf_clk cell_6873 ( .C ( clk ), .D ( signal_12464 ), .Q ( signal_12465 ) ) ;
    buf_clk cell_6877 ( .C ( clk ), .D ( signal_12468 ), .Q ( signal_12469 ) ) ;
    buf_clk cell_6879 ( .C ( clk ), .D ( signal_2373 ), .Q ( signal_12471 ) ) ;
    buf_clk cell_6881 ( .C ( clk ), .D ( signal_5270 ), .Q ( signal_12473 ) ) ;
    buf_clk cell_6883 ( .C ( clk ), .D ( signal_5271 ), .Q ( signal_12475 ) ) ;
    buf_clk cell_6903 ( .C ( clk ), .D ( signal_12494 ), .Q ( signal_12495 ) ) ;
    buf_clk cell_6923 ( .C ( clk ), .D ( signal_12514 ), .Q ( signal_12515 ) ) ;
    buf_clk cell_6943 ( .C ( clk ), .D ( signal_12534 ), .Q ( signal_12535 ) ) ;
    buf_clk cell_6949 ( .C ( clk ), .D ( signal_12540 ), .Q ( signal_12541 ) ) ;
    buf_clk cell_6957 ( .C ( clk ), .D ( signal_12548 ), .Q ( signal_12549 ) ) ;
    buf_clk cell_6965 ( .C ( clk ), .D ( signal_12556 ), .Q ( signal_12557 ) ) ;
    buf_clk cell_6977 ( .C ( clk ), .D ( signal_12568 ), .Q ( signal_12569 ) ) ;
    buf_clk cell_6989 ( .C ( clk ), .D ( signal_12580 ), .Q ( signal_12581 ) ) ;
    buf_clk cell_7001 ( .C ( clk ), .D ( signal_12592 ), .Q ( signal_12593 ) ) ;
    buf_clk cell_7013 ( .C ( clk ), .D ( signal_12604 ), .Q ( signal_12605 ) ) ;
    buf_clk cell_7027 ( .C ( clk ), .D ( signal_12618 ), .Q ( signal_12619 ) ) ;
    buf_clk cell_7041 ( .C ( clk ), .D ( signal_12632 ), .Q ( signal_12633 ) ) ;
    buf_clk cell_7053 ( .C ( clk ), .D ( signal_12644 ), .Q ( signal_12645 ) ) ;
    buf_clk cell_7067 ( .C ( clk ), .D ( signal_12658 ), .Q ( signal_12659 ) ) ;
    buf_clk cell_7081 ( .C ( clk ), .D ( signal_12672 ), .Q ( signal_12673 ) ) ;

    /* cells in depth 26 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2355 ( .a ({signal_12200, signal_12194, signal_12188}), .b ({signal_5245, signal_5244, signal_2360}), .clk ( clk ), .r ({Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({signal_5265, signal_5264, signal_2370}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2356 ( .a ({signal_12230, signal_12220, signal_12210}), .b ({signal_5249, signal_5248, signal_2362}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589]}), .c ({signal_5267, signal_5266, signal_2371}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2362 ( .a ({signal_12248, signal_12242, signal_12236}), .b ({signal_5261, signal_5260, signal_2368}), .clk ( clk ), .r ({Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({signal_5279, signal_5278, signal_2377}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2363 ( .a ({signal_12278, signal_12268, signal_12258}), .b ({signal_5263, signal_5262, signal_2369}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595]}), .c ({signal_5281, signal_5280, signal_2378}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2365 ( .a ({signal_5281, signal_5280, signal_2378}), .b ({signal_5285, signal_5284, signal_26}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2368 ( .a ({signal_12326, signal_12310, signal_12294}), .b ({signal_5269, signal_5268, signal_2372}), .clk ( clk ), .r ({Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({signal_5291, signal_5290, signal_2381}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2369 ( .a ({signal_12380, signal_12362, signal_12344}), .b ({signal_5273, signal_5272, signal_2374}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601]}), .c ({signal_5293, signal_5292, signal_2382}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2370 ( .a ({signal_12392, signal_12388, signal_12384}), .b ({signal_5275, signal_5274, signal_2375}), .clk ( clk ), .r ({Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({signal_5295, signal_5294, signal_2383}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2371 ( .a ({signal_12416, signal_12408, signal_12400}), .b ({signal_5277, signal_5276, signal_2376}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607]}), .c ({signal_5297, signal_5296, signal_2384}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2374 ( .a ({signal_5295, signal_5294, signal_2383}), .b ({signal_5303, signal_5302, signal_28}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2375 ( .a ({signal_5297, signal_5296, signal_2384}), .b ({signal_5305, signal_5304, signal_29}) ) ;
    buf_clk cell_6832 ( .C ( clk ), .D ( signal_12423 ), .Q ( signal_12424 ) ) ;
    buf_clk cell_6840 ( .C ( clk ), .D ( signal_12431 ), .Q ( signal_12432 ) ) ;
    buf_clk cell_6848 ( .C ( clk ), .D ( signal_12439 ), .Q ( signal_12440 ) ) ;
    buf_clk cell_6854 ( .C ( clk ), .D ( signal_12445 ), .Q ( signal_12446 ) ) ;
    buf_clk cell_6860 ( .C ( clk ), .D ( signal_12451 ), .Q ( signal_12452 ) ) ;
    buf_clk cell_6866 ( .C ( clk ), .D ( signal_12457 ), .Q ( signal_12458 ) ) ;
    buf_clk cell_6870 ( .C ( clk ), .D ( signal_12461 ), .Q ( signal_12462 ) ) ;
    buf_clk cell_6874 ( .C ( clk ), .D ( signal_12465 ), .Q ( signal_12466 ) ) ;
    buf_clk cell_6878 ( .C ( clk ), .D ( signal_12469 ), .Q ( signal_12470 ) ) ;
    buf_clk cell_6880 ( .C ( clk ), .D ( signal_12471 ), .Q ( signal_12472 ) ) ;
    buf_clk cell_6882 ( .C ( clk ), .D ( signal_12473 ), .Q ( signal_12474 ) ) ;
    buf_clk cell_6884 ( .C ( clk ), .D ( signal_12475 ), .Q ( signal_12476 ) ) ;
    buf_clk cell_6904 ( .C ( clk ), .D ( signal_12495 ), .Q ( signal_12496 ) ) ;
    buf_clk cell_6924 ( .C ( clk ), .D ( signal_12515 ), .Q ( signal_12516 ) ) ;
    buf_clk cell_6944 ( .C ( clk ), .D ( signal_12535 ), .Q ( signal_12536 ) ) ;
    buf_clk cell_6950 ( .C ( clk ), .D ( signal_12541 ), .Q ( signal_12542 ) ) ;
    buf_clk cell_6958 ( .C ( clk ), .D ( signal_12549 ), .Q ( signal_12550 ) ) ;
    buf_clk cell_6966 ( .C ( clk ), .D ( signal_12557 ), .Q ( signal_12558 ) ) ;
    buf_clk cell_6978 ( .C ( clk ), .D ( signal_12569 ), .Q ( signal_12570 ) ) ;
    buf_clk cell_6990 ( .C ( clk ), .D ( signal_12581 ), .Q ( signal_12582 ) ) ;
    buf_clk cell_7002 ( .C ( clk ), .D ( signal_12593 ), .Q ( signal_12594 ) ) ;
    buf_clk cell_7014 ( .C ( clk ), .D ( signal_12605 ), .Q ( signal_12606 ) ) ;
    buf_clk cell_7028 ( .C ( clk ), .D ( signal_12619 ), .Q ( signal_12620 ) ) ;
    buf_clk cell_7042 ( .C ( clk ), .D ( signal_12633 ), .Q ( signal_12634 ) ) ;
    buf_clk cell_7054 ( .C ( clk ), .D ( signal_12645 ), .Q ( signal_12646 ) ) ;
    buf_clk cell_7068 ( .C ( clk ), .D ( signal_12659 ), .Q ( signal_12660 ) ) ;
    buf_clk cell_7082 ( .C ( clk ), .D ( signal_12673 ), .Q ( signal_12674 ) ) ;

    /* cells in depth 27 */
    buf_clk cell_6951 ( .C ( clk ), .D ( signal_12542 ), .Q ( signal_12543 ) ) ;
    buf_clk cell_6959 ( .C ( clk ), .D ( signal_12550 ), .Q ( signal_12551 ) ) ;
    buf_clk cell_6967 ( .C ( clk ), .D ( signal_12558 ), .Q ( signal_12559 ) ) ;
    buf_clk cell_6979 ( .C ( clk ), .D ( signal_12570 ), .Q ( signal_12571 ) ) ;
    buf_clk cell_6991 ( .C ( clk ), .D ( signal_12582 ), .Q ( signal_12583 ) ) ;
    buf_clk cell_7003 ( .C ( clk ), .D ( signal_12594 ), .Q ( signal_12595 ) ) ;
    buf_clk cell_7015 ( .C ( clk ), .D ( signal_12606 ), .Q ( signal_12607 ) ) ;
    buf_clk cell_7029 ( .C ( clk ), .D ( signal_12620 ), .Q ( signal_12621 ) ) ;
    buf_clk cell_7043 ( .C ( clk ), .D ( signal_12634 ), .Q ( signal_12635 ) ) ;
    buf_clk cell_7055 ( .C ( clk ), .D ( signal_12646 ), .Q ( signal_12647 ) ) ;
    buf_clk cell_7069 ( .C ( clk ), .D ( signal_12660 ), .Q ( signal_12661 ) ) ;
    buf_clk cell_7083 ( .C ( clk ), .D ( signal_12674 ), .Q ( signal_12675 ) ) ;
    buf_clk cell_7137 ( .C ( clk ), .D ( signal_26 ), .Q ( signal_12729 ) ) ;
    buf_clk cell_7145 ( .C ( clk ), .D ( signal_5284 ), .Q ( signal_12737 ) ) ;
    buf_clk cell_7153 ( .C ( clk ), .D ( signal_5285 ), .Q ( signal_12745 ) ) ;
    buf_clk cell_7161 ( .C ( clk ), .D ( signal_28 ), .Q ( signal_12753 ) ) ;
    buf_clk cell_7169 ( .C ( clk ), .D ( signal_5302 ), .Q ( signal_12761 ) ) ;
    buf_clk cell_7177 ( .C ( clk ), .D ( signal_5303 ), .Q ( signal_12769 ) ) ;
    buf_clk cell_7185 ( .C ( clk ), .D ( signal_29 ), .Q ( signal_12777 ) ) ;
    buf_clk cell_7193 ( .C ( clk ), .D ( signal_5304 ), .Q ( signal_12785 ) ) ;
    buf_clk cell_7201 ( .C ( clk ), .D ( signal_5305 ), .Q ( signal_12793 ) ) ;

    /* cells in depth 28 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2364 ( .a ({signal_12440, signal_12432, signal_12424}), .b ({signal_5265, signal_5264, signal_2370}), .clk ( clk ), .r ({Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_5283, signal_5282, signal_2379}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2366 ( .a ({signal_5283, signal_5282, signal_2379}), .b ({signal_5287, signal_5286, signal_23}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2367 ( .a ({signal_12458, signal_12452, signal_12446}), .b ({signal_5267, signal_5266, signal_2371}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613]}), .c ({signal_5289, signal_5288, signal_2380}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2372 ( .a ({signal_12470, signal_12466, signal_12462}), .b ({signal_5279, signal_5278, signal_2377}), .clk ( clk ), .r ({Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({signal_5299, signal_5298, signal_2385}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2373 ( .a ({signal_5289, signal_5288, signal_2380}), .b ({signal_5301, signal_5300, signal_30}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2376 ( .a ({signal_5299, signal_5298, signal_2385}), .b ({signal_5307, signal_5306, signal_24}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2377 ( .a ({signal_12476, signal_12474, signal_12472}), .b ({signal_5291, signal_5290, signal_2381}), .clk ( clk ), .r ({Fresh[2621], Fresh[2620], Fresh[2619]}), .c ({signal_5309, signal_5308, signal_2386}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2378 ( .a ({signal_12536, signal_12516, signal_12496}), .b ({signal_5293, signal_5292, signal_2382}), .clk ( clk ), .r ({Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({signal_5311, signal_5310, signal_2387}) ) ;
    buf_clk cell_6952 ( .C ( clk ), .D ( signal_12543 ), .Q ( signal_12544 ) ) ;
    buf_clk cell_6960 ( .C ( clk ), .D ( signal_12551 ), .Q ( signal_12552 ) ) ;
    buf_clk cell_6968 ( .C ( clk ), .D ( signal_12559 ), .Q ( signal_12560 ) ) ;
    buf_clk cell_6980 ( .C ( clk ), .D ( signal_12571 ), .Q ( signal_12572 ) ) ;
    buf_clk cell_6992 ( .C ( clk ), .D ( signal_12583 ), .Q ( signal_12584 ) ) ;
    buf_clk cell_7004 ( .C ( clk ), .D ( signal_12595 ), .Q ( signal_12596 ) ) ;
    buf_clk cell_7016 ( .C ( clk ), .D ( signal_12607 ), .Q ( signal_12608 ) ) ;
    buf_clk cell_7030 ( .C ( clk ), .D ( signal_12621 ), .Q ( signal_12622 ) ) ;
    buf_clk cell_7044 ( .C ( clk ), .D ( signal_12635 ), .Q ( signal_12636 ) ) ;
    buf_clk cell_7056 ( .C ( clk ), .D ( signal_12647 ), .Q ( signal_12648 ) ) ;
    buf_clk cell_7070 ( .C ( clk ), .D ( signal_12661 ), .Q ( signal_12662 ) ) ;
    buf_clk cell_7084 ( .C ( clk ), .D ( signal_12675 ), .Q ( signal_12676 ) ) ;
    buf_clk cell_7138 ( .C ( clk ), .D ( signal_12729 ), .Q ( signal_12730 ) ) ;
    buf_clk cell_7146 ( .C ( clk ), .D ( signal_12737 ), .Q ( signal_12738 ) ) ;
    buf_clk cell_7154 ( .C ( clk ), .D ( signal_12745 ), .Q ( signal_12746 ) ) ;
    buf_clk cell_7162 ( .C ( clk ), .D ( signal_12753 ), .Q ( signal_12754 ) ) ;
    buf_clk cell_7170 ( .C ( clk ), .D ( signal_12761 ), .Q ( signal_12762 ) ) ;
    buf_clk cell_7178 ( .C ( clk ), .D ( signal_12769 ), .Q ( signal_12770 ) ) ;
    buf_clk cell_7186 ( .C ( clk ), .D ( signal_12777 ), .Q ( signal_12778 ) ) ;
    buf_clk cell_7194 ( .C ( clk ), .D ( signal_12785 ), .Q ( signal_12786 ) ) ;
    buf_clk cell_7202 ( .C ( clk ), .D ( signal_12793 ), .Q ( signal_12794 ) ) ;

    /* cells in depth 29 */
    buf_clk cell_7017 ( .C ( clk ), .D ( signal_12608 ), .Q ( signal_12609 ) ) ;
    buf_clk cell_7031 ( .C ( clk ), .D ( signal_12622 ), .Q ( signal_12623 ) ) ;
    buf_clk cell_7045 ( .C ( clk ), .D ( signal_12636 ), .Q ( signal_12637 ) ) ;
    buf_clk cell_7057 ( .C ( clk ), .D ( signal_12648 ), .Q ( signal_12649 ) ) ;
    buf_clk cell_7071 ( .C ( clk ), .D ( signal_12662 ), .Q ( signal_12663 ) ) ;
    buf_clk cell_7085 ( .C ( clk ), .D ( signal_12676 ), .Q ( signal_12677 ) ) ;
    buf_clk cell_7089 ( .C ( clk ), .D ( signal_23 ), .Q ( signal_12681 ) ) ;
    buf_clk cell_7095 ( .C ( clk ), .D ( signal_5286 ), .Q ( signal_12687 ) ) ;
    buf_clk cell_7101 ( .C ( clk ), .D ( signal_5287 ), .Q ( signal_12693 ) ) ;
    buf_clk cell_7107 ( .C ( clk ), .D ( signal_24 ), .Q ( signal_12699 ) ) ;
    buf_clk cell_7113 ( .C ( clk ), .D ( signal_5306 ), .Q ( signal_12705 ) ) ;
    buf_clk cell_7119 ( .C ( clk ), .D ( signal_5307 ), .Q ( signal_12711 ) ) ;
    buf_clk cell_7139 ( .C ( clk ), .D ( signal_12730 ), .Q ( signal_12731 ) ) ;
    buf_clk cell_7147 ( .C ( clk ), .D ( signal_12738 ), .Q ( signal_12739 ) ) ;
    buf_clk cell_7155 ( .C ( clk ), .D ( signal_12746 ), .Q ( signal_12747 ) ) ;
    buf_clk cell_7163 ( .C ( clk ), .D ( signal_12754 ), .Q ( signal_12755 ) ) ;
    buf_clk cell_7171 ( .C ( clk ), .D ( signal_12762 ), .Q ( signal_12763 ) ) ;
    buf_clk cell_7179 ( .C ( clk ), .D ( signal_12770 ), .Q ( signal_12771 ) ) ;
    buf_clk cell_7187 ( .C ( clk ), .D ( signal_12778 ), .Q ( signal_12779 ) ) ;
    buf_clk cell_7195 ( .C ( clk ), .D ( signal_12786 ), .Q ( signal_12787 ) ) ;
    buf_clk cell_7203 ( .C ( clk ), .D ( signal_12794 ), .Q ( signal_12795 ) ) ;
    buf_clk cell_7209 ( .C ( clk ), .D ( signal_30 ), .Q ( signal_12801 ) ) ;
    buf_clk cell_7215 ( .C ( clk ), .D ( signal_5300 ), .Q ( signal_12807 ) ) ;
    buf_clk cell_7221 ( .C ( clk ), .D ( signal_5301 ), .Q ( signal_12813 ) ) ;

    /* cells in depth 30 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2379 ( .a ({signal_12560, signal_12552, signal_12544}), .b ({signal_5309, signal_5308, signal_2386}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625]}), .c ({signal_5313, signal_5312, signal_2388}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2380 ( .a ({signal_12596, signal_12584, signal_12572}), .b ({signal_5311, signal_5310, signal_2387}), .clk ( clk ), .r ({Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({signal_5315, signal_5314, signal_2389}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2381 ( .a ({signal_5313, signal_5312, signal_2388}), .b ({signal_5317, signal_5316, signal_25}) ) ;
    buf_clk cell_7018 ( .C ( clk ), .D ( signal_12609 ), .Q ( signal_12610 ) ) ;
    buf_clk cell_7032 ( .C ( clk ), .D ( signal_12623 ), .Q ( signal_12624 ) ) ;
    buf_clk cell_7046 ( .C ( clk ), .D ( signal_12637 ), .Q ( signal_12638 ) ) ;
    buf_clk cell_7058 ( .C ( clk ), .D ( signal_12649 ), .Q ( signal_12650 ) ) ;
    buf_clk cell_7072 ( .C ( clk ), .D ( signal_12663 ), .Q ( signal_12664 ) ) ;
    buf_clk cell_7086 ( .C ( clk ), .D ( signal_12677 ), .Q ( signal_12678 ) ) ;
    buf_clk cell_7090 ( .C ( clk ), .D ( signal_12681 ), .Q ( signal_12682 ) ) ;
    buf_clk cell_7096 ( .C ( clk ), .D ( signal_12687 ), .Q ( signal_12688 ) ) ;
    buf_clk cell_7102 ( .C ( clk ), .D ( signal_12693 ), .Q ( signal_12694 ) ) ;
    buf_clk cell_7108 ( .C ( clk ), .D ( signal_12699 ), .Q ( signal_12700 ) ) ;
    buf_clk cell_7114 ( .C ( clk ), .D ( signal_12705 ), .Q ( signal_12706 ) ) ;
    buf_clk cell_7120 ( .C ( clk ), .D ( signal_12711 ), .Q ( signal_12712 ) ) ;
    buf_clk cell_7140 ( .C ( clk ), .D ( signal_12731 ), .Q ( signal_12732 ) ) ;
    buf_clk cell_7148 ( .C ( clk ), .D ( signal_12739 ), .Q ( signal_12740 ) ) ;
    buf_clk cell_7156 ( .C ( clk ), .D ( signal_12747 ), .Q ( signal_12748 ) ) ;
    buf_clk cell_7164 ( .C ( clk ), .D ( signal_12755 ), .Q ( signal_12756 ) ) ;
    buf_clk cell_7172 ( .C ( clk ), .D ( signal_12763 ), .Q ( signal_12764 ) ) ;
    buf_clk cell_7180 ( .C ( clk ), .D ( signal_12771 ), .Q ( signal_12772 ) ) ;
    buf_clk cell_7188 ( .C ( clk ), .D ( signal_12779 ), .Q ( signal_12780 ) ) ;
    buf_clk cell_7196 ( .C ( clk ), .D ( signal_12787 ), .Q ( signal_12788 ) ) ;
    buf_clk cell_7204 ( .C ( clk ), .D ( signal_12795 ), .Q ( signal_12796 ) ) ;
    buf_clk cell_7210 ( .C ( clk ), .D ( signal_12801 ), .Q ( signal_12802 ) ) ;
    buf_clk cell_7216 ( .C ( clk ), .D ( signal_12807 ), .Q ( signal_12808 ) ) ;
    buf_clk cell_7222 ( .C ( clk ), .D ( signal_12813 ), .Q ( signal_12814 ) ) ;

    /* cells in depth 31 */
    buf_clk cell_7059 ( .C ( clk ), .D ( signal_12650 ), .Q ( signal_12651 ) ) ;
    buf_clk cell_7073 ( .C ( clk ), .D ( signal_12664 ), .Q ( signal_12665 ) ) ;
    buf_clk cell_7087 ( .C ( clk ), .D ( signal_12678 ), .Q ( signal_12679 ) ) ;
    buf_clk cell_7091 ( .C ( clk ), .D ( signal_12682 ), .Q ( signal_12683 ) ) ;
    buf_clk cell_7097 ( .C ( clk ), .D ( signal_12688 ), .Q ( signal_12689 ) ) ;
    buf_clk cell_7103 ( .C ( clk ), .D ( signal_12694 ), .Q ( signal_12695 ) ) ;
    buf_clk cell_7109 ( .C ( clk ), .D ( signal_12700 ), .Q ( signal_12701 ) ) ;
    buf_clk cell_7115 ( .C ( clk ), .D ( signal_12706 ), .Q ( signal_12707 ) ) ;
    buf_clk cell_7121 ( .C ( clk ), .D ( signal_12712 ), .Q ( signal_12713 ) ) ;
    buf_clk cell_7125 ( .C ( clk ), .D ( signal_25 ), .Q ( signal_12717 ) ) ;
    buf_clk cell_7129 ( .C ( clk ), .D ( signal_5316 ), .Q ( signal_12721 ) ) ;
    buf_clk cell_7133 ( .C ( clk ), .D ( signal_5317 ), .Q ( signal_12725 ) ) ;
    buf_clk cell_7141 ( .C ( clk ), .D ( signal_12732 ), .Q ( signal_12733 ) ) ;
    buf_clk cell_7149 ( .C ( clk ), .D ( signal_12740 ), .Q ( signal_12741 ) ) ;
    buf_clk cell_7157 ( .C ( clk ), .D ( signal_12748 ), .Q ( signal_12749 ) ) ;
    buf_clk cell_7165 ( .C ( clk ), .D ( signal_12756 ), .Q ( signal_12757 ) ) ;
    buf_clk cell_7173 ( .C ( clk ), .D ( signal_12764 ), .Q ( signal_12765 ) ) ;
    buf_clk cell_7181 ( .C ( clk ), .D ( signal_12772 ), .Q ( signal_12773 ) ) ;
    buf_clk cell_7189 ( .C ( clk ), .D ( signal_12780 ), .Q ( signal_12781 ) ) ;
    buf_clk cell_7197 ( .C ( clk ), .D ( signal_12788 ), .Q ( signal_12789 ) ) ;
    buf_clk cell_7205 ( .C ( clk ), .D ( signal_12796 ), .Q ( signal_12797 ) ) ;
    buf_clk cell_7211 ( .C ( clk ), .D ( signal_12802 ), .Q ( signal_12803 ) ) ;
    buf_clk cell_7217 ( .C ( clk ), .D ( signal_12808 ), .Q ( signal_12809 ) ) ;
    buf_clk cell_7223 ( .C ( clk ), .D ( signal_12814 ), .Q ( signal_12815 ) ) ;

    /* cells in depth 32 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2382 ( .a ({signal_12638, signal_12624, signal_12610}), .b ({signal_5315, signal_5314, signal_2389}), .clk ( clk ), .r ({Fresh[2633], Fresh[2632], Fresh[2631]}), .c ({signal_5319, signal_5318, signal_2390}) ) ;
    buf_clk cell_7060 ( .C ( clk ), .D ( signal_12651 ), .Q ( signal_12652 ) ) ;
    buf_clk cell_7074 ( .C ( clk ), .D ( signal_12665 ), .Q ( signal_12666 ) ) ;
    buf_clk cell_7088 ( .C ( clk ), .D ( signal_12679 ), .Q ( signal_12680 ) ) ;
    buf_clk cell_7092 ( .C ( clk ), .D ( signal_12683 ), .Q ( signal_12684 ) ) ;
    buf_clk cell_7098 ( .C ( clk ), .D ( signal_12689 ), .Q ( signal_12690 ) ) ;
    buf_clk cell_7104 ( .C ( clk ), .D ( signal_12695 ), .Q ( signal_12696 ) ) ;
    buf_clk cell_7110 ( .C ( clk ), .D ( signal_12701 ), .Q ( signal_12702 ) ) ;
    buf_clk cell_7116 ( .C ( clk ), .D ( signal_12707 ), .Q ( signal_12708 ) ) ;
    buf_clk cell_7122 ( .C ( clk ), .D ( signal_12713 ), .Q ( signal_12714 ) ) ;
    buf_clk cell_7126 ( .C ( clk ), .D ( signal_12717 ), .Q ( signal_12718 ) ) ;
    buf_clk cell_7130 ( .C ( clk ), .D ( signal_12721 ), .Q ( signal_12722 ) ) ;
    buf_clk cell_7134 ( .C ( clk ), .D ( signal_12725 ), .Q ( signal_12726 ) ) ;
    buf_clk cell_7142 ( .C ( clk ), .D ( signal_12733 ), .Q ( signal_12734 ) ) ;
    buf_clk cell_7150 ( .C ( clk ), .D ( signal_12741 ), .Q ( signal_12742 ) ) ;
    buf_clk cell_7158 ( .C ( clk ), .D ( signal_12749 ), .Q ( signal_12750 ) ) ;
    buf_clk cell_7166 ( .C ( clk ), .D ( signal_12757 ), .Q ( signal_12758 ) ) ;
    buf_clk cell_7174 ( .C ( clk ), .D ( signal_12765 ), .Q ( signal_12766 ) ) ;
    buf_clk cell_7182 ( .C ( clk ), .D ( signal_12773 ), .Q ( signal_12774 ) ) ;
    buf_clk cell_7190 ( .C ( clk ), .D ( signal_12781 ), .Q ( signal_12782 ) ) ;
    buf_clk cell_7198 ( .C ( clk ), .D ( signal_12789 ), .Q ( signal_12790 ) ) ;
    buf_clk cell_7206 ( .C ( clk ), .D ( signal_12797 ), .Q ( signal_12798 ) ) ;
    buf_clk cell_7212 ( .C ( clk ), .D ( signal_12803 ), .Q ( signal_12804 ) ) ;
    buf_clk cell_7218 ( .C ( clk ), .D ( signal_12809 ), .Q ( signal_12810 ) ) ;
    buf_clk cell_7224 ( .C ( clk ), .D ( signal_12815 ), .Q ( signal_12816 ) ) ;

    /* cells in depth 33 */
    buf_clk cell_7093 ( .C ( clk ), .D ( signal_12684 ), .Q ( signal_12685 ) ) ;
    buf_clk cell_7099 ( .C ( clk ), .D ( signal_12690 ), .Q ( signal_12691 ) ) ;
    buf_clk cell_7105 ( .C ( clk ), .D ( signal_12696 ), .Q ( signal_12697 ) ) ;
    buf_clk cell_7111 ( .C ( clk ), .D ( signal_12702 ), .Q ( signal_12703 ) ) ;
    buf_clk cell_7117 ( .C ( clk ), .D ( signal_12708 ), .Q ( signal_12709 ) ) ;
    buf_clk cell_7123 ( .C ( clk ), .D ( signal_12714 ), .Q ( signal_12715 ) ) ;
    buf_clk cell_7127 ( .C ( clk ), .D ( signal_12718 ), .Q ( signal_12719 ) ) ;
    buf_clk cell_7131 ( .C ( clk ), .D ( signal_12722 ), .Q ( signal_12723 ) ) ;
    buf_clk cell_7135 ( .C ( clk ), .D ( signal_12726 ), .Q ( signal_12727 ) ) ;
    buf_clk cell_7143 ( .C ( clk ), .D ( signal_12734 ), .Q ( signal_12735 ) ) ;
    buf_clk cell_7151 ( .C ( clk ), .D ( signal_12742 ), .Q ( signal_12743 ) ) ;
    buf_clk cell_7159 ( .C ( clk ), .D ( signal_12750 ), .Q ( signal_12751 ) ) ;
    buf_clk cell_7167 ( .C ( clk ), .D ( signal_12758 ), .Q ( signal_12759 ) ) ;
    buf_clk cell_7175 ( .C ( clk ), .D ( signal_12766 ), .Q ( signal_12767 ) ) ;
    buf_clk cell_7183 ( .C ( clk ), .D ( signal_12774 ), .Q ( signal_12775 ) ) ;
    buf_clk cell_7191 ( .C ( clk ), .D ( signal_12782 ), .Q ( signal_12783 ) ) ;
    buf_clk cell_7199 ( .C ( clk ), .D ( signal_12790 ), .Q ( signal_12791 ) ) ;
    buf_clk cell_7207 ( .C ( clk ), .D ( signal_12798 ), .Q ( signal_12799 ) ) ;
    buf_clk cell_7213 ( .C ( clk ), .D ( signal_12804 ), .Q ( signal_12805 ) ) ;
    buf_clk cell_7219 ( .C ( clk ), .D ( signal_12810 ), .Q ( signal_12811 ) ) ;
    buf_clk cell_7225 ( .C ( clk ), .D ( signal_12816 ), .Q ( signal_12817 ) ) ;

    /* cells in depth 34 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_2383 ( .a ({signal_12680, signal_12666, signal_12652}), .b ({signal_5319, signal_5318, signal_2390}), .clk ( clk ), .r ({Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({signal_5321, signal_5320, signal_2391}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_2384 ( .a ({signal_5321, signal_5320, signal_2391}), .b ({signal_5323, signal_5322, signal_27}) ) ;
    buf_clk cell_7094 ( .C ( clk ), .D ( signal_12685 ), .Q ( signal_12686 ) ) ;
    buf_clk cell_7100 ( .C ( clk ), .D ( signal_12691 ), .Q ( signal_12692 ) ) ;
    buf_clk cell_7106 ( .C ( clk ), .D ( signal_12697 ), .Q ( signal_12698 ) ) ;
    buf_clk cell_7112 ( .C ( clk ), .D ( signal_12703 ), .Q ( signal_12704 ) ) ;
    buf_clk cell_7118 ( .C ( clk ), .D ( signal_12709 ), .Q ( signal_12710 ) ) ;
    buf_clk cell_7124 ( .C ( clk ), .D ( signal_12715 ), .Q ( signal_12716 ) ) ;
    buf_clk cell_7128 ( .C ( clk ), .D ( signal_12719 ), .Q ( signal_12720 ) ) ;
    buf_clk cell_7132 ( .C ( clk ), .D ( signal_12723 ), .Q ( signal_12724 ) ) ;
    buf_clk cell_7136 ( .C ( clk ), .D ( signal_12727 ), .Q ( signal_12728 ) ) ;
    buf_clk cell_7144 ( .C ( clk ), .D ( signal_12735 ), .Q ( signal_12736 ) ) ;
    buf_clk cell_7152 ( .C ( clk ), .D ( signal_12743 ), .Q ( signal_12744 ) ) ;
    buf_clk cell_7160 ( .C ( clk ), .D ( signal_12751 ), .Q ( signal_12752 ) ) ;
    buf_clk cell_7168 ( .C ( clk ), .D ( signal_12759 ), .Q ( signal_12760 ) ) ;
    buf_clk cell_7176 ( .C ( clk ), .D ( signal_12767 ), .Q ( signal_12768 ) ) ;
    buf_clk cell_7184 ( .C ( clk ), .D ( signal_12775 ), .Q ( signal_12776 ) ) ;
    buf_clk cell_7192 ( .C ( clk ), .D ( signal_12783 ), .Q ( signal_12784 ) ) ;
    buf_clk cell_7200 ( .C ( clk ), .D ( signal_12791 ), .Q ( signal_12792 ) ) ;
    buf_clk cell_7208 ( .C ( clk ), .D ( signal_12799 ), .Q ( signal_12800 ) ) ;
    buf_clk cell_7214 ( .C ( clk ), .D ( signal_12805 ), .Q ( signal_12806 ) ) ;
    buf_clk cell_7220 ( .C ( clk ), .D ( signal_12811 ), .Q ( signal_12812 ) ) ;
    buf_clk cell_7226 ( .C ( clk ), .D ( signal_12817 ), .Q ( signal_12818 ) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_12698, signal_12692, signal_12686}), .Q ({SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_12716, signal_12710, signal_12704}), .Q ({SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_12728, signal_12724, signal_12720}), .Q ({SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_12752, signal_12744, signal_12736}), .Q ({SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_5323, signal_5322, signal_27}), .Q ({SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_12776, signal_12768, signal_12760}), .Q ({SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_12800, signal_12792, signal_12784}), .Q ({SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_12818, signal_12812, signal_12806}), .Q ({SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
