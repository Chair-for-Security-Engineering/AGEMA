/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_AIG_ClockGating_d1 (X_s0, clk, X_s1, Fresh, rst, Y_s0, Y_s1, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input rst ;
    input [87:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output Synch ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_441 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_794 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(0)) cell_176 ( .a ({X_s1[0], X_s0[0]}), .b ({signal_438, signal_192}) ) ;
    INV_X1 cell_177 ( .A ( 1'b1 ), .ZN ( signal_193 ) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_178 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[4], X_s0[4]}), .c ({signal_441, signal_194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[5], X_s0[5]}), .c ({signal_444, signal_195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[4], X_s0[4]}), .c ({signal_445, signal_196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_446, signal_197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .a ({X_s1[3], X_s0[3]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_448, signal_198}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_183 ( .a ({signal_445, signal_196}), .b ({signal_449, signal_199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .a ({X_s1[6], X_s0[6]}), .b ({signal_445, signal_196}), .c ({signal_452, signal_202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_187 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_444, signal_195}), .c ({signal_454, signal_203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_188 ( .a ({signal_444, signal_195}), .b ({signal_446, signal_197}), .c ({signal_455, signal_204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_189 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_446, signal_197}), .c ({signal_457, signal_205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_190 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_448, signal_198}), .c ({signal_458, signal_206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_191 ( .a ({X_s1[5], X_s0[5]}), .b ({signal_446, signal_197}), .c ({signal_459, signal_207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_192 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_448, signal_198}), .c ({signal_460, signal_208}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_193 ( .a ({signal_455, signal_204}), .b ({signal_461, signal_209}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_194 ( .a ({signal_459, signal_207}), .b ({signal_462, signal_210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_201 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_459, signal_207}), .c ({signal_469, signal_217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_202 ( .a ({signal_454, signal_203}), .b ({signal_457, signal_205}), .c ({signal_470, signal_218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_203 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_457, signal_205}), .c ({signal_471, signal_219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_204 ( .a ({X_s1[3], X_s0[3]}), .b ({signal_457, signal_205}), .c ({signal_472, signal_220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_205 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_459, signal_207}), .c ({signal_473, signal_221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_206 ( .a ({signal_445, signal_196}), .b ({signal_460, signal_208}), .c ({signal_474, signal_222}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_208 ( .a ({signal_469, signal_217}), .b ({signal_476, signal_224}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_209 ( .a ({signal_470, signal_218}), .b ({signal_477, signal_225}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_210 ( .a ({signal_473, signal_221}), .b ({signal_478, signal_226}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_211 ( .a ({signal_474, signal_222}), .b ({signal_479, signal_227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_219 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_472, signal_220}), .c ({signal_487, signal_235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_220 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_473, signal_221}), .c ({signal_488, signal_236}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_222 ( .a ({signal_487, signal_235}), .b ({signal_490, signal_238}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_223 ( .a ({signal_488, signal_236}), .b ({signal_491, signal_239}) ) ;
    ClockGatingController #(17) cell_429 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_794 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .a ({signal_438, signal_192}), .b ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_450, signal_200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .a ({1'b0, signal_193}), .b ({signal_441, signal_194}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_451, signal_201}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_195 ( .a ({signal_450, signal_200}), .b ({signal_463, signal_211}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_196 ( .a ({signal_451, signal_201}), .b ({signal_464, signal_212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_197 ( .a ({1'b0, signal_193}), .b ({signal_454, signal_203}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_465, signal_213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_198 ( .a ({1'b0, signal_193}), .b ({signal_458, signal_206}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_466, signal_214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_199 ( .a ({1'b0, signal_193}), .b ({signal_449, signal_199}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_467, signal_215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_200 ( .a ({1'b0, signal_193}), .b ({signal_452, signal_202}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_468, signal_216}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_207 ( .a ({signal_465, signal_213}), .b ({signal_475, signal_223}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_212 ( .a ({signal_466, signal_214}), .b ({signal_480, signal_228}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_213 ( .a ({signal_467, signal_215}), .b ({signal_481, signal_229}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_214 ( .a ({signal_468, signal_216}), .b ({signal_482, signal_230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_215 ( .a ({1'b0, 1'b1}), .b ({signal_462, signal_210}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_483, signal_231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_216 ( .a ({1'b0, signal_193}), .b ({signal_471, signal_219}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_484, signal_232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_217 ( .a ({1'b0, signal_193}), .b ({signal_472, signal_220}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_485, signal_233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_218 ( .a ({1'b0, 1'b1}), .b ({signal_461, signal_209}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_486, signal_234}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_221 ( .a ({signal_483, signal_231}), .b ({signal_489, signal_237}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_224 ( .a ({signal_484, signal_232}), .b ({signal_492, signal_240}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_225 ( .a ({signal_485, signal_233}), .b ({signal_493, signal_241}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_226 ( .a ({signal_486, signal_234}), .b ({signal_494, signal_242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_228 ( .a ({1'b0, 1'b1}), .b ({signal_477, signal_225}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_496, signal_244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_229 ( .a ({1'b0, 1'b1}), .b ({signal_478, signal_226}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_497, signal_245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_230 ( .a ({1'b0, 1'b1}), .b ({signal_476, signal_224}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_498, signal_246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_231 ( .a ({1'b0, 1'b1}), .b ({signal_479, signal_227}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_499, signal_247}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_232 ( .a ({signal_496, signal_244}), .b ({signal_500, signal_248}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_233 ( .a ({signal_497, signal_245}), .b ({signal_501, signal_249}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_234 ( .a ({signal_498, signal_246}), .b ({signal_502, signal_250}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_235 ( .a ({signal_499, signal_247}), .b ({signal_503, signal_251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({1'b0, signal_193}), .b ({signal_491, signal_239}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_506, signal_254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({1'b0, 1'b1}), .b ({signal_490, signal_238}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_507, signal_255}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_241 ( .a ({signal_506, signal_254}), .b ({signal_509, signal_257}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_242 ( .a ({signal_507, signal_255}), .b ({signal_510, signal_258}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_227 ( .a ({signal_475, signal_223}), .b ({signal_463, signal_211}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_495, signal_243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({signal_480, signal_228}), .b ({signal_489, signal_237}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_504, signal_252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({signal_493, signal_241}), .b ({signal_494, signal_242}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_505, signal_253}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_240 ( .a ({signal_505, signal_253}), .b ({signal_508, signal_256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({signal_481, signal_229}), .b ({signal_500, signal_248}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_511, signal_259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({signal_492, signal_240}), .b ({signal_501, signal_249}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_512, signal_260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({signal_464, signal_212}), .b ({signal_502, signal_250}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_513, signal_261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({signal_482, signal_230}), .b ({signal_503, signal_251}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_514, signal_262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({signal_509, signal_257}), .b ({signal_510, signal_258}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_515, signal_263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({signal_495, signal_243}), .b ({signal_514, signal_262}), .c ({signal_519, signal_267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({signal_504, signal_252}), .b ({signal_514, signal_262}), .c ({signal_520, signal_268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({signal_513, signal_261}), .b ({signal_505, signal_253}), .c ({signal_521, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({signal_511, signal_259}), .b ({signal_512, signal_260}), .c ({signal_522, signal_270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({signal_512, signal_260}), .b ({signal_505, signal_253}), .c ({signal_523, signal_271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({signal_511, signal_259}), .b ({signal_513, signal_261}), .c ({signal_524, signal_272}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_257 ( .a ({signal_515, signal_263}), .b ({signal_525, signal_273}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_258 ( .a ({signal_520, signal_268}), .b ({signal_526, signal_274}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_259 ( .a ({signal_521, signal_269}), .b ({signal_527, signal_275}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_260 ( .a ({signal_523, signal_271}), .b ({signal_528, signal_276}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_261 ( .a ({signal_524, signal_272}), .b ({signal_529, signal_277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({signal_504, signal_252}), .b ({signal_515, signal_263}), .c ({signal_532, signal_280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({signal_495, signal_243}), .b ({signal_515, signal_263}), .c ({signal_533, signal_281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({signal_523, signal_271}), .b ({signal_524, signal_272}), .c ({signal_534, signal_282}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_267 ( .a ({signal_532, signal_280}), .b ({signal_535, signal_283}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_268 ( .a ({signal_533, signal_281}), .b ({signal_536, signal_284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({signal_520, signal_268}), .b ({signal_533, signal_281}), .c ({signal_541, signal_289}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({signal_511, signal_259}), .b ({signal_514, signal_262}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_516, signal_264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({signal_495, signal_243}), .b ({signal_512, signal_260}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_517, signal_265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({signal_504, signal_252}), .b ({signal_513, signal_261}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_518, signal_266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({signal_519, signal_267}), .b ({signal_522, signal_270}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_530, signal_278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({signal_520, signal_268}), .b ({signal_524, signal_272}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_531, signal_279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({signal_526, signal_274}), .b ({signal_529, signal_277}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_537, signal_285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({signal_508, signal_256}), .b ({signal_525, signal_273}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_538, signal_286}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({signal_521, signal_269}), .b ({signal_532, signal_280}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_539, signal_287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({signal_523, signal_271}), .b ({signal_533, signal_281}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_540, signal_288}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({signal_528, signal_276}), .b ({signal_536, signal_284}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_542, signal_290}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({signal_527, signal_275}), .b ({signal_535, signal_283}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_543, signal_291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({signal_534, signal_282}), .b ({signal_541, signal_289}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_544, signal_292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({signal_517, signal_265}), .b ({signal_537, signal_285}), .c ({signal_545, signal_293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({signal_530, signal_278}), .b ({signal_540, signal_288}), .c ({signal_546, signal_294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({signal_538, signal_286}), .b ({signal_539, signal_287}), .c ({signal_547, signal_295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_280 ( .a ({signal_516, signal_264}), .b ({signal_542, signal_290}), .c ({signal_548, signal_296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_281 ( .a ({signal_518, signal_266}), .b ({signal_543, signal_291}), .c ({signal_549, signal_297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_282 ( .a ({signal_530, signal_278}), .b ({signal_544, signal_292}), .c ({signal_550, signal_298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_283 ( .a ({signal_545, signal_293}), .b ({signal_546, signal_294}), .c ({signal_551, signal_299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_284 ( .a ({signal_540, signal_288}), .b ({signal_544, signal_292}), .c ({signal_552, signal_300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_285 ( .a ({signal_531, signal_279}), .b ({signal_547, signal_295}), .c ({signal_553, signal_301}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_286 ( .a ({signal_551, signal_299}), .b ({signal_554, signal_302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_287 ( .a ({signal_548, signal_296}), .b ({signal_550, signal_298}), .c ({signal_555, signal_303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_288 ( .a ({signal_549, signal_297}), .b ({signal_552, signal_300}), .c ({signal_556, signal_304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_289 ( .a ({signal_540, signal_288}), .b ({signal_553, signal_301}), .c ({signal_557, signal_305}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_290 ( .a ({signal_555, signal_303}), .b ({signal_558, signal_306}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_291 ( .a ({signal_556, signal_304}), .b ({signal_559, signal_307}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_292 ( .a ({signal_557, signal_305}), .b ({signal_560, signal_308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_294 ( .a ({signal_551, signal_299}), .b ({signal_555, signal_303}), .c ({signal_562, signal_310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_295 ( .a ({signal_556, signal_304}), .b ({signal_557, signal_305}), .c ({signal_563, signal_311}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_296 ( .a ({signal_562, signal_310}), .b ({signal_564, signal_312}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_297 ( .a ({signal_563, signal_311}), .b ({signal_565, signal_313}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_293 ( .a ({signal_555, signal_303}), .b ({signal_556, signal_304}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_561, signal_309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_298 ( .a ({signal_554, signal_302}), .b ({signal_560, signal_308}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_566, signal_314}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_299 ( .a ({signal_562, signal_310}), .b ({signal_563, signal_311}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_567, signal_315}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_300 ( .a ({signal_564, signal_312}), .b ({signal_565, signal_313}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_568, signal_316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_301 ( .a ({signal_561, signal_309}), .b ({signal_567, signal_315}), .c ({signal_569, signal_317}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_302 ( .a ({signal_569, signal_317}), .b ({signal_570, signal_318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_303 ( .a ({signal_566, signal_314}), .b ({signal_568, signal_316}), .c ({signal_571, signal_319}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_304 ( .a ({signal_571, signal_319}), .b ({signal_572, signal_320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_307 ( .a ({signal_569, signal_317}), .b ({signal_571, signal_319}), .c ({signal_575, signal_323}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_305 ( .a ({signal_560, signal_308}), .b ({signal_570, signal_318}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_573, signal_321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_306 ( .a ({signal_554, signal_302}), .b ({signal_570, signal_318}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_574, signal_322}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_308 ( .a ({signal_559, signal_307}), .b ({signal_572, signal_320}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_576, signal_324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_309 ( .a ({signal_558, signal_306}), .b ({signal_572, signal_320}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_577, signal_325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_310 ( .a ({signal_563, signal_311}), .b ({signal_575, signal_323}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_578, signal_326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_311 ( .a ({signal_562, signal_310}), .b ({signal_575, signal_323}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_579, signal_327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_312 ( .a ({signal_576, signal_324}), .b ({signal_578, signal_326}), .c ({signal_580, signal_328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_313 ( .a ({signal_573, signal_321}), .b ({signal_578, signal_326}), .c ({signal_581, signal_329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_314 ( .a ({signal_577, signal_325}), .b ({signal_579, signal_327}), .c ({signal_582, signal_330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_315 ( .a ({signal_574, signal_322}), .b ({signal_579, signal_327}), .c ({signal_583, signal_331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_324 ( .a ({signal_582, signal_330}), .b ({signal_583, signal_331}), .c ({signal_592, signal_340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_325 ( .a ({signal_580, signal_328}), .b ({signal_581, signal_329}), .c ({signal_593, signal_341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_326 ( .a ({signal_581, signal_329}), .b ({signal_583, signal_331}), .c ({signal_594, signal_342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_327 ( .a ({signal_580, signal_328}), .b ({signal_582, signal_330}), .c ({signal_595, signal_343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_336 ( .a ({signal_594, signal_342}), .b ({signal_595, signal_343}), .c ({signal_604, signal_352}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_316 ( .a ({signal_514, signal_262}), .b ({signal_580, signal_328}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_584, signal_332}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_317 ( .a ({signal_495, signal_243}), .b ({signal_581, signal_329}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_585, signal_333}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_318 ( .a ({signal_504, signal_252}), .b ({signal_582, signal_330}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_586, signal_334}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_319 ( .a ({signal_515, signal_263}), .b ({signal_583, signal_331}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_587, signal_335}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_320 ( .a ({signal_511, signal_259}), .b ({signal_580, signal_328}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_588, signal_336}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_321 ( .a ({signal_512, signal_260}), .b ({signal_581, signal_329}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_589, signal_337}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_322 ( .a ({signal_513, signal_261}), .b ({signal_582, signal_330}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_590, signal_338}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_323 ( .a ({signal_505, signal_253}), .b ({signal_583, signal_331}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_591, signal_339}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_328 ( .a ({signal_519, signal_267}), .b ({signal_593, signal_341}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_596, signal_344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_329 ( .a ({signal_532, signal_280}), .b ({signal_592, signal_340}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_597, signal_345}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_330 ( .a ({signal_520, signal_268}), .b ({signal_595, signal_343}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_598, signal_346}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_331 ( .a ({signal_533, signal_281}), .b ({signal_594, signal_342}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_599, signal_347}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_332 ( .a ({signal_522, signal_270}), .b ({signal_593, signal_341}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_600, signal_348}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_333 ( .a ({signal_521, signal_269}), .b ({signal_592, signal_340}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_601, signal_349}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_334 ( .a ({signal_524, signal_272}), .b ({signal_595, signal_343}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_602, signal_350}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_335 ( .a ({signal_523, signal_271}), .b ({signal_594, signal_342}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_603, signal_351}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_337 ( .a ({signal_541, signal_289}), .b ({signal_604, signal_352}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_605, signal_353}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_338 ( .a ({signal_534, signal_282}), .b ({signal_604, signal_352}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_606, signal_354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_339 ( .a ({signal_584, signal_332}), .b ({signal_596, signal_344}), .c ({signal_607, signal_355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_340 ( .a ({signal_585, signal_333}), .b ({signal_596, signal_344}), .c ({signal_608, signal_356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_341 ( .a ({signal_586, signal_334}), .b ({signal_597, signal_345}), .c ({signal_609, signal_357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_342 ( .a ({signal_587, signal_335}), .b ({signal_597, signal_345}), .c ({signal_610, signal_358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_343 ( .a ({signal_598, signal_346}), .b ({signal_599, signal_347}), .c ({signal_611, signal_359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_344 ( .a ({signal_588, signal_336}), .b ({signal_600, signal_348}), .c ({signal_612, signal_360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_345 ( .a ({signal_589, signal_337}), .b ({signal_600, signal_348}), .c ({signal_613, signal_361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_346 ( .a ({signal_590, signal_338}), .b ({signal_601, signal_349}), .c ({signal_614, signal_362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_347 ( .a ({signal_591, signal_339}), .b ({signal_601, signal_349}), .c ({signal_615, signal_363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_348 ( .a ({signal_602, signal_350}), .b ({signal_603, signal_351}), .c ({signal_616, signal_364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_349 ( .a ({signal_608, signal_356}), .b ({signal_611, signal_359}), .c ({signal_617, signal_365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_350 ( .a ({signal_610, signal_358}), .b ({signal_611, signal_359}), .c ({signal_618, signal_366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_351 ( .a ({signal_599, signal_347}), .b ({signal_605, signal_353}), .c ({signal_619, signal_367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_352 ( .a ({signal_613, signal_361}), .b ({signal_616, signal_364}), .c ({signal_620, signal_368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_353 ( .a ({signal_615, signal_363}), .b ({signal_616, signal_364}), .c ({signal_621, signal_369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_354 ( .a ({signal_603, signal_351}), .b ({signal_606, signal_354}), .c ({signal_622, signal_370}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_355 ( .a ({signal_620, signal_368}), .b ({signal_623, signal_371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_356 ( .a ({signal_617, signal_365}), .b ({signal_621, signal_369}), .c ({signal_624, signal_372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_357 ( .a ({signal_617, signal_365}), .b ({signal_618, signal_366}), .c ({signal_625, signal_373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_358 ( .a ({signal_607, signal_355}), .b ({signal_619, signal_367}), .c ({signal_626, signal_374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_359 ( .a ({signal_609, signal_357}), .b ({signal_619, signal_367}), .c ({signal_627, signal_375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_360 ( .a ({signal_612, signal_360}), .b ({signal_622, signal_370}), .c ({signal_628, signal_376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_361 ( .a ({signal_614, signal_362}), .b ({signal_622, signal_370}), .c ({signal_629, signal_377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_364 ( .a ({signal_627, signal_375}), .b ({signal_629, signal_377}), .c ({signal_632, signal_380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_365 ( .a ({signal_618, signal_366}), .b ({signal_629, signal_377}), .c ({signal_633, signal_381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_366 ( .a ({signal_617, signal_365}), .b ({signal_629, signal_377}), .c ({signal_634, signal_382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_367 ( .a ({signal_626, signal_374}), .b ({signal_628, signal_376}), .c ({signal_635, signal_383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_368 ( .a ({signal_627, signal_375}), .b ({signal_628, signal_376}), .c ({signal_636, signal_384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_369 ( .a ({signal_625, signal_373}), .b ({signal_629, signal_377}), .c ({signal_637, signal_385}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_370 ( .a ({signal_632, signal_380}), .b ({signal_638, signal_386}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_371 ( .a ({signal_633, signal_381}), .b ({signal_639, signal_387}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_372 ( .a ({signal_634, signal_382}), .b ({signal_640, signal_388}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_373 ( .a ({signal_636, signal_384}), .b ({signal_641, signal_389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_378 ( .a ({signal_618, signal_366}), .b ({signal_632, signal_380}), .c ({signal_646, signal_394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_379 ( .a ({signal_627, signal_375}), .b ({signal_635, signal_383}), .c ({signal_647, signal_395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_380 ( .a ({signal_620, signal_368}), .b ({signal_636, signal_384}), .c ({signal_648, signal_396}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_381 ( .a ({signal_647, signal_395}), .b ({signal_649, signal_397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_389 ( .a ({signal_626, signal_374}), .b ({signal_646, signal_394}), .c ({signal_657, signal_405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_390 ( .a ({signal_624, signal_372}), .b ({signal_647, signal_395}), .c ({signal_658, signal_406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_391 ( .a ({signal_637, signal_385}), .b ({signal_648, signal_396}), .c ({signal_659, signal_407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_392 ( .a ({signal_625, signal_373}), .b ({signal_647, signal_395}), .c ({signal_660, signal_408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_393 ( .a ({signal_624, signal_372}), .b ({signal_648, signal_396}), .c ({signal_661, signal_409}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_396 ( .a ({signal_657, signal_405}), .b ({signal_664, signal_412}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_397 ( .a ({signal_659, signal_407}), .b ({signal_665, signal_413}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_398 ( .a ({signal_660, signal_408}), .b ({signal_666, signal_414}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_399 ( .a ({signal_661, signal_409}), .b ({signal_667, signal_415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_405 ( .a ({signal_629, signal_377}), .b ({signal_658, signal_406}), .c ({signal_673, signal_420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_406 ( .a ({signal_620, signal_368}), .b ({signal_658, signal_406}), .c ({signal_674, signal_421}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_408 ( .a ({signal_673, signal_420}), .b ({signal_676, signal_423}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_409 ( .a ({signal_674, signal_421}), .b ({signal_677, signal_424}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_362 ( .a ({1'b0, signal_193}), .b ({signal_623, signal_371}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_630, signal_378}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_363 ( .a ({1'b0, 1'b1}), .b ({signal_624, signal_372}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_631, signal_379}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_374 ( .a ({signal_630, signal_378}), .b ({signal_642, signal_390}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_375 ( .a ({signal_631, signal_379}), .b ({signal_643, signal_391}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_637, signal_385}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_644, signal_392}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_377 ( .a ({1'b0, 1'b1}), .b ({signal_635, signal_383}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_645, signal_393}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_382 ( .a ({signal_644, signal_392}), .b ({signal_650, signal_398}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_383 ( .a ({signal_645, signal_393}), .b ({signal_651, signal_399}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_384 ( .a ({1'b0, signal_193}), .b ({signal_639, signal_387}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_652, signal_400}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_385 ( .a ({1'b0, 1'b1}), .b ({signal_641, signal_389}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_653, signal_401}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_386 ( .a ({1'b0, signal_193}), .b ({signal_640, signal_388}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_654, signal_402}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_387 ( .a ({1'b0, signal_193}), .b ({signal_638, signal_386}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_655, signal_403}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_388 ( .a ({1'b0, 1'b1}), .b ({signal_646, signal_394}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_656, signal_404}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_394 ( .a ({signal_652, signal_400}), .b ({signal_662, signal_410}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_395 ( .a ({signal_653, signal_401}), .b ({signal_663, signal_411}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_400 ( .a ({signal_654, signal_402}), .b ({signal_668, signal_416}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_401 ( .a ({signal_655, signal_403}), .b ({signal_669, signal_417}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_402 ( .a ({signal_656, signal_404}), .b ({signal_670, signal_418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_404 ( .a ({1'b0, 1'b1}), .b ({signal_649, signal_397}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_672, signal_419}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_407 ( .a ({signal_672, signal_419}), .b ({signal_675, signal_422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_412 ( .a ({1'b0, signal_193}), .b ({signal_665, signal_413}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_680, signal_425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_413 ( .a ({1'b0, 1'b1}), .b ({signal_666, signal_414}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_681, signal_426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_414 ( .a ({1'b0, signal_193}), .b ({signal_664, signal_412}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_682, signal_427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_415 ( .a ({1'b0, 1'b1}), .b ({signal_667, signal_415}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_683, signal_428}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_416 ( .a ({signal_680, signal_425}), .b ({signal_684, signal_429}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_417 ( .a ({signal_681, signal_426}), .b ({signal_685, signal_430}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_418 ( .a ({signal_682, signal_427}), .b ({signal_686, signal_431}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_419 ( .a ({signal_683, signal_428}), .b ({signal_687, signal_432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_421 ( .a ({1'b0, signal_193}), .b ({signal_676, signal_423}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_689, signal_433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_422 ( .a ({1'b0, signal_193}), .b ({signal_677, signal_424}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_690, signal_434}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_423 ( .a ({signal_689, signal_433}), .b ({signal_691, signal_435}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_424 ( .a ({signal_690, signal_434}), .b ({signal_692, signal_436}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_403 ( .a ({signal_642, signal_390}), .b ({signal_650, signal_398}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_671, signal_167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_410 ( .a ({signal_662, signal_410}), .b ({signal_663, signal_411}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_678, signal_160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_411 ( .a ({signal_669, signal_417}), .b ({signal_670, signal_418}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_679, signal_166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_420 ( .a ({signal_668, signal_416}), .b ({signal_675, signal_422}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_688, signal_163}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_425 ( .a ({signal_684, signal_429}), .b ({signal_685, signal_430}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_693, signal_164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_426 ( .a ({signal_686, signal_431}), .b ({signal_687, signal_432}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_694, signal_165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_427 ( .a ({signal_691, signal_435}), .b ({signal_651, signal_399}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_695, signal_161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_428 ( .a ({signal_692, signal_436}), .b ({signal_643, signal_391}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_696, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_0 ( .clk ( signal_794 ), .D ({signal_678, signal_160}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1 ( .clk ( signal_794 ), .D ({signal_695, signal_161}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_2 ( .clk ( signal_794 ), .D ({signal_696, signal_162}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3 ( .clk ( signal_794 ), .D ({signal_688, signal_163}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_4 ( .clk ( signal_794 ), .D ({signal_693, signal_164}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_5 ( .clk ( signal_794 ), .D ({signal_694, signal_165}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_6 ( .clk ( signal_794 ), .D ({signal_679, signal_166}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_7 ( .clk ( signal_794 ), .D ({signal_671, signal_167}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
