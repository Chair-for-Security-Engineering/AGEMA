/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module Midori64_HPC2_AIG_ClockGating_d1 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, DataIn_s1, Fresh, DataOut_s0, done, DataOut_s1, Synch);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [63:0] DataIn_s1 ;
    input [255:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output Synch ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1954 ;
    wire signal_1957 ;
    wire signal_1960 ;
    wire signal_1963 ;
    wire signal_1966 ;
    wire signal_1969 ;
    wire signal_1972 ;
    wire signal_1975 ;
    wire signal_1978 ;
    wire signal_1981 ;
    wire signal_1984 ;
    wire signal_1987 ;
    wire signal_1990 ;
    wire signal_1993 ;
    wire signal_1996 ;
    wire signal_1999 ;
    wire signal_2002 ;
    wire signal_2005 ;
    wire signal_2008 ;
    wire signal_2011 ;
    wire signal_2014 ;
    wire signal_2017 ;
    wire signal_2020 ;
    wire signal_2023 ;
    wire signal_2026 ;
    wire signal_2029 ;
    wire signal_2032 ;
    wire signal_2035 ;
    wire signal_2038 ;
    wire signal_2041 ;
    wire signal_2044 ;
    wire signal_2047 ;
    wire signal_2050 ;
    wire signal_2053 ;
    wire signal_2056 ;
    wire signal_2059 ;
    wire signal_2062 ;
    wire signal_2065 ;
    wire signal_2068 ;
    wire signal_2071 ;
    wire signal_2074 ;
    wire signal_2077 ;
    wire signal_2080 ;
    wire signal_2083 ;
    wire signal_2086 ;
    wire signal_2089 ;
    wire signal_2092 ;
    wire signal_2095 ;
    wire signal_2098 ;
    wire signal_2101 ;
    wire signal_2104 ;
    wire signal_2107 ;
    wire signal_2110 ;
    wire signal_2113 ;
    wire signal_2116 ;
    wire signal_2119 ;
    wire signal_2122 ;
    wire signal_2125 ;
    wire signal_2128 ;
    wire signal_2131 ;
    wire signal_2134 ;
    wire signal_2137 ;
    wire signal_2140 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2318 ;
    wire signal_2320 ;
    wire signal_2322 ;
    wire signal_2324 ;
    wire signal_2326 ;
    wire signal_2328 ;
    wire signal_2330 ;
    wire signal_2332 ;
    wire signal_2334 ;
    wire signal_2336 ;
    wire signal_2338 ;
    wire signal_2340 ;
    wire signal_2342 ;
    wire signal_2344 ;
    wire signal_2346 ;
    wire signal_2348 ;
    wire signal_2350 ;
    wire signal_2352 ;
    wire signal_2354 ;
    wire signal_2356 ;
    wire signal_2358 ;
    wire signal_2360 ;
    wire signal_2362 ;
    wire signal_2364 ;
    wire signal_2366 ;
    wire signal_2368 ;
    wire signal_2370 ;
    wire signal_2372 ;
    wire signal_2374 ;
    wire signal_2376 ;
    wire signal_2378 ;
    wire signal_2380 ;
    wire signal_2382 ;
    wire signal_2384 ;
    wire signal_2386 ;
    wire signal_2388 ;
    wire signal_2390 ;
    wire signal_2392 ;
    wire signal_2394 ;
    wire signal_2396 ;
    wire signal_2398 ;
    wire signal_2400 ;
    wire signal_2402 ;
    wire signal_2404 ;
    wire signal_2406 ;
    wire signal_2408 ;
    wire signal_2410 ;
    wire signal_2412 ;
    wire signal_2414 ;
    wire signal_2416 ;
    wire signal_2418 ;
    wire signal_2420 ;
    wire signal_2422 ;
    wire signal_2424 ;
    wire signal_2426 ;
    wire signal_2428 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2434 ;
    wire signal_2436 ;
    wire signal_2438 ;
    wire signal_2440 ;
    wire signal_2442 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3712 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_0 ( .a ({key_s1[73], key_s0[73]}), .b ({key_s1[9], key_s0[9]}), .c ({signal_1954, signal_914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1 ( .a ({key_s1[72], key_s0[72]}), .b ({key_s1[8], key_s0[8]}), .c ({signal_1957, signal_915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2 ( .a ({key_s1[71], key_s0[71]}), .b ({key_s1[7], key_s0[7]}), .c ({signal_1960, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3 ( .a ({key_s1[6], key_s0[6]}), .b ({key_s1[70], key_s0[70]}), .c ({signal_1963, signal_917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4 ( .a ({key_s1[127], key_s0[127]}), .b ({key_s1[63], key_s0[63]}), .c ({signal_1966, signal_860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5 ( .a ({key_s1[126], key_s0[126]}), .b ({key_s1[62], key_s0[62]}), .c ({signal_1969, signal_861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6 ( .a ({key_s1[125], key_s0[125]}), .b ({key_s1[61], key_s0[61]}), .c ({signal_1972, signal_862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7 ( .a ({key_s1[124], key_s0[124]}), .b ({key_s1[60], key_s0[60]}), .c ({signal_1975, signal_863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_8 ( .a ({key_s1[5], key_s0[5]}), .b ({key_s1[69], key_s0[69]}), .c ({signal_1978, signal_918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_9 ( .a ({key_s1[123], key_s0[123]}), .b ({key_s1[59], key_s0[59]}), .c ({signal_1981, signal_864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_10 ( .a ({key_s1[122], key_s0[122]}), .b ({key_s1[58], key_s0[58]}), .c ({signal_1984, signal_865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_11 ( .a ({key_s1[121], key_s0[121]}), .b ({key_s1[57], key_s0[57]}), .c ({signal_1987, signal_866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_12 ( .a ({key_s1[120], key_s0[120]}), .b ({key_s1[56], key_s0[56]}), .c ({signal_1990, signal_867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_13 ( .a ({key_s1[119], key_s0[119]}), .b ({key_s1[55], key_s0[55]}), .c ({signal_1993, signal_868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_14 ( .a ({key_s1[118], key_s0[118]}), .b ({key_s1[54], key_s0[54]}), .c ({signal_1996, signal_869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_15 ( .a ({key_s1[117], key_s0[117]}), .b ({key_s1[53], key_s0[53]}), .c ({signal_1999, signal_870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_16 ( .a ({key_s1[116], key_s0[116]}), .b ({key_s1[52], key_s0[52]}), .c ({signal_2002, signal_871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_17 ( .a ({key_s1[115], key_s0[115]}), .b ({key_s1[51], key_s0[51]}), .c ({signal_2005, signal_872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_18 ( .a ({key_s1[114], key_s0[114]}), .b ({key_s1[50], key_s0[50]}), .c ({signal_2008, signal_873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_19 ( .a ({key_s1[4], key_s0[4]}), .b ({key_s1[68], key_s0[68]}), .c ({signal_2011, signal_919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_20 ( .a ({key_s1[113], key_s0[113]}), .b ({key_s1[49], key_s0[49]}), .c ({signal_2014, signal_874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_21 ( .a ({key_s1[112], key_s0[112]}), .b ({key_s1[48], key_s0[48]}), .c ({signal_2017, signal_875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_22 ( .a ({key_s1[111], key_s0[111]}), .b ({key_s1[47], key_s0[47]}), .c ({signal_2020, signal_876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_23 ( .a ({key_s1[110], key_s0[110]}), .b ({key_s1[46], key_s0[46]}), .c ({signal_2023, signal_877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_24 ( .a ({key_s1[109], key_s0[109]}), .b ({key_s1[45], key_s0[45]}), .c ({signal_2026, signal_878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_25 ( .a ({key_s1[108], key_s0[108]}), .b ({key_s1[44], key_s0[44]}), .c ({signal_2029, signal_879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_26 ( .a ({key_s1[107], key_s0[107]}), .b ({key_s1[43], key_s0[43]}), .c ({signal_2032, signal_880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_27 ( .a ({key_s1[106], key_s0[106]}), .b ({key_s1[42], key_s0[42]}), .c ({signal_2035, signal_881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_28 ( .a ({key_s1[105], key_s0[105]}), .b ({key_s1[41], key_s0[41]}), .c ({signal_2038, signal_882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_29 ( .a ({key_s1[104], key_s0[104]}), .b ({key_s1[40], key_s0[40]}), .c ({signal_2041, signal_883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_30 ( .a ({key_s1[3], key_s0[3]}), .b ({key_s1[67], key_s0[67]}), .c ({signal_2044, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_31 ( .a ({key_s1[103], key_s0[103]}), .b ({key_s1[39], key_s0[39]}), .c ({signal_2047, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_32 ( .a ({key_s1[102], key_s0[102]}), .b ({key_s1[38], key_s0[38]}), .c ({signal_2050, signal_885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_33 ( .a ({key_s1[101], key_s0[101]}), .b ({key_s1[37], key_s0[37]}), .c ({signal_2053, signal_886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_34 ( .a ({key_s1[100], key_s0[100]}), .b ({key_s1[36], key_s0[36]}), .c ({signal_2056, signal_887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_35 ( .a ({key_s1[35], key_s0[35]}), .b ({key_s1[99], key_s0[99]}), .c ({signal_2059, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_36 ( .a ({key_s1[34], key_s0[34]}), .b ({key_s1[98], key_s0[98]}), .c ({signal_2062, signal_889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_37 ( .a ({key_s1[33], key_s0[33]}), .b ({key_s1[97], key_s0[97]}), .c ({signal_2065, signal_890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_38 ( .a ({key_s1[32], key_s0[32]}), .b ({key_s1[96], key_s0[96]}), .c ({signal_2068, signal_891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_39 ( .a ({key_s1[31], key_s0[31]}), .b ({key_s1[95], key_s0[95]}), .c ({signal_2071, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_40 ( .a ({key_s1[30], key_s0[30]}), .b ({key_s1[94], key_s0[94]}), .c ({signal_2074, signal_893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_41 ( .a ({key_s1[2], key_s0[2]}), .b ({key_s1[66], key_s0[66]}), .c ({signal_2077, signal_921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_42 ( .a ({key_s1[29], key_s0[29]}), .b ({key_s1[93], key_s0[93]}), .c ({signal_2080, signal_894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_43 ( .a ({key_s1[28], key_s0[28]}), .b ({key_s1[92], key_s0[92]}), .c ({signal_2083, signal_895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_44 ( .a ({key_s1[27], key_s0[27]}), .b ({key_s1[91], key_s0[91]}), .c ({signal_2086, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_45 ( .a ({key_s1[26], key_s0[26]}), .b ({key_s1[90], key_s0[90]}), .c ({signal_2089, signal_897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_46 ( .a ({key_s1[25], key_s0[25]}), .b ({key_s1[89], key_s0[89]}), .c ({signal_2092, signal_898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_47 ( .a ({key_s1[24], key_s0[24]}), .b ({key_s1[88], key_s0[88]}), .c ({signal_2095, signal_899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_48 ( .a ({key_s1[23], key_s0[23]}), .b ({key_s1[87], key_s0[87]}), .c ({signal_2098, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_49 ( .a ({key_s1[22], key_s0[22]}), .b ({key_s1[86], key_s0[86]}), .c ({signal_2101, signal_901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_50 ( .a ({key_s1[21], key_s0[21]}), .b ({key_s1[85], key_s0[85]}), .c ({signal_2104, signal_902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_51 ( .a ({key_s1[20], key_s0[20]}), .b ({key_s1[84], key_s0[84]}), .c ({signal_2107, signal_903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_52 ( .a ({key_s1[1], key_s0[1]}), .b ({key_s1[65], key_s0[65]}), .c ({signal_2110, signal_922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_53 ( .a ({key_s1[19], key_s0[19]}), .b ({key_s1[83], key_s0[83]}), .c ({signal_2113, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_54 ( .a ({key_s1[18], key_s0[18]}), .b ({key_s1[82], key_s0[82]}), .c ({signal_2116, signal_905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_55 ( .a ({key_s1[17], key_s0[17]}), .b ({key_s1[81], key_s0[81]}), .c ({signal_2119, signal_906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_56 ( .a ({key_s1[16], key_s0[16]}), .b ({key_s1[80], key_s0[80]}), .c ({signal_2122, signal_907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_57 ( .a ({key_s1[15], key_s0[15]}), .b ({key_s1[79], key_s0[79]}), .c ({signal_2125, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_58 ( .a ({key_s1[14], key_s0[14]}), .b ({key_s1[78], key_s0[78]}), .c ({signal_2128, signal_909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_59 ( .a ({key_s1[13], key_s0[13]}), .b ({key_s1[77], key_s0[77]}), .c ({signal_2131, signal_910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_60 ( .a ({key_s1[12], key_s0[12]}), .b ({key_s1[76], key_s0[76]}), .c ({signal_2134, signal_911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_61 ( .a ({key_s1[11], key_s0[11]}), .b ({key_s1[75], key_s0[75]}), .c ({signal_2137, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_62 ( .a ({key_s1[10], key_s0[10]}), .b ({key_s1[74], key_s0[74]}), .c ({signal_2140, signal_913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_63 ( .a ({key_s1[0], key_s0[0]}), .b ({key_s1[64], key_s0[64]}), .c ({signal_2143, signal_923}) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_266), .A2 (signal_267), .ZN (done) ) ;
    NAND2_X1 cell_65 ( .A1 (signal_927), .A2 (signal_926), .ZN (signal_267) ) ;
    NAND2_X1 cell_66 ( .A1 (signal_925), .A2 (signal_924), .ZN (signal_266) ) ;
    INV_X1 cell_67 ( .A (signal_268), .ZN (signal_278) ) ;
    MUX2_X1 cell_68 ( .S (signal_281), .A (signal_269), .B (signal_270), .Z (signal_268) ) ;
    NOR2_X1 cell_69 ( .A1 (reset), .A2 (signal_271), .ZN (signal_282) ) ;
    XNOR2_X1 cell_70 ( .A (signal_927), .B (signal_926), .ZN (signal_271) ) ;
    MUX2_X1 cell_71 ( .S (signal_924), .A (signal_272), .B (signal_273), .Z (signal_280) ) ;
    NAND2_X1 cell_72 ( .A1 (signal_269), .A2 (signal_274), .ZN (signal_273) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_281), .A2 (signal_277), .ZN (signal_274) ) ;
    NOR2_X1 cell_74 ( .A1 (signal_275), .A2 (signal_283), .ZN (signal_269) ) ;
    NOR2_X1 cell_75 ( .A1 (signal_926), .A2 (reset), .ZN (signal_275) ) ;
    NOR2_X1 cell_76 ( .A1 (signal_281), .A2 (signal_270), .ZN (signal_272) ) ;
    NAND2_X1 cell_77 ( .A1 (signal_926), .A2 (signal_276), .ZN (signal_270) ) ;
    NOR2_X1 cell_78 ( .A1 (reset), .A2 (signal_279), .ZN (signal_276) ) ;
    NOR2_X1 cell_79 ( .A1 (reset), .A2 (signal_927), .ZN (signal_283) ) ;
    INV_X1 cell_80 ( .A (reset), .ZN (signal_277) ) ;
    INV_X1 cell_81 ( .A (signal_927), .ZN (signal_279) ) ;
    INV_X1 cell_85 ( .A (signal_925), .ZN (signal_281) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_153 ( .a ({signal_1954, signal_914}), .b ({DataIn_s1[9], DataIn_s0[9]}), .c ({signal_2318, signal_982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_154 ( .a ({signal_1957, signal_915}), .b ({DataIn_s1[8], DataIn_s0[8]}), .c ({signal_2320, signal_983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_155 ( .a ({signal_1960, signal_916}), .b ({DataIn_s1[7], DataIn_s0[7]}), .c ({signal_2322, signal_984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_156 ( .a ({signal_1963, signal_917}), .b ({DataIn_s1[6], DataIn_s0[6]}), .c ({signal_2324, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_157 ( .a ({signal_1966, signal_860}), .b ({DataIn_s1[63], DataIn_s0[63]}), .c ({signal_2326, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_158 ( .a ({signal_1969, signal_861}), .b ({DataIn_s1[62], DataIn_s0[62]}), .c ({signal_2328, signal_929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_159 ( .a ({signal_1972, signal_862}), .b ({DataIn_s1[61], DataIn_s0[61]}), .c ({signal_2330, signal_930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_160 ( .a ({signal_1975, signal_863}), .b ({DataIn_s1[60], DataIn_s0[60]}), .c ({signal_2332, signal_931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_161 ( .a ({signal_1978, signal_918}), .b ({DataIn_s1[5], DataIn_s0[5]}), .c ({signal_2334, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_162 ( .a ({signal_1981, signal_864}), .b ({DataIn_s1[59], DataIn_s0[59]}), .c ({signal_2336, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_163 ( .a ({signal_1984, signal_865}), .b ({DataIn_s1[58], DataIn_s0[58]}), .c ({signal_2338, signal_933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_164 ( .a ({signal_1987, signal_866}), .b ({DataIn_s1[57], DataIn_s0[57]}), .c ({signal_2340, signal_934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_165 ( .a ({signal_1990, signal_867}), .b ({DataIn_s1[56], DataIn_s0[56]}), .c ({signal_2342, signal_935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_166 ( .a ({signal_1993, signal_868}), .b ({DataIn_s1[55], DataIn_s0[55]}), .c ({signal_2344, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_167 ( .a ({signal_1996, signal_869}), .b ({DataIn_s1[54], DataIn_s0[54]}), .c ({signal_2346, signal_937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_168 ( .a ({signal_1999, signal_870}), .b ({DataIn_s1[53], DataIn_s0[53]}), .c ({signal_2348, signal_938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_169 ( .a ({signal_2002, signal_871}), .b ({DataIn_s1[52], DataIn_s0[52]}), .c ({signal_2350, signal_939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_170 ( .a ({signal_2005, signal_872}), .b ({DataIn_s1[51], DataIn_s0[51]}), .c ({signal_2352, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_171 ( .a ({signal_2008, signal_873}), .b ({DataIn_s1[50], DataIn_s0[50]}), .c ({signal_2354, signal_941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_172 ( .a ({signal_2011, signal_919}), .b ({DataIn_s1[4], DataIn_s0[4]}), .c ({signal_2356, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_173 ( .a ({signal_2014, signal_874}), .b ({DataIn_s1[49], DataIn_s0[49]}), .c ({signal_2358, signal_942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_174 ( .a ({signal_2017, signal_875}), .b ({DataIn_s1[48], DataIn_s0[48]}), .c ({signal_2360, signal_943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_175 ( .a ({signal_2020, signal_876}), .b ({DataIn_s1[47], DataIn_s0[47]}), .c ({signal_2362, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_176 ( .a ({signal_2023, signal_877}), .b ({DataIn_s1[46], DataIn_s0[46]}), .c ({signal_2364, signal_945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_177 ( .a ({signal_2026, signal_878}), .b ({DataIn_s1[45], DataIn_s0[45]}), .c ({signal_2366, signal_946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_178 ( .a ({signal_2029, signal_879}), .b ({DataIn_s1[44], DataIn_s0[44]}), .c ({signal_2368, signal_947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .a ({signal_2032, signal_880}), .b ({DataIn_s1[43], DataIn_s0[43]}), .c ({signal_2370, signal_948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .a ({signal_2035, signal_881}), .b ({DataIn_s1[42], DataIn_s0[42]}), .c ({signal_2372, signal_949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .a ({signal_2038, signal_882}), .b ({DataIn_s1[41], DataIn_s0[41]}), .c ({signal_2374, signal_950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .a ({signal_2041, signal_883}), .b ({DataIn_s1[40], DataIn_s0[40]}), .c ({signal_2376, signal_951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_183 ( .a ({signal_2044, signal_920}), .b ({DataIn_s1[3], DataIn_s0[3]}), .c ({signal_2378, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .a ({signal_2047, signal_884}), .b ({DataIn_s1[39], DataIn_s0[39]}), .c ({signal_2380, signal_952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .a ({signal_2050, signal_885}), .b ({DataIn_s1[38], DataIn_s0[38]}), .c ({signal_2382, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .a ({signal_2053, signal_886}), .b ({DataIn_s1[37], DataIn_s0[37]}), .c ({signal_2384, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_187 ( .a ({signal_2056, signal_887}), .b ({DataIn_s1[36], DataIn_s0[36]}), .c ({signal_2386, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_188 ( .a ({signal_2059, signal_888}), .b ({DataIn_s1[35], DataIn_s0[35]}), .c ({signal_2388, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_189 ( .a ({signal_2062, signal_889}), .b ({DataIn_s1[34], DataIn_s0[34]}), .c ({signal_2390, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_190 ( .a ({signal_2065, signal_890}), .b ({DataIn_s1[33], DataIn_s0[33]}), .c ({signal_2392, signal_958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_191 ( .a ({signal_2068, signal_891}), .b ({DataIn_s1[32], DataIn_s0[32]}), .c ({signal_2394, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_192 ( .a ({signal_2071, signal_892}), .b ({DataIn_s1[31], DataIn_s0[31]}), .c ({signal_2396, signal_960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_193 ( .a ({signal_2074, signal_893}), .b ({DataIn_s1[30], DataIn_s0[30]}), .c ({signal_2398, signal_961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_194 ( .a ({signal_2077, signal_921}), .b ({DataIn_s1[2], DataIn_s0[2]}), .c ({signal_2400, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_195 ( .a ({signal_2080, signal_894}), .b ({DataIn_s1[29], DataIn_s0[29]}), .c ({signal_2402, signal_962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_196 ( .a ({signal_2083, signal_895}), .b ({DataIn_s1[28], DataIn_s0[28]}), .c ({signal_2404, signal_963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_197 ( .a ({signal_2086, signal_896}), .b ({DataIn_s1[27], DataIn_s0[27]}), .c ({signal_2406, signal_964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_198 ( .a ({signal_2089, signal_897}), .b ({DataIn_s1[26], DataIn_s0[26]}), .c ({signal_2408, signal_965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_199 ( .a ({signal_2092, signal_898}), .b ({DataIn_s1[25], DataIn_s0[25]}), .c ({signal_2410, signal_966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_200 ( .a ({signal_2095, signal_899}), .b ({DataIn_s1[24], DataIn_s0[24]}), .c ({signal_2412, signal_967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_201 ( .a ({signal_2098, signal_900}), .b ({DataIn_s1[23], DataIn_s0[23]}), .c ({signal_2414, signal_968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_202 ( .a ({signal_2101, signal_901}), .b ({DataIn_s1[22], DataIn_s0[22]}), .c ({signal_2416, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_203 ( .a ({signal_2104, signal_902}), .b ({DataIn_s1[21], DataIn_s0[21]}), .c ({signal_2418, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_204 ( .a ({signal_2107, signal_903}), .b ({DataIn_s1[20], DataIn_s0[20]}), .c ({signal_2420, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_205 ( .a ({signal_2110, signal_922}), .b ({DataIn_s1[1], DataIn_s0[1]}), .c ({signal_2422, signal_990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_206 ( .a ({signal_2113, signal_904}), .b ({DataIn_s1[19], DataIn_s0[19]}), .c ({signal_2424, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_207 ( .a ({signal_2116, signal_905}), .b ({DataIn_s1[18], DataIn_s0[18]}), .c ({signal_2426, signal_973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_208 ( .a ({signal_2119, signal_906}), .b ({DataIn_s1[17], DataIn_s0[17]}), .c ({signal_2428, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_209 ( .a ({signal_2122, signal_907}), .b ({DataIn_s1[16], DataIn_s0[16]}), .c ({signal_2430, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_210 ( .a ({signal_2125, signal_908}), .b ({DataIn_s1[15], DataIn_s0[15]}), .c ({signal_2432, signal_976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_211 ( .a ({signal_2128, signal_909}), .b ({DataIn_s1[14], DataIn_s0[14]}), .c ({signal_2434, signal_977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_212 ( .a ({signal_2131, signal_910}), .b ({DataIn_s1[13], DataIn_s0[13]}), .c ({signal_2436, signal_978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_213 ( .a ({signal_2134, signal_911}), .b ({DataIn_s1[12], DataIn_s0[12]}), .c ({signal_2438, signal_979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_214 ( .a ({signal_2137, signal_912}), .b ({DataIn_s1[11], DataIn_s0[11]}), .c ({signal_2440, signal_980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_215 ( .a ({signal_2140, signal_913}), .b ({DataIn_s1[10], DataIn_s0[10]}), .c ({signal_2442, signal_981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_216 ( .a ({signal_2143, signal_923}), .b ({DataIn_s1[0], DataIn_s0[0]}), .c ({signal_2444, signal_991}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_283 ( .a ({signal_2149, signal_310}), .b ({1'b0, signal_1453}), .c ({signal_3088, signal_286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_290 ( .a ({signal_2588, signal_362}), .b ({1'b0, signal_1440}), .c ({signal_3120, signal_287}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_296 ( .a ({signal_2584, signal_358}), .b ({1'b0, signal_1441}), .c ({signal_3121, signal_288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_301 ( .a ({signal_2580, signal_354}), .b ({1'b0, signal_1442}), .c ({signal_3122, signal_289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_305 ( .a ({signal_2148, signal_306}), .b ({1'b0, signal_1454}), .c ({signal_3123, signal_290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_308 ( .a ({signal_2576, signal_350}), .b ({1'b0, signal_1443}), .c ({signal_3232, signal_291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_313 ( .a ({signal_2572, signal_346}), .b ({1'b0, signal_1444}), .c ({signal_3089, signal_292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_318 ( .a ({signal_2568, signal_342}), .b ({1'b0, signal_1445}), .c ({signal_3124, signal_293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_324 ( .a ({signal_2564, signal_338}), .b ({1'b0, signal_1446}), .c ({signal_3090, signal_294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_329 ( .a ({signal_2560, signal_334}), .b ({1'b0, signal_1447}), .c ({signal_3125, signal_295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_335 ( .a ({signal_2556, signal_330}), .b ({1'b0, signal_1448}), .c ({signal_3191, signal_296}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_340 ( .a ({signal_2553, signal_326}), .b ({1'b0, signal_1449}), .c ({signal_3126, signal_297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_345 ( .a ({signal_2549, signal_322}), .b ({1'b0, signal_1450}), .c ({signal_3091, signal_298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_351 ( .a ({signal_2545, signal_318}), .b ({1'b0, signal_1451}), .c ({signal_3127, signal_299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_356 ( .a ({signal_2544, signal_314}), .b ({1'b0, signal_1452}), .c ({signal_3128, signal_300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_360 ( .a ({signal_2144, signal_302}), .b ({1'b0, signal_1455}), .c ({signal_3129, signal_301}) ) ;
    NAND2_X1 cell_361 ( .A1 (signal_366), .A2 (signal_367), .ZN (signal_1446) ) ;
    NOR2_X1 cell_362 ( .A1 (signal_368), .A2 (signal_369), .ZN (signal_366) ) ;
    OR2_X1 cell_363 ( .A1 (signal_370), .A2 (signal_371), .ZN (signal_369) ) ;
    NAND2_X1 cell_364 ( .A1 (signal_372), .A2 (signal_373), .ZN (signal_1447) ) ;
    NAND2_X1 cell_365 ( .A1 (signal_374), .A2 (signal_375), .ZN (signal_1448) ) ;
    NOR2_X1 cell_366 ( .A1 (signal_1444), .A2 (signal_376), .ZN (signal_375) ) ;
    NAND2_X1 cell_367 ( .A1 (signal_377), .A2 (signal_378), .ZN (signal_376) ) ;
    NOR2_X1 cell_368 ( .A1 (signal_379), .A2 (signal_380), .ZN (signal_377) ) ;
    NAND2_X1 cell_369 ( .A1 (signal_381), .A2 (signal_382), .ZN (signal_1449) ) ;
    NOR2_X1 cell_370 ( .A1 (signal_383), .A2 (signal_384), .ZN (signal_382) ) ;
    NAND2_X1 cell_371 ( .A1 (signal_385), .A2 (signal_386), .ZN (signal_1450) ) ;
    NOR2_X1 cell_372 ( .A1 (signal_371), .A2 (signal_387), .ZN (signal_386) ) ;
    NAND2_X1 cell_373 ( .A1 (signal_388), .A2 (signal_378), .ZN (signal_387) ) ;
    NAND2_X1 cell_374 ( .A1 (signal_389), .A2 (signal_388), .ZN (signal_1451) ) ;
    NOR2_X1 cell_375 ( .A1 (signal_390), .A2 (signal_391), .ZN (signal_388) ) ;
    NAND2_X1 cell_376 ( .A1 (signal_392), .A2 (signal_393), .ZN (signal_1452) ) ;
    NOR2_X1 cell_377 ( .A1 (signal_368), .A2 (signal_394), .ZN (signal_392) ) ;
    NAND2_X1 cell_378 ( .A1 (signal_395), .A2 (signal_378), .ZN (signal_394) ) ;
    INV_X1 cell_379 ( .A (signal_396), .ZN (signal_395) ) ;
    OR2_X1 cell_380 ( .A1 (signal_368), .A2 (signal_397), .ZN (signal_1453) ) ;
    NAND2_X1 cell_381 ( .A1 (signal_381), .A2 (signal_398), .ZN (signal_397) ) ;
    NOR2_X1 cell_382 ( .A1 (signal_399), .A2 (signal_371), .ZN (signal_381) ) ;
    NAND2_X1 cell_383 ( .A1 (signal_400), .A2 (signal_373), .ZN (signal_368) ) ;
    NAND2_X1 cell_384 ( .A1 (signal_401), .A2 (signal_402), .ZN (signal_1454) ) ;
    NOR2_X1 cell_385 ( .A1 (signal_396), .A2 (signal_403), .ZN (signal_402) ) ;
    OR2_X1 cell_386 ( .A1 (signal_371), .A2 (signal_379), .ZN (signal_403) ) ;
    INV_X1 cell_387 ( .A (signal_400), .ZN (signal_379) ) ;
    NAND2_X1 cell_388 ( .A1 (signal_404), .A2 (signal_405), .ZN (signal_400) ) ;
    NAND2_X1 cell_389 ( .A1 (signal_406), .A2 (signal_407), .ZN (signal_405) ) ;
    NOR2_X1 cell_390 ( .A1 (signal_455), .A2 (signal_408), .ZN (signal_371) ) ;
    MUX2_X1 cell_391 ( .S (signal_925), .A (signal_409), .B (signal_410), .Z (signal_408) ) ;
    NAND2_X1 cell_392 ( .A1 (signal_411), .A2 (signal_412), .ZN (signal_1440) ) ;
    NOR2_X1 cell_393 ( .A1 (signal_383), .A2 (signal_396), .ZN (signal_411) ) ;
    NAND2_X1 cell_394 ( .A1 (signal_413), .A2 (signal_389), .ZN (signal_1441) ) ;
    NOR2_X1 cell_395 ( .A1 (signal_414), .A2 (signal_415), .ZN (signal_389) ) ;
    NAND2_X1 cell_396 ( .A1 (signal_367), .A2 (signal_378), .ZN (signal_415) ) ;
    OR2_X1 cell_397 ( .A1 (signal_454), .A2 (signal_416), .ZN (signal_378) ) ;
    MUX2_X1 cell_398 ( .S (signal_925), .A (signal_417), .B (signal_418), .Z (signal_416) ) ;
    NAND2_X1 cell_399 ( .A1 (signal_398), .A2 (signal_419), .ZN (signal_1442) ) ;
    NOR2_X1 cell_400 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_419) ) ;
    INV_X1 cell_401 ( .A (signal_413), .ZN (signal_421) ) ;
    NOR2_X1 cell_402 ( .A1 (signal_422), .A2 (signal_391), .ZN (signal_398) ) ;
    NAND2_X1 cell_403 ( .A1 (signal_423), .A2 (signal_393), .ZN (signal_1443) ) ;
    INV_X1 cell_404 ( .A (signal_399), .ZN (signal_393) ) ;
    NOR2_X1 cell_405 ( .A1 (signal_380), .A2 (signal_424), .ZN (signal_423) ) ;
    NAND2_X1 cell_406 ( .A1 (signal_372), .A2 (signal_413), .ZN (signal_424) ) ;
    NOR2_X1 cell_407 ( .A1 (signal_390), .A2 (signal_414), .ZN (signal_372) ) ;
    NAND2_X1 cell_408 ( .A1 (signal_385), .A2 (signal_425), .ZN (signal_414) ) ;
    NAND2_X1 cell_409 ( .A1 (signal_454), .A2 (signal_426), .ZN (signal_425) ) ;
    NAND2_X1 cell_410 ( .A1 (signal_418), .A2 (signal_406), .ZN (signal_426) ) ;
    NOR2_X1 cell_411 ( .A1 (signal_383), .A2 (signal_427), .ZN (signal_385) ) ;
    NOR2_X1 cell_412 ( .A1 (signal_455), .A2 (signal_428), .ZN (signal_427) ) ;
    MUX2_X1 cell_413 ( .S (signal_925), .A (signal_407), .B (signal_417), .Z (signal_428) ) ;
    NOR2_X1 cell_414 ( .A1 (signal_454), .A2 (signal_429), .ZN (signal_383) ) ;
    MUX2_X1 cell_415 ( .S (signal_925), .A (signal_409), .B (signal_430), .Z (signal_429) ) ;
    OR2_X1 cell_416 ( .A1 (signal_384), .A2 (signal_370), .ZN (signal_1444) ) ;
    NAND2_X1 cell_417 ( .A1 (signal_413), .A2 (signal_373), .ZN (signal_384) ) ;
    NAND2_X1 cell_418 ( .A1 (signal_431), .A2 (signal_432), .ZN (signal_373) ) ;
    AND2_X1 cell_419 ( .A1 (signal_455), .A2 (signal_925), .ZN (signal_432) ) ;
    NOR2_X1 cell_420 ( .A1 (signal_433), .A2 (signal_396), .ZN (signal_413) ) ;
    NOR2_X1 cell_421 ( .A1 (signal_454), .A2 (signal_434), .ZN (signal_396) ) ;
    MUX2_X1 cell_422 ( .S (signal_925), .A (signal_418), .B (signal_417), .Z (signal_434) ) ;
    NOR2_X1 cell_423 ( .A1 (signal_454), .A2 (signal_435), .ZN (signal_433) ) ;
    MUX2_X1 cell_424 ( .S (signal_925), .A (signal_430), .B (signal_409), .Z (signal_435) ) ;
    NAND2_X1 cell_425 ( .A1 (signal_436), .A2 (signal_412), .ZN (signal_1445) ) ;
    NOR2_X1 cell_426 ( .A1 (signal_437), .A2 (signal_370), .ZN (signal_412) ) ;
    NOR2_X1 cell_427 ( .A1 (signal_455), .A2 (signal_438), .ZN (signal_370) ) ;
    MUX2_X1 cell_428 ( .S (signal_925), .A (signal_418), .B (signal_406), .Z (signal_438) ) ;
    INV_X1 cell_429 ( .A (signal_439), .ZN (signal_437) ) ;
    INV_X1 cell_430 ( .A (signal_390), .ZN (signal_436) ) ;
    NAND2_X1 cell_431 ( .A1 (signal_401), .A2 (signal_439), .ZN (signal_1455) ) ;
    NOR2_X1 cell_432 ( .A1 (signal_380), .A2 (signal_391), .ZN (signal_439) ) ;
    NOR2_X1 cell_433 ( .A1 (signal_455), .A2 (signal_440), .ZN (signal_391) ) ;
    MUX2_X1 cell_434 ( .S (signal_925), .A (signal_410), .B (signal_409), .Z (signal_440) ) ;
    NAND2_X1 cell_435 ( .A1 (signal_441), .A2 (signal_442), .ZN (signal_409) ) ;
    NAND2_X1 cell_436 ( .A1 (signal_443), .A2 (signal_926), .ZN (signal_410) ) ;
    NOR2_X1 cell_437 ( .A1 (signal_455), .A2 (signal_444), .ZN (signal_380) ) ;
    MUX2_X1 cell_438 ( .S (signal_925), .A (signal_417), .B (signal_407), .Z (signal_444) ) ;
    NAND2_X1 cell_439 ( .A1 (enc_dec), .A2 (signal_431), .ZN (signal_407) ) ;
    NOR2_X1 cell_440 ( .A1 (signal_924), .A2 (signal_442), .ZN (signal_431) ) ;
    NAND2_X1 cell_441 ( .A1 (signal_445), .A2 (signal_442), .ZN (signal_417) ) ;
    NOR2_X1 cell_442 ( .A1 (signal_399), .A2 (signal_446), .ZN (signal_401) ) ;
    NAND2_X1 cell_443 ( .A1 (signal_374), .A2 (signal_367), .ZN (signal_446) ) ;
    NAND2_X1 cell_444 ( .A1 (signal_420), .A2 (signal_447), .ZN (signal_367) ) ;
    OR2_X1 cell_445 ( .A1 (signal_443), .A2 (signal_441), .ZN (signal_447) ) ;
    AND2_X1 cell_446 ( .A1 (signal_926), .A2 (signal_404), .ZN (signal_420) ) ;
    NOR2_X1 cell_447 ( .A1 (signal_454), .A2 (signal_925), .ZN (signal_404) ) ;
    NOR2_X1 cell_448 ( .A1 (signal_390), .A2 (signal_422), .ZN (signal_374) ) ;
    NOR2_X1 cell_449 ( .A1 (signal_455), .A2 (signal_448), .ZN (signal_422) ) ;
    MUX2_X1 cell_450 ( .S (signal_925), .A (signal_406), .B (signal_418), .Z (signal_448) ) ;
    NAND2_X1 cell_451 ( .A1 (enc_dec), .A2 (signal_449), .ZN (signal_418) ) ;
    NOR2_X1 cell_452 ( .A1 (signal_924), .A2 (signal_926), .ZN (signal_449) ) ;
    NAND2_X1 cell_453 ( .A1 (signal_926), .A2 (signal_445), .ZN (signal_406) ) ;
    NOR2_X1 cell_454 ( .A1 (enc_dec), .A2 (signal_450), .ZN (signal_445) ) ;
    INV_X1 cell_455 ( .A (signal_924), .ZN (signal_450) ) ;
    NOR2_X1 cell_456 ( .A1 (signal_455), .A2 (signal_451), .ZN (signal_390) ) ;
    MUX2_X1 cell_457 ( .S (signal_925), .A (signal_430), .B (signal_452), .Z (signal_451) ) ;
    NOR2_X1 cell_458 ( .A1 (signal_455), .A2 (signal_453), .ZN (signal_399) ) ;
    MUX2_X1 cell_459 ( .S (signal_925), .A (signal_452), .B (signal_430), .Z (signal_453) ) ;
    NAND2_X1 cell_460 ( .A1 (signal_443), .A2 (signal_442), .ZN (signal_430) ) ;
    INV_X1 cell_461 ( .A (signal_926), .ZN (signal_442) ) ;
    NOR2_X1 cell_462 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_443) ) ;
    NAND2_X1 cell_463 ( .A1 (signal_441), .A2 (signal_926), .ZN (signal_452) ) ;
    AND2_X1 cell_464 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_441) ) ;
    INV_X1 cell_465 ( .A (signal_454), .ZN (signal_455) ) ;
    INV_X1 cell_466 ( .A (signal_927), .ZN (signal_454) ) ;
    INV_X1 cell_467 ( .A (signal_927), .ZN (signal_456) ) ;
    INV_X1 cell_468 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_469 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_470 ( .A (signal_456), .ZN (signal_457) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_471 ( .s (signal_927), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_2144, signal_302}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_472 ( .s (signal_927), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_2145, signal_303}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_473 ( .s (signal_927), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_2146, signal_304}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_474 ( .s (signal_927), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_2147, signal_305}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_475 ( .s (signal_927), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_2148, signal_306}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_476 ( .s (signal_459), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_2541, signal_307}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_477 ( .s (signal_457), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_2542, signal_308}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_478 ( .s (signal_458), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_2543, signal_309}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_479 ( .s (signal_927), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_2149, signal_310}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_480 ( .s (signal_927), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_2150, signal_311}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_481 ( .s (signal_927), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_2151, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_482 ( .s (signal_927), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_2152, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_483 ( .s (signal_458), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_2544, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_484 ( .s (signal_927), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_2153, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_485 ( .s (signal_927), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_2154, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_486 ( .s (signal_927), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_2155, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_487 ( .s (signal_457), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_2545, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_488 ( .s (signal_459), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_2546, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_489 ( .s (signal_457), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_2547, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_490 ( .s (signal_457), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_2548, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_491 ( .s (signal_457), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_2549, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_492 ( .s (signal_457), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_2550, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_493 ( .s (signal_458), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_2551, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_494 ( .s (signal_459), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_2552, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_495 ( .s (signal_457), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_2553, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_496 ( .s (signal_458), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_2554, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_497 ( .s (signal_927), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_2156, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_498 ( .s (signal_457), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_2555, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_499 ( .s (signal_457), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_2556, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_500 ( .s (signal_457), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_2557, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_501 ( .s (signal_457), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_2558, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_502 ( .s (signal_457), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_2559, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_503 ( .s (signal_457), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_2560, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_504 ( .s (signal_457), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_2561, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_505 ( .s (signal_457), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_2562, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_506 ( .s (signal_457), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_2563, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_507 ( .s (signal_457), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_2564, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_508 ( .s (signal_457), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_2565, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_509 ( .s (signal_457), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_2566, signal_340}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_510 ( .s (signal_457), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_2567, signal_341}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_511 ( .s (signal_458), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_2568, signal_342}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_512 ( .s (signal_458), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_2569, signal_343}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_513 ( .s (signal_458), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_2570, signal_344}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_514 ( .s (signal_458), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_2571, signal_345}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_515 ( .s (signal_458), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_2572, signal_346}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_516 ( .s (signal_458), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_2573, signal_347}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_517 ( .s (signal_458), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_2574, signal_348}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_518 ( .s (signal_458), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_2575, signal_349}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_519 ( .s (signal_458), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_2576, signal_350}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_520 ( .s (signal_458), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_2577, signal_351}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_521 ( .s (signal_458), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_2578, signal_352}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_522 ( .s (signal_458), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_2579, signal_353}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_523 ( .s (signal_459), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_2580, signal_354}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_524 ( .s (signal_459), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_2581, signal_355}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_525 ( .s (signal_459), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_2582, signal_356}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_526 ( .s (signal_459), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_2583, signal_357}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_527 ( .s (signal_459), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_2584, signal_358}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_528 ( .s (signal_459), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_2585, signal_359}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_529 ( .s (signal_459), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_2586, signal_360}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_530 ( .s (signal_459), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_2587, signal_361}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_531 ( .s (signal_459), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_2588, signal_362}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_532 ( .s (signal_459), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_2589, signal_363}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_533 ( .s (signal_459), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_2590, signal_364}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_534 ( .s (signal_459), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_2591, signal_365}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1255 ( .a ({signal_2157, signal_1312}), .b ({signal_2158, signal_1456}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1256 ( .a ({signal_2159, signal_1313}), .b ({signal_2160, signal_1457}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1257 ( .a ({signal_2161, signal_1314}), .b ({signal_2162, signal_1458}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1258 ( .a ({signal_2163, signal_1315}), .b ({signal_2164, signal_1459}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1259 ( .a ({signal_2165, signal_1316}), .b ({signal_2166, signal_1460}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1260 ( .a ({signal_2167, signal_1317}), .b ({signal_2168, signal_1461}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1261 ( .a ({signal_2169, signal_1318}), .b ({signal_2170, signal_1462}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1262 ( .a ({signal_2171, signal_1319}), .b ({signal_2172, signal_1463}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1263 ( .a ({signal_2173, signal_1320}), .b ({signal_2174, signal_1464}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1264 ( .a ({signal_2175, signal_1321}), .b ({signal_2176, signal_1465}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1265 ( .a ({signal_2177, signal_1322}), .b ({signal_2178, signal_1466}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1266 ( .a ({signal_2179, signal_1323}), .b ({signal_2180, signal_1467}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1267 ( .a ({signal_2181, signal_1324}), .b ({signal_2182, signal_1468}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1268 ( .a ({signal_2183, signal_1325}), .b ({signal_2184, signal_1469}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1269 ( .a ({signal_2185, signal_1326}), .b ({signal_2186, signal_1470}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1270 ( .a ({signal_2187, signal_1327}), .b ({signal_2188, signal_1471}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1271 ( .a ({signal_2189, signal_1328}), .b ({signal_2190, signal_1472}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1272 ( .a ({signal_2191, signal_1329}), .b ({signal_2192, signal_1473}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1273 ( .a ({signal_2193, signal_1330}), .b ({signal_2194, signal_1474}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1274 ( .a ({signal_2195, signal_1331}), .b ({signal_2196, signal_1475}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1275 ( .a ({signal_2197, signal_1332}), .b ({signal_2198, signal_1476}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1276 ( .a ({signal_2199, signal_1333}), .b ({signal_2200, signal_1477}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1277 ( .a ({signal_2201, signal_1334}), .b ({signal_2202, signal_1478}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1278 ( .a ({signal_2203, signal_1335}), .b ({signal_2204, signal_1479}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1279 ( .a ({signal_2205, signal_1336}), .b ({signal_2206, signal_1480}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1280 ( .a ({signal_2207, signal_1337}), .b ({signal_2208, signal_1481}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1281 ( .a ({signal_2209, signal_1338}), .b ({signal_2210, signal_1482}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1282 ( .a ({signal_2211, signal_1339}), .b ({signal_2212, signal_1483}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1283 ( .a ({signal_2213, signal_1340}), .b ({signal_2214, signal_1484}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1284 ( .a ({signal_2215, signal_1341}), .b ({signal_2216, signal_1485}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1285 ( .a ({signal_2217, signal_1342}), .b ({signal_2218, signal_1486}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1286 ( .a ({signal_2219, signal_1343}), .b ({signal_2220, signal_1487}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1287 ( .a ({signal_2221, signal_1344}), .b ({signal_2222, signal_1488}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1288 ( .a ({signal_2223, signal_1345}), .b ({signal_2224, signal_1489}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1289 ( .a ({signal_2225, signal_1346}), .b ({signal_2226, signal_1490}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1290 ( .a ({signal_2227, signal_1347}), .b ({signal_2228, signal_1491}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1291 ( .a ({signal_2229, signal_1348}), .b ({signal_2230, signal_1492}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1292 ( .a ({signal_2231, signal_1349}), .b ({signal_2232, signal_1493}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1293 ( .a ({signal_2233, signal_1350}), .b ({signal_2234, signal_1494}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1294 ( .a ({signal_2235, signal_1351}), .b ({signal_2236, signal_1495}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1295 ( .a ({signal_2237, signal_1352}), .b ({signal_2238, signal_1496}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1296 ( .a ({signal_2239, signal_1353}), .b ({signal_2240, signal_1497}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1297 ( .a ({signal_2241, signal_1354}), .b ({signal_2242, signal_1498}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1298 ( .a ({signal_2243, signal_1355}), .b ({signal_2244, signal_1499}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1299 ( .a ({signal_2245, signal_1356}), .b ({signal_2246, signal_1500}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1300 ( .a ({signal_2247, signal_1357}), .b ({signal_2248, signal_1501}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1301 ( .a ({signal_2249, signal_1358}), .b ({signal_2250, signal_1502}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1302 ( .a ({signal_2251, signal_1359}), .b ({signal_2252, signal_1503}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1303 ( .a ({signal_2253, signal_1360}), .b ({signal_2254, signal_1504}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1304 ( .a ({signal_2255, signal_1361}), .b ({signal_2256, signal_1505}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1305 ( .a ({signal_2257, signal_1362}), .b ({signal_2258, signal_1506}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1306 ( .a ({signal_2259, signal_1363}), .b ({signal_2260, signal_1507}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1307 ( .a ({signal_2261, signal_1364}), .b ({signal_2262, signal_1508}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1308 ( .a ({signal_2263, signal_1365}), .b ({signal_2264, signal_1509}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1309 ( .a ({signal_2265, signal_1366}), .b ({signal_2266, signal_1510}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1310 ( .a ({signal_2267, signal_1367}), .b ({signal_2268, signal_1511}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1311 ( .a ({signal_2269, signal_1368}), .b ({signal_2270, signal_1512}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1312 ( .a ({signal_2271, signal_1369}), .b ({signal_2272, signal_1513}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1313 ( .a ({signal_2273, signal_1370}), .b ({signal_2274, signal_1514}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1314 ( .a ({signal_2275, signal_1371}), .b ({signal_2276, signal_1515}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1315 ( .a ({signal_2277, signal_1372}), .b ({signal_2278, signal_1516}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1316 ( .a ({signal_2279, signal_1373}), .b ({signal_2280, signal_1517}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1317 ( .a ({signal_2281, signal_1374}), .b ({signal_2282, signal_1518}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1318 ( .a ({signal_2283, signal_1375}), .b ({signal_2284, signal_1519}) ) ;
    ClockGatingController #(9) cell_1815 ( .clk (clk), .rst (reset), .GatedClk (signal_3712), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .a ({signal_2277, signal_1372}), .b ({signal_2283, signal_1375}), .clk (clk), .r (Fresh[0]), .c ({signal_2285, signal_1520}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .a ({signal_2269, signal_1368}), .b ({signal_2275, signal_1371}), .clk (clk), .r (Fresh[1]), .c ({signal_2286, signal_1521}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .a ({signal_2261, signal_1364}), .b ({signal_2267, signal_1367}), .clk (clk), .r (Fresh[2]), .c ({signal_2287, signal_1522}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .a ({signal_2253, signal_1360}), .b ({signal_2259, signal_1363}), .clk (clk), .r (Fresh[3]), .c ({signal_2288, signal_1523}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .a ({signal_2245, signal_1356}), .b ({signal_2251, signal_1359}), .clk (clk), .r (Fresh[4]), .c ({signal_2289, signal_1524}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .a ({signal_2237, signal_1352}), .b ({signal_2243, signal_1355}), .clk (clk), .r (Fresh[5]), .c ({signal_2290, signal_1525}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .a ({signal_2229, signal_1348}), .b ({signal_2235, signal_1351}), .clk (clk), .r (Fresh[6]), .c ({signal_2291, signal_1526}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .a ({signal_2221, signal_1344}), .b ({signal_2227, signal_1347}), .clk (clk), .r (Fresh[7]), .c ({signal_2292, signal_1527}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .a ({signal_2213, signal_1340}), .b ({signal_2219, signal_1343}), .clk (clk), .r (Fresh[8]), .c ({signal_2293, signal_1528}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .a ({signal_2205, signal_1336}), .b ({signal_2211, signal_1339}), .clk (clk), .r (Fresh[9]), .c ({signal_2294, signal_1529}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .a ({signal_2197, signal_1332}), .b ({signal_2203, signal_1335}), .clk (clk), .r (Fresh[10]), .c ({signal_2295, signal_1530}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .a ({signal_2189, signal_1328}), .b ({signal_2195, signal_1331}), .clk (clk), .r (Fresh[11]), .c ({signal_2296, signal_1531}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .a ({signal_2181, signal_1324}), .b ({signal_2187, signal_1327}), .clk (clk), .r (Fresh[12]), .c ({signal_2297, signal_1532}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .a ({signal_2173, signal_1320}), .b ({signal_2179, signal_1323}), .clk (clk), .r (Fresh[13]), .c ({signal_2298, signal_1533}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .a ({signal_2165, signal_1316}), .b ({signal_2171, signal_1319}), .clk (clk), .r (Fresh[14]), .c ({signal_2299, signal_1534}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .a ({signal_2157, signal_1312}), .b ({signal_2163, signal_1315}), .clk (clk), .r (Fresh[15]), .c ({signal_2300, signal_1535}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .a ({signal_2277, signal_1372}), .b ({signal_2279, signal_1373}), .clk (clk), .r (Fresh[16]), .c ({signal_2301, signal_1536}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .a ({signal_2269, signal_1368}), .b ({signal_2271, signal_1369}), .clk (clk), .r (Fresh[17]), .c ({signal_2302, signal_1537}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .a ({signal_2261, signal_1364}), .b ({signal_2263, signal_1365}), .clk (clk), .r (Fresh[18]), .c ({signal_2303, signal_1538}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .a ({signal_2253, signal_1360}), .b ({signal_2255, signal_1361}), .clk (clk), .r (Fresh[19]), .c ({signal_2304, signal_1539}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .a ({signal_2245, signal_1356}), .b ({signal_2247, signal_1357}), .clk (clk), .r (Fresh[20]), .c ({signal_2305, signal_1540}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .a ({signal_2237, signal_1352}), .b ({signal_2239, signal_1353}), .clk (clk), .r (Fresh[21]), .c ({signal_2306, signal_1541}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .a ({signal_2229, signal_1348}), .b ({signal_2231, signal_1349}), .clk (clk), .r (Fresh[22]), .c ({signal_2307, signal_1542}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .a ({signal_2221, signal_1344}), .b ({signal_2223, signal_1345}), .clk (clk), .r (Fresh[23]), .c ({signal_2308, signal_1543}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .a ({signal_2213, signal_1340}), .b ({signal_2215, signal_1341}), .clk (clk), .r (Fresh[24]), .c ({signal_2309, signal_1544}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .a ({signal_2205, signal_1336}), .b ({signal_2207, signal_1337}), .clk (clk), .r (Fresh[25]), .c ({signal_2310, signal_1545}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .a ({signal_2197, signal_1332}), .b ({signal_2199, signal_1333}), .clk (clk), .r (Fresh[26]), .c ({signal_2311, signal_1546}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .a ({signal_2189, signal_1328}), .b ({signal_2191, signal_1329}), .clk (clk), .r (Fresh[27]), .c ({signal_2312, signal_1547}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1347 ( .a ({signal_2181, signal_1324}), .b ({signal_2183, signal_1325}), .clk (clk), .r (Fresh[28]), .c ({signal_2313, signal_1548}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1348 ( .a ({signal_2173, signal_1320}), .b ({signal_2175, signal_1321}), .clk (clk), .r (Fresh[29]), .c ({signal_2314, signal_1549}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1349 ( .a ({signal_2165, signal_1316}), .b ({signal_2167, signal_1317}), .clk (clk), .r (Fresh[30]), .c ({signal_2315, signal_1550}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1350 ( .a ({signal_2157, signal_1312}), .b ({signal_2159, signal_1313}), .clk (clk), .r (Fresh[31]), .c ({signal_2316, signal_1551}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1351 ( .a ({signal_2285, signal_1520}), .b ({signal_2445, signal_1552}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1352 ( .a ({signal_2286, signal_1521}), .b ({signal_2446, signal_1553}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1353 ( .a ({signal_2287, signal_1522}), .b ({signal_2447, signal_1554}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1354 ( .a ({signal_2288, signal_1523}), .b ({signal_2448, signal_1555}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1355 ( .a ({signal_2289, signal_1524}), .b ({signal_2449, signal_1556}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1356 ( .a ({signal_2290, signal_1525}), .b ({signal_2450, signal_1557}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1357 ( .a ({signal_2291, signal_1526}), .b ({signal_2451, signal_1558}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1358 ( .a ({signal_2292, signal_1527}), .b ({signal_2452, signal_1559}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1359 ( .a ({signal_2293, signal_1528}), .b ({signal_2453, signal_1560}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1360 ( .a ({signal_2294, signal_1529}), .b ({signal_2454, signal_1561}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1361 ( .a ({signal_2295, signal_1530}), .b ({signal_2455, signal_1562}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1362 ( .a ({signal_2296, signal_1531}), .b ({signal_2456, signal_1563}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1363 ( .a ({signal_2297, signal_1532}), .b ({signal_2457, signal_1564}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1364 ( .a ({signal_2298, signal_1533}), .b ({signal_2458, signal_1565}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1365 ( .a ({signal_2299, signal_1534}), .b ({signal_2459, signal_1566}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1366 ( .a ({signal_2300, signal_1535}), .b ({signal_2460, signal_1567}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1367 ( .a ({signal_2301, signal_1536}), .b ({signal_2461, signal_1568}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1368 ( .a ({signal_2302, signal_1537}), .b ({signal_2462, signal_1569}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1369 ( .a ({signal_2303, signal_1538}), .b ({signal_2463, signal_1570}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1370 ( .a ({signal_2304, signal_1539}), .b ({signal_2464, signal_1571}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1371 ( .a ({signal_2305, signal_1540}), .b ({signal_2465, signal_1572}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1372 ( .a ({signal_2306, signal_1541}), .b ({signal_2466, signal_1573}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1373 ( .a ({signal_2307, signal_1542}), .b ({signal_2467, signal_1574}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1374 ( .a ({signal_2308, signal_1543}), .b ({signal_2468, signal_1575}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1375 ( .a ({signal_2309, signal_1544}), .b ({signal_2469, signal_1576}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1376 ( .a ({signal_2310, signal_1545}), .b ({signal_2470, signal_1577}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1377 ( .a ({signal_2311, signal_1546}), .b ({signal_2471, signal_1578}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1378 ( .a ({signal_2312, signal_1547}), .b ({signal_2472, signal_1579}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1379 ( .a ({signal_2313, signal_1548}), .b ({signal_2473, signal_1580}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1380 ( .a ({signal_2314, signal_1549}), .b ({signal_2474, signal_1581}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1381 ( .a ({signal_2315, signal_1550}), .b ({signal_2475, signal_1582}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1382 ( .a ({signal_2316, signal_1551}), .b ({signal_2476, signal_1583}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1383 ( .a ({signal_2278, signal_1516}), .b ({signal_2280, signal_1517}), .clk (clk), .r (Fresh[32]), .c ({signal_2477, signal_1584}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .a ({signal_2270, signal_1512}), .b ({signal_2272, signal_1513}), .clk (clk), .r (Fresh[33]), .c ({signal_2478, signal_1585}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .a ({signal_2262, signal_1508}), .b ({signal_2264, signal_1509}), .clk (clk), .r (Fresh[34]), .c ({signal_2479, signal_1586}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .a ({signal_2254, signal_1504}), .b ({signal_2256, signal_1505}), .clk (clk), .r (Fresh[35]), .c ({signal_2480, signal_1587}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .a ({signal_2246, signal_1500}), .b ({signal_2248, signal_1501}), .clk (clk), .r (Fresh[36]), .c ({signal_2481, signal_1588}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .a ({signal_2238, signal_1496}), .b ({signal_2240, signal_1497}), .clk (clk), .r (Fresh[37]), .c ({signal_2482, signal_1589}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .a ({signal_2230, signal_1492}), .b ({signal_2232, signal_1493}), .clk (clk), .r (Fresh[38]), .c ({signal_2483, signal_1590}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .a ({signal_2222, signal_1488}), .b ({signal_2224, signal_1489}), .clk (clk), .r (Fresh[39]), .c ({signal_2484, signal_1591}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .a ({signal_2214, signal_1484}), .b ({signal_2216, signal_1485}), .clk (clk), .r (Fresh[40]), .c ({signal_2485, signal_1592}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .a ({signal_2206, signal_1480}), .b ({signal_2208, signal_1481}), .clk (clk), .r (Fresh[41]), .c ({signal_2486, signal_1593}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .a ({signal_2198, signal_1476}), .b ({signal_2200, signal_1477}), .clk (clk), .r (Fresh[42]), .c ({signal_2487, signal_1594}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .a ({signal_2190, signal_1472}), .b ({signal_2192, signal_1473}), .clk (clk), .r (Fresh[43]), .c ({signal_2488, signal_1595}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .a ({signal_2182, signal_1468}), .b ({signal_2184, signal_1469}), .clk (clk), .r (Fresh[44]), .c ({signal_2489, signal_1596}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .a ({signal_2174, signal_1464}), .b ({signal_2176, signal_1465}), .clk (clk), .r (Fresh[45]), .c ({signal_2490, signal_1597}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .a ({signal_2166, signal_1460}), .b ({signal_2168, signal_1461}), .clk (clk), .r (Fresh[46]), .c ({signal_2491, signal_1598}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1398 ( .a ({signal_2158, signal_1456}), .b ({signal_2160, signal_1457}), .clk (clk), .r (Fresh[47]), .c ({signal_2492, signal_1599}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1399 ( .a ({signal_2278, signal_1516}), .b ({signal_2284, signal_1519}), .clk (clk), .r (Fresh[48]), .c ({signal_2493, signal_1600}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1400 ( .a ({signal_2277, signal_1372}), .b ({signal_2280, signal_1517}), .clk (clk), .r (Fresh[49]), .c ({signal_2494, signal_1601}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1401 ( .a ({signal_2278, signal_1516}), .b ({signal_2279, signal_1373}), .clk (clk), .r (Fresh[50]), .c ({signal_2495, signal_1602}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1402 ( .a ({signal_2270, signal_1512}), .b ({signal_2276, signal_1515}), .clk (clk), .r (Fresh[51]), .c ({signal_2496, signal_1603}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1403 ( .a ({signal_2269, signal_1368}), .b ({signal_2272, signal_1513}), .clk (clk), .r (Fresh[52]), .c ({signal_2497, signal_1604}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1404 ( .a ({signal_2270, signal_1512}), .b ({signal_2271, signal_1369}), .clk (clk), .r (Fresh[53]), .c ({signal_2498, signal_1605}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1405 ( .a ({signal_2262, signal_1508}), .b ({signal_2268, signal_1511}), .clk (clk), .r (Fresh[54]), .c ({signal_2499, signal_1606}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1406 ( .a ({signal_2261, signal_1364}), .b ({signal_2264, signal_1509}), .clk (clk), .r (Fresh[55]), .c ({signal_2500, signal_1607}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1407 ( .a ({signal_2262, signal_1508}), .b ({signal_2263, signal_1365}), .clk (clk), .r (Fresh[56]), .c ({signal_2501, signal_1608}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1408 ( .a ({signal_2254, signal_1504}), .b ({signal_2260, signal_1507}), .clk (clk), .r (Fresh[57]), .c ({signal_2502, signal_1609}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1409 ( .a ({signal_2253, signal_1360}), .b ({signal_2256, signal_1505}), .clk (clk), .r (Fresh[58]), .c ({signal_2503, signal_1610}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1410 ( .a ({signal_2254, signal_1504}), .b ({signal_2255, signal_1361}), .clk (clk), .r (Fresh[59]), .c ({signal_2504, signal_1611}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1411 ( .a ({signal_2246, signal_1500}), .b ({signal_2252, signal_1503}), .clk (clk), .r (Fresh[60]), .c ({signal_2505, signal_1612}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1412 ( .a ({signal_2245, signal_1356}), .b ({signal_2248, signal_1501}), .clk (clk), .r (Fresh[61]), .c ({signal_2506, signal_1613}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1413 ( .a ({signal_2246, signal_1500}), .b ({signal_2247, signal_1357}), .clk (clk), .r (Fresh[62]), .c ({signal_2507, signal_1614}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1414 ( .a ({signal_2238, signal_1496}), .b ({signal_2244, signal_1499}), .clk (clk), .r (Fresh[63]), .c ({signal_2508, signal_1615}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1415 ( .a ({signal_2237, signal_1352}), .b ({signal_2240, signal_1497}), .clk (clk), .r (Fresh[64]), .c ({signal_2509, signal_1616}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .a ({signal_2238, signal_1496}), .b ({signal_2239, signal_1353}), .clk (clk), .r (Fresh[65]), .c ({signal_2510, signal_1617}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .a ({signal_2230, signal_1492}), .b ({signal_2236, signal_1495}), .clk (clk), .r (Fresh[66]), .c ({signal_2511, signal_1618}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .a ({signal_2229, signal_1348}), .b ({signal_2232, signal_1493}), .clk (clk), .r (Fresh[67]), .c ({signal_2512, signal_1619}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .a ({signal_2230, signal_1492}), .b ({signal_2231, signal_1349}), .clk (clk), .r (Fresh[68]), .c ({signal_2513, signal_1620}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .a ({signal_2222, signal_1488}), .b ({signal_2228, signal_1491}), .clk (clk), .r (Fresh[69]), .c ({signal_2514, signal_1621}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .a ({signal_2221, signal_1344}), .b ({signal_2224, signal_1489}), .clk (clk), .r (Fresh[70]), .c ({signal_2515, signal_1622}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .a ({signal_2222, signal_1488}), .b ({signal_2223, signal_1345}), .clk (clk), .r (Fresh[71]), .c ({signal_2516, signal_1623}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .a ({signal_2214, signal_1484}), .b ({signal_2220, signal_1487}), .clk (clk), .r (Fresh[72]), .c ({signal_2517, signal_1624}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .a ({signal_2213, signal_1340}), .b ({signal_2216, signal_1485}), .clk (clk), .r (Fresh[73]), .c ({signal_2518, signal_1625}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .a ({signal_2214, signal_1484}), .b ({signal_2215, signal_1341}), .clk (clk), .r (Fresh[74]), .c ({signal_2519, signal_1626}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .a ({signal_2206, signal_1480}), .b ({signal_2212, signal_1483}), .clk (clk), .r (Fresh[75]), .c ({signal_2520, signal_1627}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .a ({signal_2205, signal_1336}), .b ({signal_2208, signal_1481}), .clk (clk), .r (Fresh[76]), .c ({signal_2521, signal_1628}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .a ({signal_2206, signal_1480}), .b ({signal_2207, signal_1337}), .clk (clk), .r (Fresh[77]), .c ({signal_2522, signal_1629}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .a ({signal_2198, signal_1476}), .b ({signal_2204, signal_1479}), .clk (clk), .r (Fresh[78]), .c ({signal_2523, signal_1630}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .a ({signal_2197, signal_1332}), .b ({signal_2200, signal_1477}), .clk (clk), .r (Fresh[79]), .c ({signal_2524, signal_1631}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .a ({signal_2198, signal_1476}), .b ({signal_2199, signal_1333}), .clk (clk), .r (Fresh[80]), .c ({signal_2525, signal_1632}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .a ({signal_2190, signal_1472}), .b ({signal_2196, signal_1475}), .clk (clk), .r (Fresh[81]), .c ({signal_2526, signal_1633}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .a ({signal_2189, signal_1328}), .b ({signal_2192, signal_1473}), .clk (clk), .r (Fresh[82]), .c ({signal_2527, signal_1634}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .a ({signal_2190, signal_1472}), .b ({signal_2191, signal_1329}), .clk (clk), .r (Fresh[83]), .c ({signal_2528, signal_1635}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .a ({signal_2182, signal_1468}), .b ({signal_2188, signal_1471}), .clk (clk), .r (Fresh[84]), .c ({signal_2529, signal_1636}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .a ({signal_2181, signal_1324}), .b ({signal_2184, signal_1469}), .clk (clk), .r (Fresh[85]), .c ({signal_2530, signal_1637}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .a ({signal_2182, signal_1468}), .b ({signal_2183, signal_1325}), .clk (clk), .r (Fresh[86]), .c ({signal_2531, signal_1638}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .a ({signal_2174, signal_1464}), .b ({signal_2180, signal_1467}), .clk (clk), .r (Fresh[87]), .c ({signal_2532, signal_1639}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .a ({signal_2173, signal_1320}), .b ({signal_2176, signal_1465}), .clk (clk), .r (Fresh[88]), .c ({signal_2533, signal_1640}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .a ({signal_2174, signal_1464}), .b ({signal_2175, signal_1321}), .clk (clk), .r (Fresh[89]), .c ({signal_2534, signal_1641}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .a ({signal_2166, signal_1460}), .b ({signal_2172, signal_1463}), .clk (clk), .r (Fresh[90]), .c ({signal_2535, signal_1642}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .a ({signal_2165, signal_1316}), .b ({signal_2168, signal_1461}), .clk (clk), .r (Fresh[91]), .c ({signal_2536, signal_1643}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .a ({signal_2166, signal_1460}), .b ({signal_2167, signal_1317}), .clk (clk), .r (Fresh[92]), .c ({signal_2537, signal_1644}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .a ({signal_2158, signal_1456}), .b ({signal_2164, signal_1459}), .clk (clk), .r (Fresh[93]), .c ({signal_2538, signal_1645}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .a ({signal_2157, signal_1312}), .b ({signal_2160, signal_1457}), .clk (clk), .r (Fresh[94]), .c ({signal_2539, signal_1646}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .a ({signal_2158, signal_1456}), .b ({signal_2159, signal_1313}), .clk (clk), .r (Fresh[95]), .c ({signal_2540, signal_1647}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1447 ( .a ({signal_2477, signal_1584}), .b ({signal_2592, signal_1648}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1448 ( .a ({signal_2478, signal_1585}), .b ({signal_2593, signal_1649}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1449 ( .a ({signal_2479, signal_1586}), .b ({signal_2594, signal_1650}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1450 ( .a ({signal_2480, signal_1587}), .b ({signal_2595, signal_1651}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1451 ( .a ({signal_2481, signal_1588}), .b ({signal_2596, signal_1652}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1452 ( .a ({signal_2482, signal_1589}), .b ({signal_2597, signal_1653}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1453 ( .a ({signal_2483, signal_1590}), .b ({signal_2598, signal_1654}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1454 ( .a ({signal_2484, signal_1591}), .b ({signal_2599, signal_1655}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1455 ( .a ({signal_2485, signal_1592}), .b ({signal_2600, signal_1656}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1456 ( .a ({signal_2486, signal_1593}), .b ({signal_2601, signal_1657}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1457 ( .a ({signal_2487, signal_1594}), .b ({signal_2602, signal_1658}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1458 ( .a ({signal_2488, signal_1595}), .b ({signal_2603, signal_1659}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1459 ( .a ({signal_2489, signal_1596}), .b ({signal_2604, signal_1660}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1460 ( .a ({signal_2490, signal_1597}), .b ({signal_2605, signal_1661}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1461 ( .a ({signal_2491, signal_1598}), .b ({signal_2606, signal_1662}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1462 ( .a ({signal_2492, signal_1599}), .b ({signal_2607, signal_1663}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1463 ( .a ({signal_2493, signal_1600}), .b ({signal_2608, signal_1664}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1464 ( .a ({signal_2494, signal_1601}), .b ({signal_2609, signal_1665}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1465 ( .a ({signal_2495, signal_1602}), .b ({signal_2610, signal_1666}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1466 ( .a ({signal_2496, signal_1603}), .b ({signal_2611, signal_1667}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1467 ( .a ({signal_2497, signal_1604}), .b ({signal_2612, signal_1668}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1468 ( .a ({signal_2498, signal_1605}), .b ({signal_2613, signal_1669}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1469 ( .a ({signal_2499, signal_1606}), .b ({signal_2614, signal_1670}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1470 ( .a ({signal_2500, signal_1607}), .b ({signal_2615, signal_1671}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1471 ( .a ({signal_2501, signal_1608}), .b ({signal_2616, signal_1672}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1472 ( .a ({signal_2502, signal_1609}), .b ({signal_2617, signal_1673}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1473 ( .a ({signal_2503, signal_1610}), .b ({signal_2618, signal_1674}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1474 ( .a ({signal_2504, signal_1611}), .b ({signal_2619, signal_1675}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1475 ( .a ({signal_2505, signal_1612}), .b ({signal_2620, signal_1676}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1476 ( .a ({signal_2506, signal_1613}), .b ({signal_2621, signal_1677}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1477 ( .a ({signal_2507, signal_1614}), .b ({signal_2622, signal_1678}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1478 ( .a ({signal_2508, signal_1615}), .b ({signal_2623, signal_1679}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1479 ( .a ({signal_2509, signal_1616}), .b ({signal_2624, signal_1680}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1480 ( .a ({signal_2510, signal_1617}), .b ({signal_2625, signal_1681}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1481 ( .a ({signal_2511, signal_1618}), .b ({signal_2626, signal_1682}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1482 ( .a ({signal_2512, signal_1619}), .b ({signal_2627, signal_1683}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1483 ( .a ({signal_2513, signal_1620}), .b ({signal_2628, signal_1684}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1484 ( .a ({signal_2514, signal_1621}), .b ({signal_2629, signal_1685}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1485 ( .a ({signal_2515, signal_1622}), .b ({signal_2630, signal_1686}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1486 ( .a ({signal_2516, signal_1623}), .b ({signal_2631, signal_1687}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1487 ( .a ({signal_2517, signal_1624}), .b ({signal_2632, signal_1688}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1488 ( .a ({signal_2518, signal_1625}), .b ({signal_2633, signal_1689}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1489 ( .a ({signal_2519, signal_1626}), .b ({signal_2634, signal_1690}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1490 ( .a ({signal_2520, signal_1627}), .b ({signal_2635, signal_1691}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1491 ( .a ({signal_2521, signal_1628}), .b ({signal_2636, signal_1692}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1492 ( .a ({signal_2522, signal_1629}), .b ({signal_2637, signal_1693}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1493 ( .a ({signal_2523, signal_1630}), .b ({signal_2638, signal_1694}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1494 ( .a ({signal_2524, signal_1631}), .b ({signal_2639, signal_1695}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1495 ( .a ({signal_2525, signal_1632}), .b ({signal_2640, signal_1696}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1496 ( .a ({signal_2526, signal_1633}), .b ({signal_2641, signal_1697}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1497 ( .a ({signal_2527, signal_1634}), .b ({signal_2642, signal_1698}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1498 ( .a ({signal_2528, signal_1635}), .b ({signal_2643, signal_1699}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1499 ( .a ({signal_2529, signal_1636}), .b ({signal_2644, signal_1700}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1500 ( .a ({signal_2530, signal_1637}), .b ({signal_2645, signal_1701}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1501 ( .a ({signal_2531, signal_1638}), .b ({signal_2646, signal_1702}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1502 ( .a ({signal_2532, signal_1639}), .b ({signal_2647, signal_1703}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1503 ( .a ({signal_2533, signal_1640}), .b ({signal_2648, signal_1704}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1504 ( .a ({signal_2534, signal_1641}), .b ({signal_2649, signal_1705}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1505 ( .a ({signal_2535, signal_1642}), .b ({signal_2650, signal_1706}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1506 ( .a ({signal_2536, signal_1643}), .b ({signal_2651, signal_1707}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1507 ( .a ({signal_2537, signal_1644}), .b ({signal_2652, signal_1708}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1508 ( .a ({signal_2538, signal_1645}), .b ({signal_2653, signal_1709}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1509 ( .a ({signal_2539, signal_1646}), .b ({signal_2654, signal_1710}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1510 ( .a ({signal_2540, signal_1647}), .b ({signal_2655, signal_1711}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1511 ( .a ({signal_2280, signal_1517}), .b ({signal_2445, signal_1552}), .clk (clk), .r (Fresh[96]), .c ({signal_2656, signal_1712}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1512 ( .a ({signal_2272, signal_1513}), .b ({signal_2446, signal_1553}), .clk (clk), .r (Fresh[97]), .c ({signal_2657, signal_1713}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1513 ( .a ({signal_2264, signal_1509}), .b ({signal_2447, signal_1554}), .clk (clk), .r (Fresh[98]), .c ({signal_2658, signal_1714}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1514 ( .a ({signal_2256, signal_1505}), .b ({signal_2448, signal_1555}), .clk (clk), .r (Fresh[99]), .c ({signal_2659, signal_1715}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1515 ( .a ({signal_2248, signal_1501}), .b ({signal_2449, signal_1556}), .clk (clk), .r (Fresh[100]), .c ({signal_2660, signal_1716}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1516 ( .a ({signal_2240, signal_1497}), .b ({signal_2450, signal_1557}), .clk (clk), .r (Fresh[101]), .c ({signal_2661, signal_1717}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1517 ( .a ({signal_2232, signal_1493}), .b ({signal_2451, signal_1558}), .clk (clk), .r (Fresh[102]), .c ({signal_2662, signal_1718}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1518 ( .a ({signal_2224, signal_1489}), .b ({signal_2452, signal_1559}), .clk (clk), .r (Fresh[103]), .c ({signal_2663, signal_1719}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1519 ( .a ({signal_2216, signal_1485}), .b ({signal_2453, signal_1560}), .clk (clk), .r (Fresh[104]), .c ({signal_2664, signal_1720}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1520 ( .a ({signal_2208, signal_1481}), .b ({signal_2454, signal_1561}), .clk (clk), .r (Fresh[105]), .c ({signal_2665, signal_1721}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1521 ( .a ({signal_2200, signal_1477}), .b ({signal_2455, signal_1562}), .clk (clk), .r (Fresh[106]), .c ({signal_2666, signal_1722}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1522 ( .a ({signal_2192, signal_1473}), .b ({signal_2456, signal_1563}), .clk (clk), .r (Fresh[107]), .c ({signal_2667, signal_1723}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1523 ( .a ({signal_2184, signal_1469}), .b ({signal_2457, signal_1564}), .clk (clk), .r (Fresh[108]), .c ({signal_2668, signal_1724}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1524 ( .a ({signal_2176, signal_1465}), .b ({signal_2458, signal_1565}), .clk (clk), .r (Fresh[109]), .c ({signal_2669, signal_1725}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1525 ( .a ({signal_2168, signal_1461}), .b ({signal_2459, signal_1566}), .clk (clk), .r (Fresh[110]), .c ({signal_2670, signal_1726}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1526 ( .a ({signal_2160, signal_1457}), .b ({signal_2460, signal_1567}), .clk (clk), .r (Fresh[111]), .c ({signal_2671, signal_1727}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1527 ( .a ({signal_2282, signal_1518}), .b ({signal_2461, signal_1568}), .clk (clk), .r (Fresh[112]), .c ({signal_2672, signal_1728}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1528 ( .a ({signal_2274, signal_1514}), .b ({signal_2462, signal_1569}), .clk (clk), .r (Fresh[113]), .c ({signal_2673, signal_1729}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1529 ( .a ({signal_2266, signal_1510}), .b ({signal_2463, signal_1570}), .clk (clk), .r (Fresh[114]), .c ({signal_2674, signal_1730}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1530 ( .a ({signal_2258, signal_1506}), .b ({signal_2464, signal_1571}), .clk (clk), .r (Fresh[115]), .c ({signal_2675, signal_1731}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1531 ( .a ({signal_2250, signal_1502}), .b ({signal_2465, signal_1572}), .clk (clk), .r (Fresh[116]), .c ({signal_2676, signal_1732}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1532 ( .a ({signal_2242, signal_1498}), .b ({signal_2466, signal_1573}), .clk (clk), .r (Fresh[117]), .c ({signal_2677, signal_1733}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1533 ( .a ({signal_2234, signal_1494}), .b ({signal_2467, signal_1574}), .clk (clk), .r (Fresh[118]), .c ({signal_2678, signal_1734}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1534 ( .a ({signal_2226, signal_1490}), .b ({signal_2468, signal_1575}), .clk (clk), .r (Fresh[119]), .c ({signal_2679, signal_1735}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1535 ( .a ({signal_2218, signal_1486}), .b ({signal_2469, signal_1576}), .clk (clk), .r (Fresh[120]), .c ({signal_2680, signal_1736}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1536 ( .a ({signal_2210, signal_1482}), .b ({signal_2470, signal_1577}), .clk (clk), .r (Fresh[121]), .c ({signal_2681, signal_1737}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1537 ( .a ({signal_2202, signal_1478}), .b ({signal_2471, signal_1578}), .clk (clk), .r (Fresh[122]), .c ({signal_2682, signal_1738}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1538 ( .a ({signal_2194, signal_1474}), .b ({signal_2472, signal_1579}), .clk (clk), .r (Fresh[123]), .c ({signal_2683, signal_1739}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1539 ( .a ({signal_2186, signal_1470}), .b ({signal_2473, signal_1580}), .clk (clk), .r (Fresh[124]), .c ({signal_2684, signal_1740}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1540 ( .a ({signal_2178, signal_1466}), .b ({signal_2474, signal_1581}), .clk (clk), .r (Fresh[125]), .c ({signal_2685, signal_1741}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1541 ( .a ({signal_2170, signal_1462}), .b ({signal_2475, signal_1582}), .clk (clk), .r (Fresh[126]), .c ({signal_2686, signal_1742}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1542 ( .a ({signal_2162, signal_1458}), .b ({signal_2476, signal_1583}), .clk (clk), .r (Fresh[127]), .c ({signal_2687, signal_1743}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1543 ( .a ({signal_2656, signal_1712}), .b ({signal_2688, signal_1744}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1544 ( .a ({signal_2657, signal_1713}), .b ({signal_2689, signal_1745}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1545 ( .a ({signal_2658, signal_1714}), .b ({signal_2690, signal_1746}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1546 ( .a ({signal_2659, signal_1715}), .b ({signal_2691, signal_1747}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1547 ( .a ({signal_2660, signal_1716}), .b ({signal_2692, signal_1748}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1548 ( .a ({signal_2661, signal_1717}), .b ({signal_2693, signal_1749}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1549 ( .a ({signal_2662, signal_1718}), .b ({signal_2694, signal_1750}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1550 ( .a ({signal_2663, signal_1719}), .b ({signal_2695, signal_1751}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1551 ( .a ({signal_2664, signal_1720}), .b ({signal_2696, signal_1752}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1552 ( .a ({signal_2665, signal_1721}), .b ({signal_2697, signal_1753}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1553 ( .a ({signal_2666, signal_1722}), .b ({signal_2698, signal_1754}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1554 ( .a ({signal_2667, signal_1723}), .b ({signal_2699, signal_1755}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1555 ( .a ({signal_2668, signal_1724}), .b ({signal_2700, signal_1756}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1556 ( .a ({signal_2669, signal_1725}), .b ({signal_2701, signal_1757}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1557 ( .a ({signal_2670, signal_1726}), .b ({signal_2702, signal_1758}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1558 ( .a ({signal_2671, signal_1727}), .b ({signal_2703, signal_1759}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1559 ( .a ({signal_2672, signal_1728}), .b ({signal_2704, signal_1760}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1560 ( .a ({signal_2673, signal_1729}), .b ({signal_2705, signal_1761}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1561 ( .a ({signal_2674, signal_1730}), .b ({signal_2706, signal_1762}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1562 ( .a ({signal_2675, signal_1731}), .b ({signal_2707, signal_1763}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1563 ( .a ({signal_2676, signal_1732}), .b ({signal_2708, signal_1764}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1564 ( .a ({signal_2677, signal_1733}), .b ({signal_2709, signal_1765}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1565 ( .a ({signal_2678, signal_1734}), .b ({signal_2710, signal_1766}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1566 ( .a ({signal_2679, signal_1735}), .b ({signal_2711, signal_1767}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1567 ( .a ({signal_2680, signal_1736}), .b ({signal_2712, signal_1768}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1568 ( .a ({signal_2681, signal_1737}), .b ({signal_2713, signal_1769}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1569 ( .a ({signal_2682, signal_1738}), .b ({signal_2714, signal_1770}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1570 ( .a ({signal_2683, signal_1739}), .b ({signal_2715, signal_1771}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1571 ( .a ({signal_2684, signal_1740}), .b ({signal_2716, signal_1772}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1572 ( .a ({signal_2685, signal_1741}), .b ({signal_2717, signal_1773}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1573 ( .a ({signal_2686, signal_1742}), .b ({signal_2718, signal_1774}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1574 ( .a ({signal_2687, signal_1743}), .b ({signal_2719, signal_1775}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1575 ( .a ({signal_2283, signal_1375}), .b ({signal_2592, signal_1648}), .clk (clk), .r (Fresh[128]), .c ({signal_2720, signal_1776}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1576 ( .a ({signal_2275, signal_1371}), .b ({signal_2593, signal_1649}), .clk (clk), .r (Fresh[129]), .c ({signal_2721, signal_1777}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1577 ( .a ({signal_2267, signal_1367}), .b ({signal_2594, signal_1650}), .clk (clk), .r (Fresh[130]), .c ({signal_2722, signal_1778}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1578 ( .a ({signal_2259, signal_1363}), .b ({signal_2595, signal_1651}), .clk (clk), .r (Fresh[131]), .c ({signal_2723, signal_1779}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1579 ( .a ({signal_2251, signal_1359}), .b ({signal_2596, signal_1652}), .clk (clk), .r (Fresh[132]), .c ({signal_2724, signal_1780}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1580 ( .a ({signal_2243, signal_1355}), .b ({signal_2597, signal_1653}), .clk (clk), .r (Fresh[133]), .c ({signal_2725, signal_1781}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1581 ( .a ({signal_2235, signal_1351}), .b ({signal_2598, signal_1654}), .clk (clk), .r (Fresh[134]), .c ({signal_2726, signal_1782}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1582 ( .a ({signal_2227, signal_1347}), .b ({signal_2599, signal_1655}), .clk (clk), .r (Fresh[135]), .c ({signal_2727, signal_1783}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1583 ( .a ({signal_2219, signal_1343}), .b ({signal_2600, signal_1656}), .clk (clk), .r (Fresh[136]), .c ({signal_2728, signal_1784}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1584 ( .a ({signal_2211, signal_1339}), .b ({signal_2601, signal_1657}), .clk (clk), .r (Fresh[137]), .c ({signal_2729, signal_1785}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1585 ( .a ({signal_2203, signal_1335}), .b ({signal_2602, signal_1658}), .clk (clk), .r (Fresh[138]), .c ({signal_2730, signal_1786}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1586 ( .a ({signal_2195, signal_1331}), .b ({signal_2603, signal_1659}), .clk (clk), .r (Fresh[139]), .c ({signal_2731, signal_1787}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1587 ( .a ({signal_2187, signal_1327}), .b ({signal_2604, signal_1660}), .clk (clk), .r (Fresh[140]), .c ({signal_2732, signal_1788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1588 ( .a ({signal_2179, signal_1323}), .b ({signal_2605, signal_1661}), .clk (clk), .r (Fresh[141]), .c ({signal_2733, signal_1789}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1589 ( .a ({signal_2171, signal_1319}), .b ({signal_2606, signal_1662}), .clk (clk), .r (Fresh[142]), .c ({signal_2734, signal_1790}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1590 ( .a ({signal_2163, signal_1315}), .b ({signal_2607, signal_1663}), .clk (clk), .r (Fresh[143]), .c ({signal_2735, signal_1791}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1591 ( .a ({signal_2283, signal_1375}), .b ({signal_2609, signal_1665}), .clk (clk), .r (Fresh[144]), .c ({signal_2736, signal_1792}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1592 ( .a ({signal_2275, signal_1371}), .b ({signal_2612, signal_1668}), .clk (clk), .r (Fresh[145]), .c ({signal_2737, signal_1793}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1593 ( .a ({signal_2267, signal_1367}), .b ({signal_2615, signal_1671}), .clk (clk), .r (Fresh[146]), .c ({signal_2738, signal_1794}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1594 ( .a ({signal_2259, signal_1363}), .b ({signal_2618, signal_1674}), .clk (clk), .r (Fresh[147]), .c ({signal_2739, signal_1795}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1595 ( .a ({signal_2251, signal_1359}), .b ({signal_2621, signal_1677}), .clk (clk), .r (Fresh[148]), .c ({signal_2740, signal_1796}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1596 ( .a ({signal_2243, signal_1355}), .b ({signal_2624, signal_1680}), .clk (clk), .r (Fresh[149]), .c ({signal_2741, signal_1797}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1597 ( .a ({signal_2235, signal_1351}), .b ({signal_2627, signal_1683}), .clk (clk), .r (Fresh[150]), .c ({signal_2742, signal_1798}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1598 ( .a ({signal_2227, signal_1347}), .b ({signal_2630, signal_1686}), .clk (clk), .r (Fresh[151]), .c ({signal_2743, signal_1799}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1599 ( .a ({signal_2219, signal_1343}), .b ({signal_2633, signal_1689}), .clk (clk), .r (Fresh[152]), .c ({signal_2744, signal_1800}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1600 ( .a ({signal_2211, signal_1339}), .b ({signal_2636, signal_1692}), .clk (clk), .r (Fresh[153]), .c ({signal_2745, signal_1801}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1601 ( .a ({signal_2203, signal_1335}), .b ({signal_2639, signal_1695}), .clk (clk), .r (Fresh[154]), .c ({signal_2746, signal_1802}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1602 ( .a ({signal_2195, signal_1331}), .b ({signal_2642, signal_1698}), .clk (clk), .r (Fresh[155]), .c ({signal_2747, signal_1803}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1603 ( .a ({signal_2187, signal_1327}), .b ({signal_2645, signal_1701}), .clk (clk), .r (Fresh[156]), .c ({signal_2748, signal_1804}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1604 ( .a ({signal_2179, signal_1323}), .b ({signal_2648, signal_1704}), .clk (clk), .r (Fresh[157]), .c ({signal_2749, signal_1805}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1605 ( .a ({signal_2171, signal_1319}), .b ({signal_2651, signal_1707}), .clk (clk), .r (Fresh[158]), .c ({signal_2750, signal_1806}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1606 ( .a ({signal_2163, signal_1315}), .b ({signal_2654, signal_1710}), .clk (clk), .r (Fresh[159]), .c ({signal_2751, signal_1807}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1607 ( .a ({signal_2720, signal_1776}), .b ({signal_2752, signal_1808}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1608 ( .a ({signal_2721, signal_1777}), .b ({signal_2753, signal_1809}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1609 ( .a ({signal_2722, signal_1778}), .b ({signal_2754, signal_1810}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1610 ( .a ({signal_2723, signal_1779}), .b ({signal_2755, signal_1811}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1611 ( .a ({signal_2724, signal_1780}), .b ({signal_2756, signal_1812}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1612 ( .a ({signal_2725, signal_1781}), .b ({signal_2757, signal_1813}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1613 ( .a ({signal_2726, signal_1782}), .b ({signal_2758, signal_1814}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1614 ( .a ({signal_2727, signal_1783}), .b ({signal_2759, signal_1815}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1615 ( .a ({signal_2728, signal_1784}), .b ({signal_2760, signal_1816}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1616 ( .a ({signal_2729, signal_1785}), .b ({signal_2761, signal_1817}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1617 ( .a ({signal_2730, signal_1786}), .b ({signal_2762, signal_1818}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1618 ( .a ({signal_2731, signal_1787}), .b ({signal_2763, signal_1819}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1619 ( .a ({signal_2732, signal_1788}), .b ({signal_2764, signal_1820}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1620 ( .a ({signal_2733, signal_1789}), .b ({signal_2765, signal_1821}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1621 ( .a ({signal_2734, signal_1790}), .b ({signal_2766, signal_1822}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1622 ( .a ({signal_2735, signal_1791}), .b ({signal_2767, signal_1823}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1623 ( .a ({signal_2736, signal_1792}), .b ({signal_2768, signal_1824}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1624 ( .a ({signal_2737, signal_1793}), .b ({signal_2769, signal_1825}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1625 ( .a ({signal_2738, signal_1794}), .b ({signal_2770, signal_1826}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1626 ( .a ({signal_2739, signal_1795}), .b ({signal_2771, signal_1827}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1627 ( .a ({signal_2740, signal_1796}), .b ({signal_2772, signal_1828}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1628 ( .a ({signal_2741, signal_1797}), .b ({signal_2773, signal_1829}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1629 ( .a ({signal_2742, signal_1798}), .b ({signal_2774, signal_1830}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1630 ( .a ({signal_2743, signal_1799}), .b ({signal_2775, signal_1831}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1631 ( .a ({signal_2744, signal_1800}), .b ({signal_2776, signal_1832}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1632 ( .a ({signal_2745, signal_1801}), .b ({signal_2777, signal_1833}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1633 ( .a ({signal_2746, signal_1802}), .b ({signal_2778, signal_1834}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1634 ( .a ({signal_2747, signal_1803}), .b ({signal_2779, signal_1835}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1635 ( .a ({signal_2748, signal_1804}), .b ({signal_2780, signal_1836}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1636 ( .a ({signal_2749, signal_1805}), .b ({signal_2781, signal_1837}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1637 ( .a ({signal_2750, signal_1806}), .b ({signal_2782, signal_1838}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1638 ( .a ({signal_2751, signal_1807}), .b ({signal_2783, signal_1839}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_89 ( .a ({signal_1954, signal_914}), .b ({signal_2930, signal_1302}), .c ({DataOut_s1[9], DataOut_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_91 ( .a ({signal_1960, signal_916}), .b ({signal_2833, signal_1264}), .c ({DataOut_s1[7], DataOut_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_93 ( .a ({signal_1966, signal_860}), .b ({signal_2847, signal_1248}), .c ({DataOut_s1[63], DataOut_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_95 ( .a ({signal_1972, signal_862}), .b ({signal_2943, signal_1250}), .c ({DataOut_s1[61], DataOut_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_97 ( .a ({signal_1978, signal_918}), .b ({signal_2929, signal_1266}), .c ({DataOut_s1[5], DataOut_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_98 ( .a ({signal_1981, signal_864}), .b ({signal_2846, signal_1276}), .c ({DataOut_s1[59], DataOut_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_100 ( .a ({signal_1987, signal_866}), .b ({signal_2942, signal_1278}), .c ({DataOut_s1[57], DataOut_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_102 ( .a ({signal_1993, signal_868}), .b ({signal_2845, signal_1304}), .c ({DataOut_s1[55], DataOut_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_104 ( .a ({signal_1999, signal_870}), .b ({signal_2941, signal_1306}), .c ({DataOut_s1[53], DataOut_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_106 ( .a ({signal_2005, signal_872}), .b ({signal_2844, signal_1284}), .c ({DataOut_s1[51], DataOut_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_109 ( .a ({signal_2014, signal_874}), .b ({signal_2940, signal_1286}), .c ({DataOut_s1[49], DataOut_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_111 ( .a ({signal_2020, signal_876}), .b ({signal_2843, signal_1268}), .c ({DataOut_s1[47], DataOut_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_113 ( .a ({signal_2026, signal_878}), .b ({signal_2939, signal_1270}), .c ({DataOut_s1[45], DataOut_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_115 ( .a ({signal_2032, signal_880}), .b ({signal_2842, signal_1256}), .c ({DataOut_s1[43], DataOut_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_117 ( .a ({signal_2038, signal_882}), .b ({signal_2938, signal_1258}), .c ({DataOut_s1[41], DataOut_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_119 ( .a ({signal_2044, signal_920}), .b ({signal_2832, signal_1260}), .c ({DataOut_s1[3], DataOut_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_120 ( .a ({signal_2047, signal_884}), .b ({signal_2841, signal_1292}), .c ({DataOut_s1[39], DataOut_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_122 ( .a ({signal_2053, signal_886}), .b ({signal_2937, signal_1294}), .c ({DataOut_s1[37], DataOut_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_124 ( .a ({signal_2059, signal_888}), .b ({signal_2840, signal_1296}), .c ({DataOut_s1[35], DataOut_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_126 ( .a ({signal_2065, signal_890}), .b ({signal_2936, signal_1298}), .c ({DataOut_s1[33], DataOut_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_128 ( .a ({signal_2071, signal_892}), .b ({signal_2839, signal_1308}), .c ({DataOut_s1[31], DataOut_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_131 ( .a ({signal_2080, signal_894}), .b ({signal_2935, signal_1310}), .c ({DataOut_s1[29], DataOut_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_133 ( .a ({signal_2086, signal_896}), .b ({signal_2838, signal_1280}), .c ({DataOut_s1[27], DataOut_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_135 ( .a ({signal_2092, signal_898}), .b ({signal_2934, signal_1282}), .c ({DataOut_s1[25], DataOut_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_137 ( .a ({signal_2098, signal_900}), .b ({signal_2837, signal_1252}), .c ({DataOut_s1[23], DataOut_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_139 ( .a ({signal_2104, signal_902}), .b ({signal_2933, signal_1254}), .c ({DataOut_s1[21], DataOut_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_141 ( .a ({signal_2110, signal_922}), .b ({signal_2928, signal_1262}), .c ({DataOut_s1[1], DataOut_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_142 ( .a ({signal_2113, signal_904}), .b ({signal_2836, signal_1272}), .c ({DataOut_s1[19], DataOut_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_144 ( .a ({signal_2119, signal_906}), .b ({signal_2932, signal_1274}), .c ({DataOut_s1[17], DataOut_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_146 ( .a ({signal_2125, signal_908}), .b ({signal_2835, signal_1288}), .c ({DataOut_s1[15], DataOut_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_148 ( .a ({signal_2131, signal_910}), .b ({signal_2931, signal_1290}), .c ({DataOut_s1[13], DataOut_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_150 ( .a ({signal_2137, signal_912}), .b ({signal_2834, signal_1300}), .c ({DataOut_s1[11], DataOut_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_217 ( .a ({signal_2150, signal_311}), .b ({signal_2930, signal_1302}), .c ({signal_2976, signal_1238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_219 ( .a ({signal_2543, signal_309}), .b ({signal_2833, signal_1264}), .c ({signal_2896, signal_1240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_221 ( .a ({signal_2591, signal_365}), .b ({signal_2847, signal_1248}), .c ({signal_2897, signal_1184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_223 ( .a ({signal_2589, signal_363}), .b ({signal_2943, signal_1250}), .c ({signal_2977, signal_1186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_225 ( .a ({signal_2541, signal_307}), .b ({signal_2929, signal_1266}), .c ({signal_2978, signal_1242}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_226 ( .a ({signal_2587, signal_361}), .b ({signal_2846, signal_1276}), .c ({signal_2898, signal_1188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_228 ( .a ({signal_2585, signal_359}), .b ({signal_2942, signal_1278}), .c ({signal_2979, signal_1190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_230 ( .a ({signal_2583, signal_357}), .b ({signal_2845, signal_1304}), .c ({signal_2899, signal_1192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_232 ( .a ({signal_2581, signal_355}), .b ({signal_2941, signal_1306}), .c ({signal_2980, signal_1194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_234 ( .a ({signal_2579, signal_353}), .b ({signal_2844, signal_1284}), .c ({signal_2900, signal_1196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({signal_2577, signal_351}), .b ({signal_2940, signal_1286}), .c ({signal_2981, signal_1198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({signal_2575, signal_349}), .b ({signal_2843, signal_1268}), .c ({signal_2901, signal_1200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({signal_2573, signal_347}), .b ({signal_2939, signal_1270}), .c ({signal_2982, signal_1202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({signal_2571, signal_345}), .b ({signal_2842, signal_1256}), .c ({signal_2902, signal_1204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({signal_2569, signal_343}), .b ({signal_2938, signal_1258}), .c ({signal_2983, signal_1206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({signal_2147, signal_305}), .b ({signal_2832, signal_1260}), .c ({signal_2903, signal_1244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({signal_2567, signal_341}), .b ({signal_2841, signal_1292}), .c ({signal_2904, signal_1208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({signal_2565, signal_339}), .b ({signal_2937, signal_1294}), .c ({signal_2984, signal_1210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({signal_2563, signal_337}), .b ({signal_2840, signal_1296}), .c ({signal_2905, signal_1212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({signal_2561, signal_335}), .b ({signal_2936, signal_1298}), .c ({signal_2985, signal_1214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({signal_2559, signal_333}), .b ({signal_2839, signal_1308}), .c ({signal_2906, signal_1216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .a ({signal_2557, signal_331}), .b ({signal_2935, signal_1310}), .c ({signal_2986, signal_1218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .a ({signal_2555, signal_329}), .b ({signal_2838, signal_1280}), .c ({signal_2907, signal_1220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({signal_2554, signal_327}), .b ({signal_2934, signal_1282}), .c ({signal_2987, signal_1222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({signal_2552, signal_325}), .b ({signal_2837, signal_1252}), .c ({signal_2908, signal_1224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .a ({signal_2550, signal_323}), .b ({signal_2933, signal_1254}), .c ({signal_2988, signal_1226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({signal_2145, signal_303}), .b ({signal_2928, signal_1262}), .c ({signal_2989, signal_1246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({signal_2548, signal_321}), .b ({signal_2836, signal_1272}), .c ({signal_2909, signal_1228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({signal_2546, signal_319}), .b ({signal_2932, signal_1274}), .c ({signal_2990, signal_1230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({signal_2155, signal_317}), .b ({signal_2835, signal_1288}), .c ({signal_2910, signal_1232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({signal_2153, signal_315}), .b ({signal_2931, signal_1290}), .c ({signal_2991, signal_1234}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({signal_2152, signal_313}), .b ({signal_2834, signal_1300}), .c ({signal_2911, signal_1236}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_281 ( .a ({signal_2150, signal_311}), .b ({signal_3219, signal_1110}), .c ({signal_3226, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_284 ( .a ({signal_2543, signal_309}), .b ({signal_3164, signal_1064}), .c ({signal_3180, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_286 ( .a ({signal_2591, signal_365}), .b ({signal_3149, signal_1056}), .c ({signal_3181, signal_992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_288 ( .a ({signal_2589, signal_363}), .b ({signal_3205, signal_1058}), .c ({signal_3227, signal_994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_291 ( .a ({signal_2541, signal_307}), .b ({signal_3220, signal_1066}), .c ({signal_3228, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_292 ( .a ({signal_2587, signal_361}), .b ({signal_3151, signal_1096}), .c ({signal_3182, signal_996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_294 ( .a ({signal_2585, signal_359}), .b ({signal_3201, signal_1098}), .c ({signal_3229, signal_998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_297 ( .a ({signal_2583, signal_357}), .b ({signal_3146, signal_1076}), .c ({signal_3183, signal_1000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_299 ( .a ({signal_2581, signal_355}), .b ({signal_3202, signal_1078}), .c ({signal_3230, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_302 ( .a ({signal_2579, signal_353}), .b ({signal_3147, signal_1116}), .c ({signal_3184, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_306 ( .a ({signal_2577, signal_351}), .b ({signal_3204, signal_1118}), .c ({signal_3231, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_309 ( .a ({signal_2575, signal_349}), .b ({signal_3155, signal_1112}), .c ({signal_3185, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_311 ( .a ({signal_2573, signal_347}), .b ({signal_3211, signal_1114}), .c ({signal_3233, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_314 ( .a ({signal_2571, signal_345}), .b ({signal_3157, signal_1072}), .c ({signal_3186, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_316 ( .a ({signal_2569, signal_343}), .b ({signal_3207, signal_1074}), .c ({signal_3234, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_319 ( .a ({signal_2147, signal_305}), .b ({signal_3165, signal_1088}), .c ({signal_3187, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_320 ( .a ({signal_2567, signal_341}), .b ({signal_3152, signal_1100}), .c ({signal_3188, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_322 ( .a ({signal_2565, signal_339}), .b ({signal_3208, signal_1102}), .c ({signal_3235, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_325 ( .a ({signal_2563, signal_337}), .b ({signal_3153, signal_1060}), .c ({signal_3189, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_327 ( .a ({signal_2561, signal_335}), .b ({signal_3210, signal_1062}), .c ({signal_3236, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_330 ( .a ({signal_2559, signal_333}), .b ({signal_3161, signal_1092}), .c ({signal_3190, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_333 ( .a ({signal_2557, signal_331}), .b ({signal_3217, signal_1094}), .c ({signal_3237, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_336 ( .a ({signal_2555, signal_329}), .b ({signal_3163, signal_1068}), .c ({signal_3192, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_338 ( .a ({signal_2554, signal_327}), .b ({signal_3213, signal_1070}), .c ({signal_3238, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_341 ( .a ({signal_2552, signal_325}), .b ({signal_3158, signal_1104}), .c ({signal_3193, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_343 ( .a ({signal_2550, signal_323}), .b ({signal_3214, signal_1106}), .c ({signal_3239, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_346 ( .a ({signal_2145, signal_303}), .b ({signal_3222, signal_1090}), .c ({signal_3240, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_347 ( .a ({signal_2548, signal_321}), .b ({signal_3159, signal_1080}), .c ({signal_3194, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_349 ( .a ({signal_2546, signal_319}), .b ({signal_3216, signal_1082}), .c ({signal_3241, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_352 ( .a ({signal_2155, signal_317}), .b ({signal_3167, signal_1084}), .c ({signal_3195, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_354 ( .a ({signal_2153, signal_315}), .b ({signal_3223, signal_1086}), .c ({signal_3242, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_357 ( .a ({signal_2152, signal_313}), .b ({signal_3169, signal_1108}), .c ({signal_3196, signal_1044}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_538 ( .s (reset), .b ({signal_3325, signal_1438}), .a ({signal_2422, signal_990}), .c ({signal_3341, signal_462}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_544 ( .s (reset), .b ({signal_3269, signal_1436}), .a ({signal_2378, signal_988}), .c ({signal_3302, signal_466}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_550 ( .s (reset), .b ({signal_3326, signal_1434}), .a ({signal_2334, signal_986}), .c ({signal_3342, signal_470}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_556 ( .s (reset), .b ({signal_3270, signal_1432}), .a ({signal_2322, signal_984}), .c ({signal_3303, signal_474}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_562 ( .s (reset), .b ({signal_3327, signal_1430}), .a ({signal_2318, signal_982}), .c ({signal_3343, signal_478}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_568 ( .s (reset), .b ({signal_3271, signal_1428}), .a ({signal_2440, signal_980}), .c ({signal_3304, signal_482}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_574 ( .s (reset), .b ({signal_3328, signal_1426}), .a ({signal_2436, signal_978}), .c ({signal_3344, signal_486}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_580 ( .s (reset), .b ({signal_3272, signal_1424}), .a ({signal_2432, signal_976}), .c ({signal_3305, signal_490}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_586 ( .s (reset), .b ({signal_3329, signal_1422}), .a ({signal_2428, signal_974}), .c ({signal_3345, signal_494}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_592 ( .s (reset), .b ({signal_3273, signal_1420}), .a ({signal_2424, signal_972}), .c ({signal_3306, signal_498}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_598 ( .s (reset), .b ({signal_3330, signal_1418}), .a ({signal_2418, signal_970}), .c ({signal_3346, signal_502}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_604 ( .s (reset), .b ({signal_3274, signal_1416}), .a ({signal_2414, signal_968}), .c ({signal_3307, signal_506}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_610 ( .s (reset), .b ({signal_3331, signal_1414}), .a ({signal_2410, signal_966}), .c ({signal_3347, signal_510}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_616 ( .s (reset), .b ({signal_3275, signal_1412}), .a ({signal_2406, signal_964}), .c ({signal_3308, signal_514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_622 ( .s (reset), .b ({signal_3332, signal_1410}), .a ({signal_2402, signal_962}), .c ({signal_3348, signal_518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_628 ( .s (reset), .b ({signal_3276, signal_1408}), .a ({signal_2396, signal_960}), .c ({signal_3309, signal_522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_634 ( .s (reset), .b ({signal_3333, signal_1406}), .a ({signal_2392, signal_958}), .c ({signal_3349, signal_526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_640 ( .s (reset), .b ({signal_3277, signal_1404}), .a ({signal_2388, signal_956}), .c ({signal_3310, signal_530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_646 ( .s (reset), .b ({signal_3334, signal_1402}), .a ({signal_2384, signal_954}), .c ({signal_3350, signal_534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_652 ( .s (reset), .b ({signal_3278, signal_1400}), .a ({signal_2380, signal_952}), .c ({signal_3311, signal_538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_658 ( .s (reset), .b ({signal_3335, signal_1398}), .a ({signal_2374, signal_950}), .c ({signal_3351, signal_542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_664 ( .s (reset), .b ({signal_3279, signal_1396}), .a ({signal_2370, signal_948}), .c ({signal_3312, signal_546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_670 ( .s (reset), .b ({signal_3336, signal_1394}), .a ({signal_2366, signal_946}), .c ({signal_3352, signal_550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_676 ( .s (reset), .b ({signal_3280, signal_1392}), .a ({signal_2362, signal_944}), .c ({signal_3313, signal_554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_682 ( .s (reset), .b ({signal_3337, signal_1390}), .a ({signal_2358, signal_942}), .c ({signal_3353, signal_558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_688 ( .s (reset), .b ({signal_3281, signal_1388}), .a ({signal_2352, signal_940}), .c ({signal_3314, signal_562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_694 ( .s (reset), .b ({signal_3338, signal_1386}), .a ({signal_2348, signal_938}), .c ({signal_3354, signal_566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_700 ( .s (reset), .b ({signal_3282, signal_1384}), .a ({signal_2344, signal_936}), .c ({signal_3315, signal_570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_706 ( .s (reset), .b ({signal_3339, signal_1382}), .a ({signal_2340, signal_934}), .c ({signal_3355, signal_574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_712 ( .s (reset), .b ({signal_3283, signal_1380}), .a ({signal_2336, signal_932}), .c ({signal_3316, signal_578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_718 ( .s (reset), .b ({signal_3340, signal_1378}), .a ({signal_2330, signal_930}), .c ({signal_3356, signal_582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_724 ( .s (reset), .b ({signal_3284, signal_1376}), .a ({signal_2326, signal_928}), .c ({signal_3317, signal_586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1032 ( .s (enc_dec), .b ({signal_2935, signal_1310}), .a ({signal_2989, signal_1246}), .c ({signal_3092, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1034 ( .s (enc_dec), .b ({signal_2839, signal_1308}), .a ({signal_2903, signal_1244}), .c ({signal_2992, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1036 ( .s (enc_dec), .b ({signal_2941, signal_1306}), .a ({signal_2978, signal_1242}), .c ({signal_3093, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1038 ( .s (enc_dec), .b ({signal_2845, signal_1304}), .a ({signal_2896, signal_1240}), .c ({signal_2993, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1040 ( .s (enc_dec), .b ({signal_2930, signal_1302}), .a ({signal_2976, signal_1238}), .c ({signal_3094, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1042 ( .s (enc_dec), .b ({signal_2834, signal_1300}), .a ({signal_2911, signal_1236}), .c ({signal_2994, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1044 ( .s (enc_dec), .b ({signal_2936, signal_1298}), .a ({signal_2991, signal_1234}), .c ({signal_3095, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1046 ( .s (enc_dec), .b ({signal_2840, signal_1296}), .a ({signal_2910, signal_1232}), .c ({signal_2995, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1048 ( .s (enc_dec), .b ({signal_2937, signal_1294}), .a ({signal_2990, signal_1230}), .c ({signal_3096, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1050 ( .s (enc_dec), .b ({signal_2841, signal_1292}), .a ({signal_2909, signal_1228}), .c ({signal_2996, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1052 ( .s (enc_dec), .b ({signal_2931, signal_1290}), .a ({signal_2988, signal_1226}), .c ({signal_3097, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1054 ( .s (enc_dec), .b ({signal_2835, signal_1288}), .a ({signal_2908, signal_1224}), .c ({signal_2997, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1056 ( .s (enc_dec), .b ({signal_2940, signal_1286}), .a ({signal_2987, signal_1222}), .c ({signal_3098, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1058 ( .s (enc_dec), .b ({signal_2844, signal_1284}), .a ({signal_2907, signal_1220}), .c ({signal_2998, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1060 ( .s (enc_dec), .b ({signal_2934, signal_1282}), .a ({signal_2986, signal_1218}), .c ({signal_3099, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1062 ( .s (enc_dec), .b ({signal_2838, signal_1280}), .a ({signal_2906, signal_1216}), .c ({signal_2999, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1064 ( .s (enc_dec), .b ({signal_2942, signal_1278}), .a ({signal_2985, signal_1214}), .c ({signal_3100, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1066 ( .s (enc_dec), .b ({signal_2846, signal_1276}), .a ({signal_2905, signal_1212}), .c ({signal_3000, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1068 ( .s (enc_dec), .b ({signal_2932, signal_1274}), .a ({signal_2984, signal_1210}), .c ({signal_3101, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1070 ( .s (enc_dec), .b ({signal_2836, signal_1272}), .a ({signal_2904, signal_1208}), .c ({signal_3001, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1072 ( .s (enc_dec), .b ({signal_2939, signal_1270}), .a ({signal_2983, signal_1206}), .c ({signal_3102, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1074 ( .s (enc_dec), .b ({signal_2843, signal_1268}), .a ({signal_2902, signal_1204}), .c ({signal_3002, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1076 ( .s (enc_dec), .b ({signal_2929, signal_1266}), .a ({signal_2982, signal_1202}), .c ({signal_3103, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1078 ( .s (enc_dec), .b ({signal_2833, signal_1264}), .a ({signal_2901, signal_1200}), .c ({signal_3003, signal_1136}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1080 ( .s (enc_dec), .b ({signal_2928, signal_1262}), .a ({signal_2981, signal_1198}), .c ({signal_3104, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1082 ( .s (enc_dec), .b ({signal_2832, signal_1260}), .a ({signal_2900, signal_1196}), .c ({signal_3004, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1084 ( .s (enc_dec), .b ({signal_2938, signal_1258}), .a ({signal_2980, signal_1194}), .c ({signal_3105, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1086 ( .s (enc_dec), .b ({signal_2842, signal_1256}), .a ({signal_2899, signal_1192}), .c ({signal_3005, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1088 ( .s (enc_dec), .b ({signal_2933, signal_1254}), .a ({signal_2979, signal_1190}), .c ({signal_3106, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1090 ( .s (enc_dec), .b ({signal_2837, signal_1252}), .a ({signal_2898, signal_1188}), .c ({signal_3006, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1092 ( .s (enc_dec), .b ({signal_2943, signal_1250}), .a ({signal_2977, signal_1186}), .c ({signal_3107, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1094 ( .s (enc_dec), .b ({signal_2847, signal_1248}), .a ({signal_2897, signal_1184}), .c ({signal_3007, signal_1120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .a ({signal_3107, signal_1122}), .b ({signal_3150, signal_828}), .c ({signal_3201, signal_1098}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .a ({signal_3004, signal_1132}), .b ({signal_3108, signal_830}), .c ({signal_3146, signal_1076}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .a ({signal_3104, signal_1134}), .b ({signal_3148, signal_832}), .c ({signal_3202, signal_1078}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .a ({signal_3005, signal_1128}), .b ({signal_3108, signal_830}), .c ({signal_3147, signal_1116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .a ({signal_3007, signal_1120}), .b ({signal_3006, signal_1124}), .c ({signal_3108, signal_830}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .a ({signal_3105, signal_1130}), .b ({signal_3148, signal_832}), .c ({signal_3204, signal_1118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .a ({signal_3106, signal_1126}), .b ({signal_3107, signal_1122}), .c ({signal_3148, signal_832}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1107 ( .a ({signal_3006, signal_1124}), .b ({signal_3109, signal_834}), .c ({signal_3149, signal_1056}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1109 ( .a ({signal_3106, signal_1126}), .b ({signal_3150, signal_828}), .c ({signal_3205, signal_1058}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1110 ( .a ({signal_3104, signal_1134}), .b ({signal_3105, signal_1130}), .c ({signal_3150, signal_828}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1113 ( .a ({signal_3007, signal_1120}), .b ({signal_3109, signal_834}), .c ({signal_3151, signal_1096}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1114 ( .a ({signal_3004, signal_1132}), .b ({signal_3005, signal_1128}), .c ({signal_3109, signal_834}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1119 ( .a ({signal_3103, signal_1138}), .b ({signal_3156, signal_836}), .c ({signal_3207, signal_1074}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1121 ( .a ({signal_3000, signal_1148}), .b ({signal_3110, signal_838}), .c ({signal_3152, signal_1100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1123 ( .a ({signal_3100, signal_1150}), .b ({signal_3154, signal_840}), .c ({signal_3208, signal_1102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1125 ( .a ({signal_3001, signal_1144}), .b ({signal_3110, signal_838}), .c ({signal_3153, signal_1060}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1126 ( .a ({signal_3003, signal_1136}), .b ({signal_3002, signal_1140}), .c ({signal_3110, signal_838}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1129 ( .a ({signal_3101, signal_1146}), .b ({signal_3154, signal_840}), .c ({signal_3210, signal_1062}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1130 ( .a ({signal_3102, signal_1142}), .b ({signal_3103, signal_1138}), .c ({signal_3154, signal_840}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1131 ( .a ({signal_3002, signal_1140}), .b ({signal_3111, signal_842}), .c ({signal_3155, signal_1112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1133 ( .a ({signal_3102, signal_1142}), .b ({signal_3156, signal_836}), .c ({signal_3211, signal_1114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1134 ( .a ({signal_3100, signal_1150}), .b ({signal_3101, signal_1146}), .c ({signal_3156, signal_836}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1137 ( .a ({signal_3003, signal_1136}), .b ({signal_3111, signal_842}), .c ({signal_3157, signal_1072}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1138 ( .a ({signal_3000, signal_1148}), .b ({signal_3001, signal_1144}), .c ({signal_3111, signal_842}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .a ({signal_3099, signal_1154}), .b ({signal_3162, signal_844}), .c ({signal_3213, signal_1070}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .a ({signal_2996, signal_1164}), .b ({signal_3112, signal_846}), .c ({signal_3158, signal_1104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .a ({signal_3096, signal_1166}), .b ({signal_3160, signal_848}), .c ({signal_3214, signal_1106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .a ({signal_2997, signal_1160}), .b ({signal_3112, signal_846}), .c ({signal_3159, signal_1080}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .a ({signal_2999, signal_1152}), .b ({signal_2998, signal_1156}), .c ({signal_3112, signal_846}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .a ({signal_3097, signal_1162}), .b ({signal_3160, signal_848}), .c ({signal_3216, signal_1082}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .a ({signal_3098, signal_1158}), .b ({signal_3099, signal_1154}), .c ({signal_3160, signal_848}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .a ({signal_2998, signal_1156}), .b ({signal_3113, signal_850}), .c ({signal_3161, signal_1092}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .a ({signal_3098, signal_1158}), .b ({signal_3162, signal_844}), .c ({signal_3217, signal_1094}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .a ({signal_3096, signal_1166}), .b ({signal_3097, signal_1162}), .c ({signal_3162, signal_844}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .a ({signal_2999, signal_1152}), .b ({signal_3113, signal_850}), .c ({signal_3163, signal_1068}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .a ({signal_2996, signal_1164}), .b ({signal_2997, signal_1160}), .c ({signal_3113, signal_850}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .a ({signal_3095, signal_1170}), .b ({signal_3168, signal_852}), .c ({signal_3219, signal_1110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .a ({signal_2992, signal_1180}), .b ({signal_3114, signal_854}), .c ({signal_3164, signal_1064}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .a ({signal_3092, signal_1182}), .b ({signal_3166, signal_856}), .c ({signal_3220, signal_1066}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .a ({signal_2993, signal_1176}), .b ({signal_3114, signal_854}), .c ({signal_3165, signal_1088}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .a ({signal_2995, signal_1168}), .b ({signal_2994, signal_1172}), .c ({signal_3114, signal_854}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .a ({signal_3093, signal_1178}), .b ({signal_3166, signal_856}), .c ({signal_3222, signal_1090}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .a ({signal_3094, signal_1174}), .b ({signal_3095, signal_1170}), .c ({signal_3166, signal_856}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .a ({signal_2994, signal_1172}), .b ({signal_3115, signal_858}), .c ({signal_3167, signal_1084}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_3094, signal_1174}), .b ({signal_3168, signal_852}), .c ({signal_3223, signal_1086}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .a ({signal_3092, signal_1182}), .b ({signal_3093, signal_1178}), .c ({signal_3168, signal_852}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .a ({signal_2995, signal_1168}), .b ({signal_3115, signal_858}), .c ({signal_3169, signal_1108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .a ({signal_2992, signal_1180}), .b ({signal_2993, signal_1176}), .c ({signal_3115, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1192 ( .s (enc_dec), .b ({signal_3240, signal_1054}), .a ({signal_3204, signal_1118}), .c ({signal_3325, signal_1438}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1194 ( .s (enc_dec), .b ({signal_3187, signal_1052}), .a ({signal_3147, signal_1116}), .c ({signal_3269, signal_1436}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1196 ( .s (enc_dec), .b ({signal_3228, signal_1050}), .a ({signal_3211, signal_1114}), .c ({signal_3326, signal_1434}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1198 ( .s (enc_dec), .b ({signal_3180, signal_1048}), .a ({signal_3155, signal_1112}), .c ({signal_3270, signal_1432}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1200 ( .s (enc_dec), .b ({signal_3226, signal_1046}), .a ({signal_3219, signal_1110}), .c ({signal_3327, signal_1430}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1202 ( .s (enc_dec), .b ({signal_3196, signal_1044}), .a ({signal_3169, signal_1108}), .c ({signal_3271, signal_1428}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1204 ( .s (enc_dec), .b ({signal_3242, signal_1042}), .a ({signal_3214, signal_1106}), .c ({signal_3328, signal_1426}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1206 ( .s (enc_dec), .b ({signal_3195, signal_1040}), .a ({signal_3158, signal_1104}), .c ({signal_3272, signal_1424}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1208 ( .s (enc_dec), .b ({signal_3241, signal_1038}), .a ({signal_3208, signal_1102}), .c ({signal_3329, signal_1422}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1210 ( .s (enc_dec), .b ({signal_3194, signal_1036}), .a ({signal_3152, signal_1100}), .c ({signal_3273, signal_1420}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1212 ( .s (enc_dec), .b ({signal_3239, signal_1034}), .a ({signal_3201, signal_1098}), .c ({signal_3330, signal_1418}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1214 ( .s (enc_dec), .b ({signal_3193, signal_1032}), .a ({signal_3151, signal_1096}), .c ({signal_3274, signal_1416}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1216 ( .s (enc_dec), .b ({signal_3238, signal_1030}), .a ({signal_3217, signal_1094}), .c ({signal_3331, signal_1414}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1218 ( .s (enc_dec), .b ({signal_3192, signal_1028}), .a ({signal_3161, signal_1092}), .c ({signal_3275, signal_1412}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1220 ( .s (enc_dec), .b ({signal_3237, signal_1026}), .a ({signal_3222, signal_1090}), .c ({signal_3332, signal_1410}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1222 ( .s (enc_dec), .b ({signal_3190, signal_1024}), .a ({signal_3165, signal_1088}), .c ({signal_3276, signal_1408}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1224 ( .s (enc_dec), .b ({signal_3236, signal_1022}), .a ({signal_3223, signal_1086}), .c ({signal_3333, signal_1406}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1226 ( .s (enc_dec), .b ({signal_3189, signal_1020}), .a ({signal_3167, signal_1084}), .c ({signal_3277, signal_1404}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1228 ( .s (enc_dec), .b ({signal_3235, signal_1018}), .a ({signal_3216, signal_1082}), .c ({signal_3334, signal_1402}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1230 ( .s (enc_dec), .b ({signal_3188, signal_1016}), .a ({signal_3159, signal_1080}), .c ({signal_3278, signal_1400}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1232 ( .s (enc_dec), .b ({signal_3234, signal_1014}), .a ({signal_3202, signal_1078}), .c ({signal_3335, signal_1398}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1234 ( .s (enc_dec), .b ({signal_3186, signal_1012}), .a ({signal_3146, signal_1076}), .c ({signal_3279, signal_1396}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1236 ( .s (enc_dec), .b ({signal_3233, signal_1010}), .a ({signal_3207, signal_1074}), .c ({signal_3336, signal_1394}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1238 ( .s (enc_dec), .b ({signal_3185, signal_1008}), .a ({signal_3157, signal_1072}), .c ({signal_3280, signal_1392}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1240 ( .s (enc_dec), .b ({signal_3231, signal_1006}), .a ({signal_3213, signal_1070}), .c ({signal_3337, signal_1390}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1242 ( .s (enc_dec), .b ({signal_3184, signal_1004}), .a ({signal_3163, signal_1068}), .c ({signal_3281, signal_1388}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1244 ( .s (enc_dec), .b ({signal_3230, signal_1002}), .a ({signal_3220, signal_1066}), .c ({signal_3338, signal_1386}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1246 ( .s (enc_dec), .b ({signal_3183, signal_1000}), .a ({signal_3164, signal_1064}), .c ({signal_3282, signal_1384}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1248 ( .s (enc_dec), .b ({signal_3229, signal_998}), .a ({signal_3210, signal_1062}), .c ({signal_3339, signal_1382}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1250 ( .s (enc_dec), .b ({signal_3182, signal_996}), .a ({signal_3153, signal_1060}), .c ({signal_3283, signal_1380}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1252 ( .s (enc_dec), .b ({signal_3227, signal_994}), .a ({signal_3205, signal_1058}), .c ({signal_3340, signal_1378}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1254 ( .s (enc_dec), .b ({signal_3181, signal_992}), .a ({signal_3149, signal_1056}), .c ({signal_3284, signal_1376}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1639 ( .a ({signal_2281, signal_1374}), .b ({signal_2688, signal_1744}), .clk (clk), .r (Fresh[160]), .c ({signal_2784, signal_1840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1640 ( .a ({signal_2273, signal_1370}), .b ({signal_2689, signal_1745}), .clk (clk), .r (Fresh[161]), .c ({signal_2785, signal_1841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1641 ( .a ({signal_2265, signal_1366}), .b ({signal_2690, signal_1746}), .clk (clk), .r (Fresh[162]), .c ({signal_2786, signal_1842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1642 ( .a ({signal_2257, signal_1362}), .b ({signal_2691, signal_1747}), .clk (clk), .r (Fresh[163]), .c ({signal_2787, signal_1843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1643 ( .a ({signal_2249, signal_1358}), .b ({signal_2692, signal_1748}), .clk (clk), .r (Fresh[164]), .c ({signal_2788, signal_1844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1644 ( .a ({signal_2241, signal_1354}), .b ({signal_2693, signal_1749}), .clk (clk), .r (Fresh[165]), .c ({signal_2789, signal_1845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1645 ( .a ({signal_2233, signal_1350}), .b ({signal_2694, signal_1750}), .clk (clk), .r (Fresh[166]), .c ({signal_2790, signal_1846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1646 ( .a ({signal_2225, signal_1346}), .b ({signal_2695, signal_1751}), .clk (clk), .r (Fresh[167]), .c ({signal_2791, signal_1847}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1647 ( .a ({signal_2217, signal_1342}), .b ({signal_2696, signal_1752}), .clk (clk), .r (Fresh[168]), .c ({signal_2792, signal_1848}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1648 ( .a ({signal_2209, signal_1338}), .b ({signal_2697, signal_1753}), .clk (clk), .r (Fresh[169]), .c ({signal_2793, signal_1849}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1649 ( .a ({signal_2201, signal_1334}), .b ({signal_2698, signal_1754}), .clk (clk), .r (Fresh[170]), .c ({signal_2794, signal_1850}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1650 ( .a ({signal_2193, signal_1330}), .b ({signal_2699, signal_1755}), .clk (clk), .r (Fresh[171]), .c ({signal_2795, signal_1851}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1651 ( .a ({signal_2185, signal_1326}), .b ({signal_2700, signal_1756}), .clk (clk), .r (Fresh[172]), .c ({signal_2796, signal_1852}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1652 ( .a ({signal_2177, signal_1322}), .b ({signal_2701, signal_1757}), .clk (clk), .r (Fresh[173]), .c ({signal_2797, signal_1853}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1653 ( .a ({signal_2169, signal_1318}), .b ({signal_2702, signal_1758}), .clk (clk), .r (Fresh[174]), .c ({signal_2798, signal_1854}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1654 ( .a ({signal_2161, signal_1314}), .b ({signal_2703, signal_1759}), .clk (clk), .r (Fresh[175]), .c ({signal_2799, signal_1855}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1655 ( .a ({signal_2608, signal_1664}), .b ({signal_2704, signal_1760}), .clk (clk), .r (Fresh[176]), .c ({signal_2800, signal_1856}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1656 ( .a ({signal_2611, signal_1667}), .b ({signal_2705, signal_1761}), .clk (clk), .r (Fresh[177]), .c ({signal_2801, signal_1857}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1657 ( .a ({signal_2614, signal_1670}), .b ({signal_2706, signal_1762}), .clk (clk), .r (Fresh[178]), .c ({signal_2802, signal_1858}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1658 ( .a ({signal_2617, signal_1673}), .b ({signal_2707, signal_1763}), .clk (clk), .r (Fresh[179]), .c ({signal_2803, signal_1859}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1659 ( .a ({signal_2620, signal_1676}), .b ({signal_2708, signal_1764}), .clk (clk), .r (Fresh[180]), .c ({signal_2804, signal_1860}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1660 ( .a ({signal_2623, signal_1679}), .b ({signal_2709, signal_1765}), .clk (clk), .r (Fresh[181]), .c ({signal_2805, signal_1861}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1661 ( .a ({signal_2626, signal_1682}), .b ({signal_2710, signal_1766}), .clk (clk), .r (Fresh[182]), .c ({signal_2806, signal_1862}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1662 ( .a ({signal_2629, signal_1685}), .b ({signal_2711, signal_1767}), .clk (clk), .r (Fresh[183]), .c ({signal_2807, signal_1863}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1663 ( .a ({signal_2632, signal_1688}), .b ({signal_2712, signal_1768}), .clk (clk), .r (Fresh[184]), .c ({signal_2808, signal_1864}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1664 ( .a ({signal_2635, signal_1691}), .b ({signal_2713, signal_1769}), .clk (clk), .r (Fresh[185]), .c ({signal_2809, signal_1865}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1665 ( .a ({signal_2638, signal_1694}), .b ({signal_2714, signal_1770}), .clk (clk), .r (Fresh[186]), .c ({signal_2810, signal_1866}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1666 ( .a ({signal_2641, signal_1697}), .b ({signal_2715, signal_1771}), .clk (clk), .r (Fresh[187]), .c ({signal_2811, signal_1867}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1667 ( .a ({signal_2644, signal_1700}), .b ({signal_2716, signal_1772}), .clk (clk), .r (Fresh[188]), .c ({signal_2812, signal_1868}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1668 ( .a ({signal_2647, signal_1703}), .b ({signal_2717, signal_1773}), .clk (clk), .r (Fresh[189]), .c ({signal_2813, signal_1869}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1669 ( .a ({signal_2650, signal_1706}), .b ({signal_2718, signal_1774}), .clk (clk), .r (Fresh[190]), .c ({signal_2814, signal_1870}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1670 ( .a ({signal_2653, signal_1709}), .b ({signal_2719, signal_1775}), .clk (clk), .r (Fresh[191]), .c ({signal_2815, signal_1871}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1671 ( .a ({signal_2784, signal_1840}), .b ({signal_2816, signal_1872}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1672 ( .a ({signal_2785, signal_1841}), .b ({signal_2817, signal_1873}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1673 ( .a ({signal_2786, signal_1842}), .b ({signal_2818, signal_1874}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1674 ( .a ({signal_2787, signal_1843}), .b ({signal_2819, signal_1875}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1675 ( .a ({signal_2788, signal_1844}), .b ({signal_2820, signal_1876}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1676 ( .a ({signal_2789, signal_1845}), .b ({signal_2821, signal_1877}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1677 ( .a ({signal_2790, signal_1846}), .b ({signal_2822, signal_1878}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1678 ( .a ({signal_2791, signal_1847}), .b ({signal_2823, signal_1879}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1679 ( .a ({signal_2792, signal_1848}), .b ({signal_2824, signal_1880}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1680 ( .a ({signal_2793, signal_1849}), .b ({signal_2825, signal_1881}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1681 ( .a ({signal_2794, signal_1850}), .b ({signal_2826, signal_1882}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1682 ( .a ({signal_2795, signal_1851}), .b ({signal_2827, signal_1883}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1683 ( .a ({signal_2796, signal_1852}), .b ({signal_2828, signal_1884}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1684 ( .a ({signal_2797, signal_1853}), .b ({signal_2829, signal_1885}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1685 ( .a ({signal_2798, signal_1854}), .b ({signal_2830, signal_1886}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1686 ( .a ({signal_2799, signal_1855}), .b ({signal_2831, signal_1887}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1687 ( .a ({signal_2800, signal_1856}), .b ({signal_2832, signal_1260}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1688 ( .a ({signal_2801, signal_1857}), .b ({signal_2833, signal_1264}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1689 ( .a ({signal_2802, signal_1858}), .b ({signal_2834, signal_1300}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1690 ( .a ({signal_2803, signal_1859}), .b ({signal_2835, signal_1288}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1691 ( .a ({signal_2804, signal_1860}), .b ({signal_2836, signal_1272}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1692 ( .a ({signal_2805, signal_1861}), .b ({signal_2837, signal_1252}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1693 ( .a ({signal_2806, signal_1862}), .b ({signal_2838, signal_1280}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1694 ( .a ({signal_2807, signal_1863}), .b ({signal_2839, signal_1308}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1695 ( .a ({signal_2808, signal_1864}), .b ({signal_2840, signal_1296}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1696 ( .a ({signal_2809, signal_1865}), .b ({signal_2841, signal_1292}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1697 ( .a ({signal_2810, signal_1866}), .b ({signal_2842, signal_1256}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1698 ( .a ({signal_2811, signal_1867}), .b ({signal_2843, signal_1268}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1699 ( .a ({signal_2812, signal_1868}), .b ({signal_2844, signal_1284}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1700 ( .a ({signal_2813, signal_1869}), .b ({signal_2845, signal_1304}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1701 ( .a ({signal_2814, signal_1870}), .b ({signal_2846, signal_1276}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1702 ( .a ({signal_2815, signal_1871}), .b ({signal_2847, signal_1248}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1703 ( .a ({signal_2282, signal_1518}), .b ({signal_2752, signal_1808}), .clk (clk), .r (Fresh[192]), .c ({signal_2848, signal_1888}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1704 ( .a ({signal_2274, signal_1514}), .b ({signal_2753, signal_1809}), .clk (clk), .r (Fresh[193]), .c ({signal_2849, signal_1889}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1705 ( .a ({signal_2266, signal_1510}), .b ({signal_2754, signal_1810}), .clk (clk), .r (Fresh[194]), .c ({signal_2850, signal_1890}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1706 ( .a ({signal_2258, signal_1506}), .b ({signal_2755, signal_1811}), .clk (clk), .r (Fresh[195]), .c ({signal_2851, signal_1891}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1707 ( .a ({signal_2250, signal_1502}), .b ({signal_2756, signal_1812}), .clk (clk), .r (Fresh[196]), .c ({signal_2852, signal_1892}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1708 ( .a ({signal_2242, signal_1498}), .b ({signal_2757, signal_1813}), .clk (clk), .r (Fresh[197]), .c ({signal_2853, signal_1893}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1709 ( .a ({signal_2234, signal_1494}), .b ({signal_2758, signal_1814}), .clk (clk), .r (Fresh[198]), .c ({signal_2854, signal_1894}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1710 ( .a ({signal_2226, signal_1490}), .b ({signal_2759, signal_1815}), .clk (clk), .r (Fresh[199]), .c ({signal_2855, signal_1895}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1711 ( .a ({signal_2218, signal_1486}), .b ({signal_2760, signal_1816}), .clk (clk), .r (Fresh[200]), .c ({signal_2856, signal_1896}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1712 ( .a ({signal_2210, signal_1482}), .b ({signal_2761, signal_1817}), .clk (clk), .r (Fresh[201]), .c ({signal_2857, signal_1897}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1713 ( .a ({signal_2202, signal_1478}), .b ({signal_2762, signal_1818}), .clk (clk), .r (Fresh[202]), .c ({signal_2858, signal_1898}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1714 ( .a ({signal_2194, signal_1474}), .b ({signal_2763, signal_1819}), .clk (clk), .r (Fresh[203]), .c ({signal_2859, signal_1899}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1715 ( .a ({signal_2186, signal_1470}), .b ({signal_2764, signal_1820}), .clk (clk), .r (Fresh[204]), .c ({signal_2860, signal_1900}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1716 ( .a ({signal_2178, signal_1466}), .b ({signal_2765, signal_1821}), .clk (clk), .r (Fresh[205]), .c ({signal_2861, signal_1901}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1717 ( .a ({signal_2170, signal_1462}), .b ({signal_2766, signal_1822}), .clk (clk), .r (Fresh[206]), .c ({signal_2862, signal_1902}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1718 ( .a ({signal_2162, signal_1458}), .b ({signal_2767, signal_1823}), .clk (clk), .r (Fresh[207]), .c ({signal_2863, signal_1903}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1719 ( .a ({signal_2610, signal_1666}), .b ({signal_2768, signal_1824}), .clk (clk), .r (Fresh[208]), .c ({signal_2864, signal_1904}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1720 ( .a ({signal_2613, signal_1669}), .b ({signal_2769, signal_1825}), .clk (clk), .r (Fresh[209]), .c ({signal_2865, signal_1905}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1721 ( .a ({signal_2616, signal_1672}), .b ({signal_2770, signal_1826}), .clk (clk), .r (Fresh[210]), .c ({signal_2866, signal_1906}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1722 ( .a ({signal_2619, signal_1675}), .b ({signal_2771, signal_1827}), .clk (clk), .r (Fresh[211]), .c ({signal_2867, signal_1907}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1723 ( .a ({signal_2622, signal_1678}), .b ({signal_2772, signal_1828}), .clk (clk), .r (Fresh[212]), .c ({signal_2868, signal_1908}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1724 ( .a ({signal_2625, signal_1681}), .b ({signal_2773, signal_1829}), .clk (clk), .r (Fresh[213]), .c ({signal_2869, signal_1909}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1725 ( .a ({signal_2628, signal_1684}), .b ({signal_2774, signal_1830}), .clk (clk), .r (Fresh[214]), .c ({signal_2870, signal_1910}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1726 ( .a ({signal_2631, signal_1687}), .b ({signal_2775, signal_1831}), .clk (clk), .r (Fresh[215]), .c ({signal_2871, signal_1911}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1727 ( .a ({signal_2634, signal_1690}), .b ({signal_2776, signal_1832}), .clk (clk), .r (Fresh[216]), .c ({signal_2872, signal_1912}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1728 ( .a ({signal_2637, signal_1693}), .b ({signal_2777, signal_1833}), .clk (clk), .r (Fresh[217]), .c ({signal_2873, signal_1913}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1729 ( .a ({signal_2640, signal_1696}), .b ({signal_2778, signal_1834}), .clk (clk), .r (Fresh[218]), .c ({signal_2874, signal_1914}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1730 ( .a ({signal_2643, signal_1699}), .b ({signal_2779, signal_1835}), .clk (clk), .r (Fresh[219]), .c ({signal_2875, signal_1915}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1731 ( .a ({signal_2646, signal_1702}), .b ({signal_2780, signal_1836}), .clk (clk), .r (Fresh[220]), .c ({signal_2876, signal_1916}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1732 ( .a ({signal_2649, signal_1705}), .b ({signal_2781, signal_1837}), .clk (clk), .r (Fresh[221]), .c ({signal_2877, signal_1917}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1733 ( .a ({signal_2652, signal_1708}), .b ({signal_2782, signal_1838}), .clk (clk), .r (Fresh[222]), .c ({signal_2878, signal_1918}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1734 ( .a ({signal_2655, signal_1711}), .b ({signal_2783, signal_1839}), .clk (clk), .r (Fresh[223]), .c ({signal_2879, signal_1919}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1735 ( .a ({signal_2848, signal_1888}), .b ({signal_2912, signal_1920}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1736 ( .a ({signal_2849, signal_1889}), .b ({signal_2913, signal_1921}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1737 ( .a ({signal_2850, signal_1890}), .b ({signal_2914, signal_1922}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1738 ( .a ({signal_2851, signal_1891}), .b ({signal_2915, signal_1923}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1739 ( .a ({signal_2852, signal_1892}), .b ({signal_2916, signal_1924}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1740 ( .a ({signal_2853, signal_1893}), .b ({signal_2917, signal_1925}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1741 ( .a ({signal_2854, signal_1894}), .b ({signal_2918, signal_1926}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1742 ( .a ({signal_2855, signal_1895}), .b ({signal_2919, signal_1927}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1743 ( .a ({signal_2856, signal_1896}), .b ({signal_2920, signal_1928}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1744 ( .a ({signal_2857, signal_1897}), .b ({signal_2921, signal_1929}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1745 ( .a ({signal_2858, signal_1898}), .b ({signal_2922, signal_1930}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1746 ( .a ({signal_2859, signal_1899}), .b ({signal_2923, signal_1931}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1747 ( .a ({signal_2860, signal_1900}), .b ({signal_2924, signal_1932}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1748 ( .a ({signal_2861, signal_1901}), .b ({signal_2925, signal_1933}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1749 ( .a ({signal_2862, signal_1902}), .b ({signal_2926, signal_1934}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1750 ( .a ({signal_2863, signal_1903}), .b ({signal_2927, signal_1935}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1751 ( .a ({signal_2864, signal_1904}), .b ({signal_2928, signal_1262}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1752 ( .a ({signal_2865, signal_1905}), .b ({signal_2929, signal_1266}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1753 ( .a ({signal_2866, signal_1906}), .b ({signal_2930, signal_1302}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1754 ( .a ({signal_2867, signal_1907}), .b ({signal_2931, signal_1290}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1755 ( .a ({signal_2868, signal_1908}), .b ({signal_2932, signal_1274}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1756 ( .a ({signal_2869, signal_1909}), .b ({signal_2933, signal_1254}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1757 ( .a ({signal_2870, signal_1910}), .b ({signal_2934, signal_1282}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1758 ( .a ({signal_2871, signal_1911}), .b ({signal_2935, signal_1310}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1759 ( .a ({signal_2872, signal_1912}), .b ({signal_2936, signal_1298}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1760 ( .a ({signal_2873, signal_1913}), .b ({signal_2937, signal_1294}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1761 ( .a ({signal_2874, signal_1914}), .b ({signal_2938, signal_1258}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1762 ( .a ({signal_2875, signal_1915}), .b ({signal_2939, signal_1270}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1763 ( .a ({signal_2876, signal_1916}), .b ({signal_2940, signal_1286}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1764 ( .a ({signal_2877, signal_1917}), .b ({signal_2941, signal_1306}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1765 ( .a ({signal_2878, signal_1918}), .b ({signal_2942, signal_1278}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1766 ( .a ({signal_2879, signal_1919}), .b ({signal_2943, signal_1250}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_90 ( .a ({signal_1957, signal_915}), .b ({signal_3026, signal_1303}), .c ({DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_92 ( .a ({signal_1963, signal_917}), .b ({signal_3009, signal_1265}), .c ({DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_94 ( .a ({signal_1969, signal_861}), .b ({signal_3023, signal_1249}), .c ({DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_96 ( .a ({signal_1975, signal_863}), .b ({signal_3039, signal_1251}), .c ({DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_99 ( .a ({signal_1984, signal_865}), .b ({signal_3022, signal_1277}), .c ({DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_101 ( .a ({signal_1990, signal_867}), .b ({signal_3038, signal_1279}), .c ({DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_103 ( .a ({signal_1996, signal_869}), .b ({signal_3021, signal_1305}), .c ({DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_105 ( .a ({signal_2002, signal_871}), .b ({signal_3037, signal_1307}), .c ({DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_107 ( .a ({signal_2008, signal_873}), .b ({signal_3020, signal_1285}), .c ({DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_108 ( .a ({signal_2011, signal_919}), .b ({signal_3025, signal_1267}), .c ({DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_110 ( .a ({signal_2017, signal_875}), .b ({signal_3036, signal_1287}), .c ({DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_112 ( .a ({signal_2023, signal_877}), .b ({signal_3019, signal_1269}), .c ({DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_114 ( .a ({signal_2029, signal_879}), .b ({signal_3035, signal_1271}), .c ({DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_116 ( .a ({signal_2035, signal_881}), .b ({signal_3018, signal_1257}), .c ({DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_118 ( .a ({signal_2041, signal_883}), .b ({signal_3034, signal_1259}), .c ({DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_121 ( .a ({signal_2050, signal_885}), .b ({signal_3017, signal_1293}), .c ({DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_123 ( .a ({signal_2056, signal_887}), .b ({signal_3033, signal_1295}), .c ({DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_125 ( .a ({signal_2062, signal_889}), .b ({signal_3016, signal_1297}), .c ({DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_127 ( .a ({signal_2068, signal_891}), .b ({signal_3032, signal_1299}), .c ({DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_129 ( .a ({signal_2074, signal_893}), .b ({signal_3015, signal_1309}), .c ({DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_130 ( .a ({signal_2077, signal_921}), .b ({signal_3008, signal_1261}), .c ({DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_132 ( .a ({signal_2083, signal_895}), .b ({signal_3031, signal_1311}), .c ({DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_134 ( .a ({signal_2089, signal_897}), .b ({signal_3014, signal_1281}), .c ({DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_136 ( .a ({signal_2095, signal_899}), .b ({signal_3030, signal_1283}), .c ({DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_138 ( .a ({signal_2101, signal_901}), .b ({signal_3013, signal_1253}), .c ({DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_140 ( .a ({signal_2107, signal_903}), .b ({signal_3029, signal_1255}), .c ({DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_143 ( .a ({signal_2116, signal_905}), .b ({signal_3012, signal_1273}), .c ({DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_145 ( .a ({signal_2122, signal_907}), .b ({signal_3028, signal_1275}), .c ({DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_147 ( .a ({signal_2128, signal_909}), .b ({signal_3011, signal_1289}), .c ({DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_149 ( .a ({signal_2134, signal_911}), .b ({signal_3027, signal_1291}), .c ({DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_151 ( .a ({signal_2140, signal_913}), .b ({signal_3010, signal_1301}), .c ({DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_152 ( .a ({signal_2143, signal_923}), .b ({signal_3024, signal_1263}), .c ({DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_218 ( .a ({signal_3026, signal_1303}), .b ({signal_3088, signal_286}), .c ({signal_3116, signal_1239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_220 ( .a ({signal_2542, signal_308}), .b ({signal_3009, signal_1265}), .c ({signal_3072, signal_1241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_222 ( .a ({signal_2590, signal_364}), .b ({signal_3023, signal_1249}), .c ({signal_3073, signal_1185}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_224 ( .a ({signal_3039, signal_1251}), .b ({signal_3120, signal_287}), .c ({signal_3170, signal_1187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_227 ( .a ({signal_2586, signal_360}), .b ({signal_3022, signal_1277}), .c ({signal_3074, signal_1189}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_229 ( .a ({signal_3038, signal_1279}), .b ({signal_3121, signal_288}), .c ({signal_3171, signal_1191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_231 ( .a ({signal_2582, signal_356}), .b ({signal_3021, signal_1305}), .c ({signal_3075, signal_1193}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_233 ( .a ({signal_3037, signal_1307}), .b ({signal_3122, signal_289}), .c ({signal_3172, signal_1195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({signal_2578, signal_352}), .b ({signal_3020, signal_1285}), .c ({signal_3076, signal_1197}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({signal_3025, signal_1267}), .b ({signal_3123, signal_290}), .c ({signal_3173, signal_1243}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({signal_3036, signal_1287}), .b ({signal_3232, signal_291}), .c ({signal_3285, signal_1199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({signal_2574, signal_348}), .b ({signal_3019, signal_1269}), .c ({signal_3077, signal_1201}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({signal_3035, signal_1271}), .b ({signal_3089, signal_292}), .c ({signal_3117, signal_1203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({signal_2570, signal_344}), .b ({signal_3018, signal_1257}), .c ({signal_3078, signal_1205}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({signal_3034, signal_1259}), .b ({signal_3124, signal_293}), .c ({signal_3174, signal_1207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({signal_2566, signal_340}), .b ({signal_3017, signal_1293}), .c ({signal_3079, signal_1209}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({signal_3033, signal_1295}), .b ({signal_3090, signal_294}), .c ({signal_3118, signal_1211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({signal_2562, signal_336}), .b ({signal_3016, signal_1297}), .c ({signal_3080, signal_1213}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({signal_3032, signal_1299}), .b ({signal_3125, signal_295}), .c ({signal_3175, signal_1215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .a ({signal_2558, signal_332}), .b ({signal_3015, signal_1309}), .c ({signal_3081, signal_1217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .a ({signal_2146, signal_304}), .b ({signal_3008, signal_1261}), .c ({signal_3082, signal_1245}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .a ({signal_3031, signal_1311}), .b ({signal_3191, signal_296}), .c ({signal_3225, signal_1219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({signal_2156, signal_328}), .b ({signal_3014, signal_1281}), .c ({signal_3083, signal_1221}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({signal_3030, signal_1283}), .b ({signal_3126, signal_297}), .c ({signal_3176, signal_1223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({signal_2551, signal_324}), .b ({signal_3013, signal_1253}), .c ({signal_3084, signal_1225}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .a ({signal_3029, signal_1255}), .b ({signal_3091, signal_298}), .c ({signal_3119, signal_1227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({signal_2547, signal_320}), .b ({signal_3012, signal_1273}), .c ({signal_3085, signal_1229}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({signal_3028, signal_1275}), .b ({signal_3127, signal_299}), .c ({signal_3177, signal_1231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({signal_2154, signal_316}), .b ({signal_3011, signal_1289}), .c ({signal_3086, signal_1233}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({signal_3027, signal_1291}), .b ({signal_3128, signal_300}), .c ({signal_3178, signal_1235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({signal_2151, signal_312}), .b ({signal_3010, signal_1301}), .c ({signal_3087, signal_1237}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_280 ( .a ({signal_3024, signal_1263}), .b ({signal_3129, signal_301}), .c ({signal_3179, signal_1247}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_282 ( .a ({signal_3366, signal_1111}), .b ({signal_3088, signal_286}), .c ({signal_3386, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_285 ( .a ({signal_2542, signal_308}), .b ({signal_3265, signal_1065}), .c ({signal_3286, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_287 ( .a ({signal_2590, signal_364}), .b ({signal_3255, signal_1057}), .c ({signal_3287, signal_993}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_289 ( .a ({signal_3421, signal_1059}), .b ({signal_3120, signal_287}), .c ({signal_3433, signal_995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_293 ( .a ({signal_2586, signal_360}), .b ({signal_3256, signal_1097}), .c ({signal_3288, signal_997}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_295 ( .a ({signal_3420, signal_1099}), .b ({signal_3121, signal_288}), .c ({signal_3434, signal_999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_298 ( .a ({signal_2582, signal_356}), .b ({signal_3253, signal_1077}), .c ({signal_3289, signal_1001}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_300 ( .a ({signal_3413, signal_1079}), .b ({signal_3122, signal_289}), .c ({signal_3417, signal_1003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_303 ( .a ({signal_2578, signal_352}), .b ({signal_3254, signal_1117}), .c ({signal_3290, signal_1005}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_304 ( .a ({signal_3367, signal_1067}), .b ({signal_3123, signal_290}), .c ({signal_3387, signal_1051}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_307 ( .a ({signal_3358, signal_1119}), .b ({signal_3232, signal_291}), .c ({signal_3388, signal_1007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_310 ( .a ({signal_2574, signal_348}), .b ({signal_3259, signal_1113}), .c ({signal_3291, signal_1009}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_312 ( .a ({signal_3361, signal_1115}), .b ({signal_3089, signal_292}), .c ({signal_3389, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_315 ( .a ({signal_2570, signal_344}), .b ({signal_3260, signal_1073}), .c ({signal_3292, signal_1013}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_317 ( .a ({signal_3359, signal_1075}), .b ({signal_3124, signal_293}), .c ({signal_3390, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_321 ( .a ({signal_2566, signal_340}), .b ({signal_3257, signal_1101}), .c ({signal_3293, signal_1017}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_323 ( .a ({signal_3360, signal_1103}), .b ({signal_3090, signal_294}), .c ({signal_3391, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_326 ( .a ({signal_2562, signal_336}), .b ({signal_3258, signal_1061}), .c ({signal_3294, signal_1021}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_328 ( .a ({signal_3362, signal_1063}), .b ({signal_3125, signal_295}), .c ({signal_3392, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_331 ( .a ({signal_2558, signal_332}), .b ({signal_3263, signal_1093}), .c ({signal_3295, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_332 ( .a ({signal_2146, signal_304}), .b ({signal_3266, signal_1089}), .c ({signal_3296, signal_1053}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_334 ( .a ({signal_3364, signal_1095}), .b ({signal_3191, signal_296}), .c ({signal_3393, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_337 ( .a ({signal_2156, signal_328}), .b ({signal_3264, signal_1069}), .c ({signal_3297, signal_1029}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_339 ( .a ({signal_3363, signal_1071}), .b ({signal_3126, signal_297}), .c ({signal_3394, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_342 ( .a ({signal_2551, signal_324}), .b ({signal_3261, signal_1105}), .c ({signal_3298, signal_1033}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_344 ( .a ({signal_3415, signal_1107}), .b ({signal_3091, signal_298}), .c ({signal_3418, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_348 ( .a ({signal_2547, signal_320}), .b ({signal_3262, signal_1081}), .c ({signal_3299, signal_1037}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_350 ( .a ({signal_3416, signal_1083}), .b ({signal_3127, signal_299}), .c ({signal_3419, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_353 ( .a ({signal_2154, signal_316}), .b ({signal_3267, signal_1085}), .c ({signal_3300, signal_1041}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_355 ( .a ({signal_3368, signal_1087}), .b ({signal_3128, signal_300}), .c ({signal_3395, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_358 ( .a ({signal_2151, signal_312}), .b ({signal_3268, signal_1109}), .c ({signal_3301, signal_1045}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_359 ( .a ({signal_3369, signal_1091}), .b ({signal_3129, signal_301}), .c ({signal_3396, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_535 ( .s (reset), .b ({signal_3422, signal_1439}), .a ({signal_2444, signal_991}), .c ({signal_3435, signal_460}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_541 ( .s (reset), .b ({signal_3370, signal_1437}), .a ({signal_2400, signal_989}), .c ({signal_3397, signal_464}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_547 ( .s (reset), .b ({signal_3423, signal_1435}), .a ({signal_2356, signal_987}), .c ({signal_3436, signal_468}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_553 ( .s (reset), .b ({signal_3371, signal_1433}), .a ({signal_2324, signal_985}), .c ({signal_3398, signal_472}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_559 ( .s (reset), .b ({signal_3424, signal_1431}), .a ({signal_2320, signal_983}), .c ({signal_3437, signal_476}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_565 ( .s (reset), .b ({signal_3372, signal_1429}), .a ({signal_2442, signal_981}), .c ({signal_3399, signal_480}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_571 ( .s (reset), .b ({signal_3425, signal_1427}), .a ({signal_2438, signal_979}), .c ({signal_3438, signal_484}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_577 ( .s (reset), .b ({signal_3373, signal_1425}), .a ({signal_2434, signal_977}), .c ({signal_3400, signal_488}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_583 ( .s (reset), .b ({signal_3446, signal_1423}), .a ({signal_2430, signal_975}), .c ({signal_3449, signal_492}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_589 ( .s (reset), .b ({signal_3374, signal_1421}), .a ({signal_2426, signal_973}), .c ({signal_3401, signal_496}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_595 ( .s (reset), .b ({signal_3447, signal_1419}), .a ({signal_2420, signal_971}), .c ({signal_3450, signal_500}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_601 ( .s (reset), .b ({signal_3375, signal_1417}), .a ({signal_2416, signal_969}), .c ({signal_3402, signal_504}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_607 ( .s (reset), .b ({signal_3426, signal_1415}), .a ({signal_2412, signal_967}), .c ({signal_3439, signal_508}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_613 ( .s (reset), .b ({signal_3376, signal_1413}), .a ({signal_2408, signal_965}), .c ({signal_3403, signal_512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_619 ( .s (reset), .b ({signal_3427, signal_1411}), .a ({signal_2404, signal_963}), .c ({signal_3440, signal_516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_625 ( .s (reset), .b ({signal_3377, signal_1409}), .a ({signal_2398, signal_961}), .c ({signal_3404, signal_520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_631 ( .s (reset), .b ({signal_3428, signal_1407}), .a ({signal_2394, signal_959}), .c ({signal_3441, signal_524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_637 ( .s (reset), .b ({signal_3378, signal_1405}), .a ({signal_2390, signal_957}), .c ({signal_3405, signal_528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_643 ( .s (reset), .b ({signal_3429, signal_1403}), .a ({signal_2386, signal_955}), .c ({signal_3442, signal_532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_649 ( .s (reset), .b ({signal_3379, signal_1401}), .a ({signal_2382, signal_953}), .c ({signal_3406, signal_536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_655 ( .s (reset), .b ({signal_3430, signal_1399}), .a ({signal_2376, signal_951}), .c ({signal_3443, signal_540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_661 ( .s (reset), .b ({signal_3380, signal_1397}), .a ({signal_2372, signal_949}), .c ({signal_3407, signal_544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_667 ( .s (reset), .b ({signal_3431, signal_1395}), .a ({signal_2368, signal_947}), .c ({signal_3444, signal_548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_673 ( .s (reset), .b ({signal_3381, signal_1393}), .a ({signal_2364, signal_945}), .c ({signal_3408, signal_552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_679 ( .s (reset), .b ({signal_3432, signal_1391}), .a ({signal_2360, signal_943}), .c ({signal_3445, signal_556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_685 ( .s (reset), .b ({signal_3382, signal_1389}), .a ({signal_2354, signal_941}), .c ({signal_3409, signal_560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_691 ( .s (reset), .b ({signal_3448, signal_1387}), .a ({signal_2350, signal_939}), .c ({signal_3451, signal_564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_697 ( .s (reset), .b ({signal_3383, signal_1385}), .a ({signal_2346, signal_937}), .c ({signal_3410, signal_568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_703 ( .s (reset), .b ({signal_3452, signal_1383}), .a ({signal_2342, signal_935}), .c ({signal_3454, signal_572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_709 ( .s (reset), .b ({signal_3384, signal_1381}), .a ({signal_2338, signal_933}), .c ({signal_3411, signal_576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_715 ( .s (reset), .b ({signal_3453, signal_1379}), .a ({signal_2332, signal_931}), .c ({signal_3455, signal_580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_721 ( .s (reset), .b ({signal_3385, signal_1377}), .a ({signal_2328, signal_929}), .c ({signal_3412, signal_584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1031 ( .s (enc_dec), .b ({signal_3031, signal_1311}), .a ({signal_3179, signal_1247}), .c ({signal_3243, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1033 ( .s (enc_dec), .b ({signal_3015, signal_1309}), .a ({signal_3082, signal_1245}), .c ({signal_3130, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1035 ( .s (enc_dec), .b ({signal_3037, signal_1307}), .a ({signal_3173, signal_1243}), .c ({signal_3244, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1037 ( .s (enc_dec), .b ({signal_3021, signal_1305}), .a ({signal_3072, signal_1241}), .c ({signal_3131, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1039 ( .s (enc_dec), .b ({signal_3026, signal_1303}), .a ({signal_3116, signal_1239}), .c ({signal_3197, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1041 ( .s (enc_dec), .b ({signal_3010, signal_1301}), .a ({signal_3087, signal_1237}), .c ({signal_3132, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1043 ( .s (enc_dec), .b ({signal_3032, signal_1299}), .a ({signal_3178, signal_1235}), .c ({signal_3245, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1045 ( .s (enc_dec), .b ({signal_3016, signal_1297}), .a ({signal_3086, signal_1233}), .c ({signal_3133, signal_1169}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1047 ( .s (enc_dec), .b ({signal_3033, signal_1295}), .a ({signal_3177, signal_1231}), .c ({signal_3246, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1049 ( .s (enc_dec), .b ({signal_3017, signal_1293}), .a ({signal_3085, signal_1229}), .c ({signal_3134, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1051 ( .s (enc_dec), .b ({signal_3027, signal_1291}), .a ({signal_3119, signal_1227}), .c ({signal_3198, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1053 ( .s (enc_dec), .b ({signal_3011, signal_1289}), .a ({signal_3084, signal_1225}), .c ({signal_3135, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1055 ( .s (enc_dec), .b ({signal_3036, signal_1287}), .a ({signal_3176, signal_1223}), .c ({signal_3247, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1057 ( .s (enc_dec), .b ({signal_3020, signal_1285}), .a ({signal_3083, signal_1221}), .c ({signal_3136, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1059 ( .s (enc_dec), .b ({signal_3030, signal_1283}), .a ({signal_3225, signal_1219}), .c ({signal_3318, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1061 ( .s (enc_dec), .b ({signal_3014, signal_1281}), .a ({signal_3081, signal_1217}), .c ({signal_3137, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1063 ( .s (enc_dec), .b ({signal_3038, signal_1279}), .a ({signal_3175, signal_1215}), .c ({signal_3248, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1065 ( .s (enc_dec), .b ({signal_3022, signal_1277}), .a ({signal_3080, signal_1213}), .c ({signal_3138, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1067 ( .s (enc_dec), .b ({signal_3028, signal_1275}), .a ({signal_3118, signal_1211}), .c ({signal_3199, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1069 ( .s (enc_dec), .b ({signal_3012, signal_1273}), .a ({signal_3079, signal_1209}), .c ({signal_3139, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1071 ( .s (enc_dec), .b ({signal_3035, signal_1271}), .a ({signal_3174, signal_1207}), .c ({signal_3249, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1073 ( .s (enc_dec), .b ({signal_3019, signal_1269}), .a ({signal_3078, signal_1205}), .c ({signal_3140, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1075 ( .s (enc_dec), .b ({signal_3025, signal_1267}), .a ({signal_3117, signal_1203}), .c ({signal_3200, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1077 ( .s (enc_dec), .b ({signal_3009, signal_1265}), .a ({signal_3077, signal_1201}), .c ({signal_3141, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1079 ( .s (enc_dec), .b ({signal_3024, signal_1263}), .a ({signal_3285, signal_1199}), .c ({signal_3357, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1081 ( .s (enc_dec), .b ({signal_3008, signal_1261}), .a ({signal_3076, signal_1197}), .c ({signal_3142, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1083 ( .s (enc_dec), .b ({signal_3034, signal_1259}), .a ({signal_3172, signal_1195}), .c ({signal_3250, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1085 ( .s (enc_dec), .b ({signal_3018, signal_1257}), .a ({signal_3075, signal_1193}), .c ({signal_3143, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1087 ( .s (enc_dec), .b ({signal_3029, signal_1255}), .a ({signal_3171, signal_1191}), .c ({signal_3251, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1089 ( .s (enc_dec), .b ({signal_3013, signal_1253}), .a ({signal_3074, signal_1189}), .c ({signal_3144, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1091 ( .s (enc_dec), .b ({signal_3039, signal_1251}), .a ({signal_3170, signal_1187}), .c ({signal_3252, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1093 ( .s (enc_dec), .b ({signal_3023, signal_1249}), .a ({signal_3073, signal_1185}), .c ({signal_3145, signal_1121}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .a ({signal_3252, signal_1123}), .b ({signal_3414, signal_829}), .c ({signal_3420, signal_1099}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .a ({signal_3142, signal_1133}), .b ({signal_3203, signal_831}), .c ({signal_3253, signal_1077}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .a ({signal_3357, signal_1135}), .b ({signal_3319, signal_833}), .c ({signal_3413, signal_1079}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .a ({signal_3143, signal_1129}), .b ({signal_3203, signal_831}), .c ({signal_3254, signal_1117}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .a ({signal_3145, signal_1121}), .b ({signal_3144, signal_1125}), .c ({signal_3203, signal_831}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1108 ( .a ({signal_3144, signal_1125}), .b ({signal_3206, signal_835}), .c ({signal_3255, signal_1057}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1111 ( .a ({signal_3251, signal_1127}), .b ({signal_3414, signal_829}), .c ({signal_3421, signal_1059}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1112 ( .a ({signal_3250, signal_1131}), .b ({signal_3357, signal_1135}), .c ({signal_3414, signal_829}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1115 ( .a ({signal_3145, signal_1121}), .b ({signal_3206, signal_835}), .c ({signal_3256, signal_1097}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1116 ( .a ({signal_3142, signal_1133}), .b ({signal_3143, signal_1129}), .c ({signal_3206, signal_835}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1117 ( .a ({signal_3250, signal_1131}), .b ({signal_3319, signal_833}), .c ({signal_3358, signal_1119}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1118 ( .a ({signal_3252, signal_1123}), .b ({signal_3251, signal_1127}), .c ({signal_3319, signal_833}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1120 ( .a ({signal_3200, signal_1139}), .b ({signal_3320, signal_837}), .c ({signal_3359, signal_1075}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1122 ( .a ({signal_3138, signal_1149}), .b ({signal_3209, signal_839}), .c ({signal_3257, signal_1101}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1124 ( .a ({signal_3248, signal_1151}), .b ({signal_3321, signal_841}), .c ({signal_3360, signal_1103}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1127 ( .a ({signal_3139, signal_1145}), .b ({signal_3209, signal_839}), .c ({signal_3258, signal_1061}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1128 ( .a ({signal_3141, signal_1137}), .b ({signal_3140, signal_1141}), .c ({signal_3209, signal_839}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1132 ( .a ({signal_3140, signal_1141}), .b ({signal_3212, signal_843}), .c ({signal_3259, signal_1113}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1135 ( .a ({signal_3249, signal_1143}), .b ({signal_3320, signal_837}), .c ({signal_3361, signal_1115}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1136 ( .a ({signal_3199, signal_1147}), .b ({signal_3248, signal_1151}), .c ({signal_3320, signal_837}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .a ({signal_3141, signal_1137}), .b ({signal_3212, signal_843}), .c ({signal_3260, signal_1073}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .a ({signal_3138, signal_1149}), .b ({signal_3139, signal_1145}), .c ({signal_3212, signal_843}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .a ({signal_3199, signal_1147}), .b ({signal_3321, signal_841}), .c ({signal_3362, signal_1063}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .a ({signal_3200, signal_1139}), .b ({signal_3249, signal_1143}), .c ({signal_3321, signal_841}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .a ({signal_3318, signal_1155}), .b ({signal_3322, signal_845}), .c ({signal_3363, signal_1071}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .a ({signal_3134, signal_1165}), .b ({signal_3215, signal_847}), .c ({signal_3261, signal_1105}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .a ({signal_3246, signal_1167}), .b ({signal_3365, signal_849}), .c ({signal_3415, signal_1107}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .a ({signal_3135, signal_1161}), .b ({signal_3215, signal_847}), .c ({signal_3262, signal_1081}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .a ({signal_3137, signal_1153}), .b ({signal_3136, signal_1157}), .c ({signal_3215, signal_847}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .a ({signal_3136, signal_1157}), .b ({signal_3218, signal_851}), .c ({signal_3263, signal_1093}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .a ({signal_3247, signal_1159}), .b ({signal_3322, signal_845}), .c ({signal_3364, signal_1095}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .a ({signal_3198, signal_1163}), .b ({signal_3246, signal_1167}), .c ({signal_3322, signal_845}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .a ({signal_3137, signal_1153}), .b ({signal_3218, signal_851}), .c ({signal_3264, signal_1069}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .a ({signal_3134, signal_1165}), .b ({signal_3135, signal_1161}), .c ({signal_3218, signal_851}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .a ({signal_3198, signal_1163}), .b ({signal_3365, signal_849}), .c ({signal_3416, signal_1083}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .a ({signal_3318, signal_1155}), .b ({signal_3247, signal_1159}), .c ({signal_3365, signal_849}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .a ({signal_3245, signal_1171}), .b ({signal_3323, signal_853}), .c ({signal_3366, signal_1111}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .a ({signal_3130, signal_1181}), .b ({signal_3221, signal_855}), .c ({signal_3265, signal_1065}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .a ({signal_3243, signal_1183}), .b ({signal_3324, signal_857}), .c ({signal_3367, signal_1067}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .a ({signal_3131, signal_1177}), .b ({signal_3221, signal_855}), .c ({signal_3266, signal_1089}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .a ({signal_3133, signal_1169}), .b ({signal_3132, signal_1173}), .c ({signal_3221, signal_855}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .a ({signal_3132, signal_1173}), .b ({signal_3224, signal_859}), .c ({signal_3267, signal_1085}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .a ({signal_3197, signal_1175}), .b ({signal_3323, signal_853}), .c ({signal_3368, signal_1087}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .a ({signal_3244, signal_1179}), .b ({signal_3243, signal_1183}), .c ({signal_3323, signal_853}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .a ({signal_3133, signal_1169}), .b ({signal_3224, signal_859}), .c ({signal_3268, signal_1109}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .a ({signal_3130, signal_1181}), .b ({signal_3131, signal_1177}), .c ({signal_3224, signal_859}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .a ({signal_3244, signal_1179}), .b ({signal_3324, signal_857}), .c ({signal_3369, signal_1091}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .a ({signal_3245, signal_1171}), .b ({signal_3197, signal_1175}), .c ({signal_3324, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1191 ( .s (enc_dec), .b ({signal_3396, signal_1055}), .a ({signal_3358, signal_1119}), .c ({signal_3422, signal_1439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1193 ( .s (enc_dec), .b ({signal_3296, signal_1053}), .a ({signal_3254, signal_1117}), .c ({signal_3370, signal_1437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1195 ( .s (enc_dec), .b ({signal_3387, signal_1051}), .a ({signal_3361, signal_1115}), .c ({signal_3423, signal_1435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1197 ( .s (enc_dec), .b ({signal_3286, signal_1049}), .a ({signal_3259, signal_1113}), .c ({signal_3371, signal_1433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1199 ( .s (enc_dec), .b ({signal_3386, signal_1047}), .a ({signal_3366, signal_1111}), .c ({signal_3424, signal_1431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1201 ( .s (enc_dec), .b ({signal_3301, signal_1045}), .a ({signal_3268, signal_1109}), .c ({signal_3372, signal_1429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1203 ( .s (enc_dec), .b ({signal_3395, signal_1043}), .a ({signal_3415, signal_1107}), .c ({signal_3425, signal_1427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1205 ( .s (enc_dec), .b ({signal_3300, signal_1041}), .a ({signal_3261, signal_1105}), .c ({signal_3373, signal_1425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1207 ( .s (enc_dec), .b ({signal_3419, signal_1039}), .a ({signal_3360, signal_1103}), .c ({signal_3446, signal_1423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1209 ( .s (enc_dec), .b ({signal_3299, signal_1037}), .a ({signal_3257, signal_1101}), .c ({signal_3374, signal_1421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1211 ( .s (enc_dec), .b ({signal_3418, signal_1035}), .a ({signal_3420, signal_1099}), .c ({signal_3447, signal_1419}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1213 ( .s (enc_dec), .b ({signal_3298, signal_1033}), .a ({signal_3256, signal_1097}), .c ({signal_3375, signal_1417}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1215 ( .s (enc_dec), .b ({signal_3394, signal_1031}), .a ({signal_3364, signal_1095}), .c ({signal_3426, signal_1415}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1217 ( .s (enc_dec), .b ({signal_3297, signal_1029}), .a ({signal_3263, signal_1093}), .c ({signal_3376, signal_1413}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1219 ( .s (enc_dec), .b ({signal_3393, signal_1027}), .a ({signal_3369, signal_1091}), .c ({signal_3427, signal_1411}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1221 ( .s (enc_dec), .b ({signal_3295, signal_1025}), .a ({signal_3266, signal_1089}), .c ({signal_3377, signal_1409}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1223 ( .s (enc_dec), .b ({signal_3392, signal_1023}), .a ({signal_3368, signal_1087}), .c ({signal_3428, signal_1407}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1225 ( .s (enc_dec), .b ({signal_3294, signal_1021}), .a ({signal_3267, signal_1085}), .c ({signal_3378, signal_1405}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1227 ( .s (enc_dec), .b ({signal_3391, signal_1019}), .a ({signal_3416, signal_1083}), .c ({signal_3429, signal_1403}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1229 ( .s (enc_dec), .b ({signal_3293, signal_1017}), .a ({signal_3262, signal_1081}), .c ({signal_3379, signal_1401}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1231 ( .s (enc_dec), .b ({signal_3390, signal_1015}), .a ({signal_3413, signal_1079}), .c ({signal_3430, signal_1399}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1233 ( .s (enc_dec), .b ({signal_3292, signal_1013}), .a ({signal_3253, signal_1077}), .c ({signal_3380, signal_1397}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1235 ( .s (enc_dec), .b ({signal_3389, signal_1011}), .a ({signal_3359, signal_1075}), .c ({signal_3431, signal_1395}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1237 ( .s (enc_dec), .b ({signal_3291, signal_1009}), .a ({signal_3260, signal_1073}), .c ({signal_3381, signal_1393}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1239 ( .s (enc_dec), .b ({signal_3388, signal_1007}), .a ({signal_3363, signal_1071}), .c ({signal_3432, signal_1391}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1241 ( .s (enc_dec), .b ({signal_3290, signal_1005}), .a ({signal_3264, signal_1069}), .c ({signal_3382, signal_1389}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1243 ( .s (enc_dec), .b ({signal_3417, signal_1003}), .a ({signal_3367, signal_1067}), .c ({signal_3448, signal_1387}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1245 ( .s (enc_dec), .b ({signal_3289, signal_1001}), .a ({signal_3265, signal_1065}), .c ({signal_3383, signal_1385}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1247 ( .s (enc_dec), .b ({signal_3434, signal_999}), .a ({signal_3362, signal_1063}), .c ({signal_3452, signal_1383}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1249 ( .s (enc_dec), .b ({signal_3288, signal_997}), .a ({signal_3258, signal_1061}), .c ({signal_3384, signal_1381}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1251 ( .s (enc_dec), .b ({signal_3433, signal_995}), .a ({signal_3421, signal_1059}), .c ({signal_3453, signal_1379}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1253 ( .s (enc_dec), .b ({signal_3287, signal_993}), .a ({signal_3255, signal_1057}), .c ({signal_3385, signal_1377}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1767 ( .a ({signal_2608, signal_1664}), .b ({signal_2816, signal_1872}), .clk (clk), .r (Fresh[224]), .c ({signal_2944, signal_1936}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1768 ( .a ({signal_2611, signal_1667}), .b ({signal_2817, signal_1873}), .clk (clk), .r (Fresh[225]), .c ({signal_2945, signal_1937}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1769 ( .a ({signal_2614, signal_1670}), .b ({signal_2818, signal_1874}), .clk (clk), .r (Fresh[226]), .c ({signal_2946, signal_1938}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1770 ( .a ({signal_2617, signal_1673}), .b ({signal_2819, signal_1875}), .clk (clk), .r (Fresh[227]), .c ({signal_2947, signal_1939}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1771 ( .a ({signal_2620, signal_1676}), .b ({signal_2820, signal_1876}), .clk (clk), .r (Fresh[228]), .c ({signal_2948, signal_1940}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1772 ( .a ({signal_2623, signal_1679}), .b ({signal_2821, signal_1877}), .clk (clk), .r (Fresh[229]), .c ({signal_2949, signal_1941}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1773 ( .a ({signal_2626, signal_1682}), .b ({signal_2822, signal_1878}), .clk (clk), .r (Fresh[230]), .c ({signal_2950, signal_1942}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1774 ( .a ({signal_2629, signal_1685}), .b ({signal_2823, signal_1879}), .clk (clk), .r (Fresh[231]), .c ({signal_2951, signal_1943}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1775 ( .a ({signal_2632, signal_1688}), .b ({signal_2824, signal_1880}), .clk (clk), .r (Fresh[232]), .c ({signal_2952, signal_1944}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1776 ( .a ({signal_2635, signal_1691}), .b ({signal_2825, signal_1881}), .clk (clk), .r (Fresh[233]), .c ({signal_2953, signal_1945}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1777 ( .a ({signal_2638, signal_1694}), .b ({signal_2826, signal_1882}), .clk (clk), .r (Fresh[234]), .c ({signal_2954, signal_1946}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1778 ( .a ({signal_2641, signal_1697}), .b ({signal_2827, signal_1883}), .clk (clk), .r (Fresh[235]), .c ({signal_2955, signal_1947}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1779 ( .a ({signal_2644, signal_1700}), .b ({signal_2828, signal_1884}), .clk (clk), .r (Fresh[236]), .c ({signal_2956, signal_1948}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1780 ( .a ({signal_2647, signal_1703}), .b ({signal_2829, signal_1885}), .clk (clk), .r (Fresh[237]), .c ({signal_2957, signal_1949}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1781 ( .a ({signal_2650, signal_1706}), .b ({signal_2830, signal_1886}), .clk (clk), .r (Fresh[238]), .c ({signal_2958, signal_1950}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1782 ( .a ({signal_2653, signal_1709}), .b ({signal_2831, signal_1887}), .clk (clk), .r (Fresh[239]), .c ({signal_2959, signal_1951}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1783 ( .a ({signal_2944, signal_1936}), .b ({signal_3008, signal_1261}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1784 ( .a ({signal_2945, signal_1937}), .b ({signal_3009, signal_1265}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1785 ( .a ({signal_2946, signal_1938}), .b ({signal_3010, signal_1301}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1786 ( .a ({signal_2947, signal_1939}), .b ({signal_3011, signal_1289}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1787 ( .a ({signal_2948, signal_1940}), .b ({signal_3012, signal_1273}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1788 ( .a ({signal_2949, signal_1941}), .b ({signal_3013, signal_1253}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1789 ( .a ({signal_2950, signal_1942}), .b ({signal_3014, signal_1281}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1790 ( .a ({signal_2951, signal_1943}), .b ({signal_3015, signal_1309}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1791 ( .a ({signal_2952, signal_1944}), .b ({signal_3016, signal_1297}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1792 ( .a ({signal_2953, signal_1945}), .b ({signal_3017, signal_1293}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1793 ( .a ({signal_2954, signal_1946}), .b ({signal_3018, signal_1257}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1794 ( .a ({signal_2955, signal_1947}), .b ({signal_3019, signal_1269}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1795 ( .a ({signal_2956, signal_1948}), .b ({signal_3020, signal_1285}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1796 ( .a ({signal_2957, signal_1949}), .b ({signal_3021, signal_1305}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1797 ( .a ({signal_2958, signal_1950}), .b ({signal_3022, signal_1277}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1798 ( .a ({signal_2959, signal_1951}), .b ({signal_3023, signal_1249}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1799 ( .a ({signal_2461, signal_1568}), .b ({signal_2912, signal_1920}), .clk (clk), .r (Fresh[240]), .c ({signal_3024, signal_1263}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1800 ( .a ({signal_2462, signal_1569}), .b ({signal_2913, signal_1921}), .clk (clk), .r (Fresh[241]), .c ({signal_3025, signal_1267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1801 ( .a ({signal_2463, signal_1570}), .b ({signal_2914, signal_1922}), .clk (clk), .r (Fresh[242]), .c ({signal_3026, signal_1303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1802 ( .a ({signal_2464, signal_1571}), .b ({signal_2915, signal_1923}), .clk (clk), .r (Fresh[243]), .c ({signal_3027, signal_1291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1803 ( .a ({signal_2465, signal_1572}), .b ({signal_2916, signal_1924}), .clk (clk), .r (Fresh[244]), .c ({signal_3028, signal_1275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1804 ( .a ({signal_2466, signal_1573}), .b ({signal_2917, signal_1925}), .clk (clk), .r (Fresh[245]), .c ({signal_3029, signal_1255}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1805 ( .a ({signal_2467, signal_1574}), .b ({signal_2918, signal_1926}), .clk (clk), .r (Fresh[246]), .c ({signal_3030, signal_1283}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1806 ( .a ({signal_2468, signal_1575}), .b ({signal_2919, signal_1927}), .clk (clk), .r (Fresh[247]), .c ({signal_3031, signal_1311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1807 ( .a ({signal_2469, signal_1576}), .b ({signal_2920, signal_1928}), .clk (clk), .r (Fresh[248]), .c ({signal_3032, signal_1299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1808 ( .a ({signal_2470, signal_1577}), .b ({signal_2921, signal_1929}), .clk (clk), .r (Fresh[249]), .c ({signal_3033, signal_1295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1809 ( .a ({signal_2471, signal_1578}), .b ({signal_2922, signal_1930}), .clk (clk), .r (Fresh[250]), .c ({signal_3034, signal_1259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1810 ( .a ({signal_2472, signal_1579}), .b ({signal_2923, signal_1931}), .clk (clk), .r (Fresh[251]), .c ({signal_3035, signal_1271}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1811 ( .a ({signal_2473, signal_1580}), .b ({signal_2924, signal_1932}), .clk (clk), .r (Fresh[252]), .c ({signal_3036, signal_1287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1812 ( .a ({signal_2474, signal_1581}), .b ({signal_2925, signal_1933}), .clk (clk), .r (Fresh[253]), .c ({signal_3037, signal_1307}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1813 ( .a ({signal_2475, signal_1582}), .b ({signal_2926, signal_1934}), .clk (clk), .r (Fresh[254]), .c ({signal_3038, signal_1279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1814 ( .a ({signal_2476, signal_1583}), .b ({signal_2927, signal_1935}), .clk (clk), .r (Fresh[255]), .c ({signal_3039, signal_1251}) ) ;

    /* register cells */
    DFF_X1 cell_82 ( .CK (signal_3712), .D (signal_283), .Q (signal_927), .QN () ) ;
    DFF_X1 cell_84 ( .CK (signal_3712), .D (signal_282), .Q (signal_926), .QN () ) ;
    DFF_X1 cell_86 ( .CK (signal_3712), .D (signal_278), .Q (signal_925), .QN () ) ;
    DFF_X1 cell_88 ( .CK (signal_3712), .D (signal_280), .Q (signal_924), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_537 ( .clk (signal_3712), .D ({signal_3435, signal_460}), .Q ({signal_2283, signal_1375}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_540 ( .clk (signal_3712), .D ({signal_3341, signal_462}), .Q ({signal_2281, signal_1374}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_543 ( .clk (signal_3712), .D ({signal_3397, signal_464}), .Q ({signal_2279, signal_1373}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_546 ( .clk (signal_3712), .D ({signal_3302, signal_466}), .Q ({signal_2277, signal_1372}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_549 ( .clk (signal_3712), .D ({signal_3436, signal_468}), .Q ({signal_2275, signal_1371}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_552 ( .clk (signal_3712), .D ({signal_3342, signal_470}), .Q ({signal_2273, signal_1370}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_555 ( .clk (signal_3712), .D ({signal_3398, signal_472}), .Q ({signal_2271, signal_1369}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_558 ( .clk (signal_3712), .D ({signal_3303, signal_474}), .Q ({signal_2269, signal_1368}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_561 ( .clk (signal_3712), .D ({signal_3437, signal_476}), .Q ({signal_2267, signal_1367}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_564 ( .clk (signal_3712), .D ({signal_3343, signal_478}), .Q ({signal_2265, signal_1366}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_567 ( .clk (signal_3712), .D ({signal_3399, signal_480}), .Q ({signal_2263, signal_1365}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_570 ( .clk (signal_3712), .D ({signal_3304, signal_482}), .Q ({signal_2261, signal_1364}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_573 ( .clk (signal_3712), .D ({signal_3438, signal_484}), .Q ({signal_2259, signal_1363}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_576 ( .clk (signal_3712), .D ({signal_3344, signal_486}), .Q ({signal_2257, signal_1362}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_579 ( .clk (signal_3712), .D ({signal_3400, signal_488}), .Q ({signal_2255, signal_1361}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_582 ( .clk (signal_3712), .D ({signal_3305, signal_490}), .Q ({signal_2253, signal_1360}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_585 ( .clk (signal_3712), .D ({signal_3449, signal_492}), .Q ({signal_2251, signal_1359}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_588 ( .clk (signal_3712), .D ({signal_3345, signal_494}), .Q ({signal_2249, signal_1358}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_591 ( .clk (signal_3712), .D ({signal_3401, signal_496}), .Q ({signal_2247, signal_1357}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_594 ( .clk (signal_3712), .D ({signal_3306, signal_498}), .Q ({signal_2245, signal_1356}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_597 ( .clk (signal_3712), .D ({signal_3450, signal_500}), .Q ({signal_2243, signal_1355}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_600 ( .clk (signal_3712), .D ({signal_3346, signal_502}), .Q ({signal_2241, signal_1354}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_603 ( .clk (signal_3712), .D ({signal_3402, signal_504}), .Q ({signal_2239, signal_1353}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_606 ( .clk (signal_3712), .D ({signal_3307, signal_506}), .Q ({signal_2237, signal_1352}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_609 ( .clk (signal_3712), .D ({signal_3439, signal_508}), .Q ({signal_2235, signal_1351}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_612 ( .clk (signal_3712), .D ({signal_3347, signal_510}), .Q ({signal_2233, signal_1350}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_615 ( .clk (signal_3712), .D ({signal_3403, signal_512}), .Q ({signal_2231, signal_1349}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_618 ( .clk (signal_3712), .D ({signal_3308, signal_514}), .Q ({signal_2229, signal_1348}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_621 ( .clk (signal_3712), .D ({signal_3440, signal_516}), .Q ({signal_2227, signal_1347}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_624 ( .clk (signal_3712), .D ({signal_3348, signal_518}), .Q ({signal_2225, signal_1346}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_627 ( .clk (signal_3712), .D ({signal_3404, signal_520}), .Q ({signal_2223, signal_1345}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_630 ( .clk (signal_3712), .D ({signal_3309, signal_522}), .Q ({signal_2221, signal_1344}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_633 ( .clk (signal_3712), .D ({signal_3441, signal_524}), .Q ({signal_2219, signal_1343}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_636 ( .clk (signal_3712), .D ({signal_3349, signal_526}), .Q ({signal_2217, signal_1342}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_639 ( .clk (signal_3712), .D ({signal_3405, signal_528}), .Q ({signal_2215, signal_1341}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_642 ( .clk (signal_3712), .D ({signal_3310, signal_530}), .Q ({signal_2213, signal_1340}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_645 ( .clk (signal_3712), .D ({signal_3442, signal_532}), .Q ({signal_2211, signal_1339}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_648 ( .clk (signal_3712), .D ({signal_3350, signal_534}), .Q ({signal_2209, signal_1338}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_651 ( .clk (signal_3712), .D ({signal_3406, signal_536}), .Q ({signal_2207, signal_1337}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_654 ( .clk (signal_3712), .D ({signal_3311, signal_538}), .Q ({signal_2205, signal_1336}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_657 ( .clk (signal_3712), .D ({signal_3443, signal_540}), .Q ({signal_2203, signal_1335}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_660 ( .clk (signal_3712), .D ({signal_3351, signal_542}), .Q ({signal_2201, signal_1334}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_663 ( .clk (signal_3712), .D ({signal_3407, signal_544}), .Q ({signal_2199, signal_1333}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_666 ( .clk (signal_3712), .D ({signal_3312, signal_546}), .Q ({signal_2197, signal_1332}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_669 ( .clk (signal_3712), .D ({signal_3444, signal_548}), .Q ({signal_2195, signal_1331}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_672 ( .clk (signal_3712), .D ({signal_3352, signal_550}), .Q ({signal_2193, signal_1330}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_675 ( .clk (signal_3712), .D ({signal_3408, signal_552}), .Q ({signal_2191, signal_1329}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_678 ( .clk (signal_3712), .D ({signal_3313, signal_554}), .Q ({signal_2189, signal_1328}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_681 ( .clk (signal_3712), .D ({signal_3445, signal_556}), .Q ({signal_2187, signal_1327}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_684 ( .clk (signal_3712), .D ({signal_3353, signal_558}), .Q ({signal_2185, signal_1326}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_687 ( .clk (signal_3712), .D ({signal_3409, signal_560}), .Q ({signal_2183, signal_1325}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_690 ( .clk (signal_3712), .D ({signal_3314, signal_562}), .Q ({signal_2181, signal_1324}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_693 ( .clk (signal_3712), .D ({signal_3451, signal_564}), .Q ({signal_2179, signal_1323}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_696 ( .clk (signal_3712), .D ({signal_3354, signal_566}), .Q ({signal_2177, signal_1322}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_699 ( .clk (signal_3712), .D ({signal_3410, signal_568}), .Q ({signal_2175, signal_1321}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_702 ( .clk (signal_3712), .D ({signal_3315, signal_570}), .Q ({signal_2173, signal_1320}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_705 ( .clk (signal_3712), .D ({signal_3454, signal_572}), .Q ({signal_2171, signal_1319}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_708 ( .clk (signal_3712), .D ({signal_3355, signal_574}), .Q ({signal_2169, signal_1318}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_711 ( .clk (signal_3712), .D ({signal_3411, signal_576}), .Q ({signal_2167, signal_1317}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_714 ( .clk (signal_3712), .D ({signal_3316, signal_578}), .Q ({signal_2165, signal_1316}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_717 ( .clk (signal_3712), .D ({signal_3455, signal_580}), .Q ({signal_2163, signal_1315}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_720 ( .clk (signal_3712), .D ({signal_3356, signal_582}), .Q ({signal_2161, signal_1314}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_723 ( .clk (signal_3712), .D ({signal_3412, signal_584}), .Q ({signal_2159, signal_1313}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_726 ( .clk (signal_3712), .D ({signal_3317, signal_586}), .Q ({signal_2157, signal_1312}) ) ;
endmodule
