/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_Pipeline_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input [399:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    wire sbe_n10 ;
    wire sbe_n9 ;
    wire sbe_n8 ;
    wire sbe_n7 ;
    wire sbe_n6 ;
    wire sbe_n5 ;
    wire sbe_n4 ;
    wire sbe_n3 ;
    wire sbe_n12 ;
    wire sbe_n11 ;
    wire sbe_n2 ;
    wire sbe_n1 ;
    wire sbe_n25 ;
    wire sbe_n24 ;
    wire sbe_n23 ;
    wire sbe_n22 ;
    wire sbe_n21 ;
    wire sbe_n20 ;
    wire sbe_n19 ;
    wire sbe_n18 ;
    wire sbe_n17 ;
    wire sbe_n16 ;
    wire sbe_n15 ;
    wire sbe_n14 ;
    wire sbe_D_0_ ;
    wire sbe_D_2_ ;
    wire sbe_D_3_ ;
    wire sbe_D_5_ ;
    wire sbe_D_6_ ;
    wire sbe_C_0_ ;
    wire sbe_C_1_ ;
    wire sbe_C_2_ ;
    wire sbe_C_3_ ;
    wire sbe_C_4_ ;
    wire sbe_C_5_ ;
    wire sbe_C_6_ ;
    wire sbe_C_7_ ;
    wire sbe_Y_0_ ;
    wire sbe_Y_1_ ;
    wire sbe_Y_2_ ;
    wire sbe_Y_4_ ;
    wire sbe_Y_5_ ;
    wire sbe_Y_6_ ;
    wire sbe_B_3_ ;
    wire sbe_B_6_ ;
    wire sbe_sel_in_m7_n8 ;
    wire sbe_sel_in_m6_n8 ;
    wire sbe_sel_in_m5_n8 ;
    wire sbe_sel_in_m4_n8 ;
    wire sbe_sel_in_m3_n8 ;
    wire sbe_sel_in_m2_n8 ;
    wire sbe_sel_in_m1_n8 ;
    wire sbe_sel_in_m0_n8 ;
    wire sbe_inv_n21 ;
    wire sbe_inv_n20 ;
    wire sbe_inv_n19 ;
    wire sbe_inv_n18 ;
    wire sbe_inv_n17 ;
    wire sbe_inv_n16 ;
    wire sbe_inv_n15 ;
    wire sbe_inv_n14 ;
    wire sbe_inv_n13 ;
    wire sbe_inv_n12 ;
    wire sbe_inv_n11 ;
    wire sbe_inv_n10 ;
    wire sbe_inv_n9 ;
    wire sbe_inv_n8 ;
    wire sbe_inv_n7 ;
    wire sbe_inv_n6 ;
    wire sbe_inv_n5 ;
    wire sbe_inv_n4 ;
    wire sbe_inv_n3 ;
    wire sbe_inv_n2 ;
    wire sbe_inv_dd ;
    wire sbe_inv_dh ;
    wire sbe_inv_dl ;
    wire sbe_inv_sd_0_ ;
    wire sbe_inv_sd_1_ ;
    wire sbe_inv_d_0_ ;
    wire sbe_inv_d_1_ ;
    wire sbe_inv_d_2_ ;
    wire sbe_inv_d_3_ ;
    wire sbe_inv_bb ;
    wire sbe_inv_bh ;
    wire sbe_inv_bl ;
    wire sbe_inv_aa ;
    wire sbe_inv_ah ;
    wire sbe_inv_al ;
    wire sbe_inv_sb_0_ ;
    wire sbe_inv_sb_1_ ;
    wire sbe_inv_sa_0_ ;
    wire sbe_inv_sa_1_ ;
    wire sbe_inv_dinv_n4 ;
    wire sbe_inv_dinv_n3 ;
    wire sbe_inv_dinv_n2 ;
    wire sbe_inv_dinv_n1 ;
    wire sbe_inv_dinv_sd ;
    wire sbe_inv_dinv_d_0_ ;
    wire sbe_inv_dinv_d_1_ ;
    wire sbe_inv_dinv_sb ;
    wire sbe_inv_dinv_sa ;
    wire sbe_inv_dinv_pmul_n9 ;
    wire sbe_inv_dinv_pmul_n8 ;
    wire sbe_inv_dinv_pmul_n7 ;
    wire sbe_inv_dinv_qmul_n9 ;
    wire sbe_inv_dinv_qmul_n8 ;
    wire sbe_inv_dinv_qmul_n7 ;
    wire sbe_inv_pmul_p_0_ ;
    wire sbe_inv_pmul_p_1_ ;
    wire sbe_inv_pmul_himul_n9 ;
    wire sbe_inv_pmul_himul_n8 ;
    wire sbe_inv_pmul_himul_n7 ;
    wire sbe_inv_pmul_lomul_n9 ;
    wire sbe_inv_pmul_lomul_n8 ;
    wire sbe_inv_pmul_lomul_n7 ;
    wire sbe_inv_pmul_summul_n9 ;
    wire sbe_inv_pmul_summul_n8 ;
    wire sbe_inv_pmul_summul_n7 ;
    wire sbe_inv_qmul_p_0_ ;
    wire sbe_inv_qmul_p_1_ ;
    wire sbe_inv_qmul_himul_n9 ;
    wire sbe_inv_qmul_himul_n8 ;
    wire sbe_inv_qmul_himul_n7 ;
    wire sbe_inv_qmul_lomul_n9 ;
    wire sbe_inv_qmul_lomul_n8 ;
    wire sbe_inv_qmul_lomul_n7 ;
    wire sbe_inv_qmul_summul_n9 ;
    wire sbe_inv_qmul_summul_n8 ;
    wire sbe_inv_qmul_summul_n7 ;
    wire sbe_sel_out_m7_n8 ;
    wire sbe_sel_out_m6_n8 ;
    wire sbe_sel_out_m5_n8 ;
    wire sbe_sel_out_m4_n8 ;
    wire sbe_sel_out_m3_n8 ;
    wire sbe_sel_out_m2_n8 ;
    wire sbe_sel_out_m1_n8 ;
    wire sbe_sel_out_m0_n8 ;
    wire [7:0] O ;
    wire [6:3] sbe_X ;
    wire [7:0] sbe_Z ;
    wire [3:0] sbe_inv_c ;
    wire [1:0] sbe_inv_pmul_pl ;
    wire [1:0] sbe_inv_pmul_ph ;
    wire [1:0] sbe_inv_qmul_pl ;
    wire [1:0] sbe_inv_qmul_ph ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;
    wire new_AGEMA_signal_593 ;
    wire new_AGEMA_signal_594 ;
    wire new_AGEMA_signal_595 ;
    wire new_AGEMA_signal_596 ;
    wire new_AGEMA_signal_597 ;
    wire new_AGEMA_signal_598 ;
    wire new_AGEMA_signal_599 ;
    wire new_AGEMA_signal_600 ;
    wire new_AGEMA_signal_601 ;
    wire new_AGEMA_signal_602 ;
    wire new_AGEMA_signal_603 ;
    wire new_AGEMA_signal_604 ;
    wire new_AGEMA_signal_605 ;
    wire new_AGEMA_signal_606 ;
    wire new_AGEMA_signal_607 ;
    wire new_AGEMA_signal_608 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;
    wire new_AGEMA_signal_656 ;
    wire new_AGEMA_signal_657 ;
    wire new_AGEMA_signal_658 ;
    wire new_AGEMA_signal_659 ;
    wire new_AGEMA_signal_660 ;
    wire new_AGEMA_signal_661 ;
    wire new_AGEMA_signal_662 ;
    wire new_AGEMA_signal_663 ;
    wire new_AGEMA_signal_664 ;
    wire new_AGEMA_signal_665 ;
    wire new_AGEMA_signal_666 ;
    wire new_AGEMA_signal_667 ;
    wire new_AGEMA_signal_668 ;
    wire new_AGEMA_signal_669 ;
    wire new_AGEMA_signal_670 ;
    wire new_AGEMA_signal_671 ;
    wire new_AGEMA_signal_672 ;
    wire new_AGEMA_signal_673 ;
    wire new_AGEMA_signal_674 ;
    wire new_AGEMA_signal_675 ;
    wire new_AGEMA_signal_676 ;
    wire new_AGEMA_signal_677 ;
    wire new_AGEMA_signal_678 ;
    wire new_AGEMA_signal_679 ;
    wire new_AGEMA_signal_680 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_699 ;
    wire new_AGEMA_signal_700 ;
    wire new_AGEMA_signal_701 ;
    wire new_AGEMA_signal_702 ;
    wire new_AGEMA_signal_703 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_709 ;
    wire new_AGEMA_signal_710 ;
    wire new_AGEMA_signal_711 ;
    wire new_AGEMA_signal_712 ;
    wire new_AGEMA_signal_713 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_718 ;
    wire new_AGEMA_signal_719 ;
    wire new_AGEMA_signal_720 ;
    wire new_AGEMA_signal_721 ;
    wire new_AGEMA_signal_722 ;
    wire new_AGEMA_signal_723 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_725 ;
    wire new_AGEMA_signal_726 ;
    wire new_AGEMA_signal_727 ;
    wire new_AGEMA_signal_728 ;
    wire new_AGEMA_signal_729 ;
    wire new_AGEMA_signal_730 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_735 ;
    wire new_AGEMA_signal_736 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_739 ;
    wire new_AGEMA_signal_740 ;
    wire new_AGEMA_signal_741 ;
    wire new_AGEMA_signal_742 ;
    wire new_AGEMA_signal_743 ;
    wire new_AGEMA_signal_744 ;
    wire new_AGEMA_signal_745 ;
    wire new_AGEMA_signal_746 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_749 ;
    wire new_AGEMA_signal_750 ;
    wire new_AGEMA_signal_751 ;
    wire new_AGEMA_signal_752 ;
    wire new_AGEMA_signal_753 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_759 ;
    wire new_AGEMA_signal_760 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_762 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_767 ;
    wire new_AGEMA_signal_768 ;
    wire new_AGEMA_signal_769 ;
    wire new_AGEMA_signal_770 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_782 ;
    wire new_AGEMA_signal_783 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_792 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_799 ;
    wire new_AGEMA_signal_800 ;
    wire new_AGEMA_signal_801 ;
    wire new_AGEMA_signal_802 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_808 ;
    wire new_AGEMA_signal_809 ;
    wire new_AGEMA_signal_810 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_833 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_839 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_842 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U39 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_n25}), .c ({new_AGEMA_signal_283, new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_n12}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U38 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_295, new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_Y_4_}), .c ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_n24}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U37 ( .a ({new_AGEMA_signal_239, new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_Y_2_}), .b ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_n10}), .c ({new_AGEMA_signal_287, new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_n23}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U36 ( .a ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_n9}), .b ({new_AGEMA_signal_215, new_AGEMA_signal_214, new_AGEMA_signal_213, new_AGEMA_signal_212, sbe_n8}), .c ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n22}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U35 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n11}), .c ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n21}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U29 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_n10}), .c ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_Y_6_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U28 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_203, new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, sbe_Y_5_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U27 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_n10}), .c ({new_AGEMA_signal_295, new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_Y_4_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U26 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_n9}), .c ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_n10}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U25 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_215, new_AGEMA_signal_214, new_AGEMA_signal_213, new_AGEMA_signal_212, sbe_n8}), .c ({new_AGEMA_signal_239, new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_Y_2_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U24 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_215, new_AGEMA_signal_214, new_AGEMA_signal_213, new_AGEMA_signal_212, sbe_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U23 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_n7}), .c ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_Y_1_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U22 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_299, new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_B_6_}), .c ({new_AGEMA_signal_319, new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_Y_0_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U8 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_n25}), .c ({new_AGEMA_signal_299, new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_B_6_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U7 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_n9}), .c ({new_AGEMA_signal_271, new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_n25}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U6 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, sbe_n2}), .c ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_n9}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U5 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_n3}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n11}), .c ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_B_3_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U4 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_n7}), .c ({new_AGEMA_signal_275, new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_n3}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U3 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, sbe_n2}), .c ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_n7}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U2 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n11}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, sbe_n2}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m7_U2 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_sel_in_m7_n8}), .b ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_Z[7]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n11}), .a ({new_AGEMA_signal_287, new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_n23}), .c ({new_AGEMA_signal_323, new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_sel_in_m7_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m6_U2 ( .a ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_sel_in_m6_n8}), .b ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_Z[6]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_Y_6_}), .a ({new_AGEMA_signal_299, new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_B_6_}), .c ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_sel_in_m6_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m5_U2 ( .a ({new_AGEMA_signal_331, new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_sel_in_m5_n8}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_Z[5]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_203, new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, sbe_Y_5_}), .a ({new_AGEMA_signal_283, new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_n12}), .c ({new_AGEMA_signal_331, new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_sel_in_m5_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m4_U2 ( .a ({new_AGEMA_signal_335, new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_sel_in_m4_n8}), .b ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_Z[4]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_295, new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_Y_4_}), .a ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n22}), .c ({new_AGEMA_signal_335, new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_sel_in_m4_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m3_U2 ( .a ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_sel_in_m3_n8}), .b ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_Z[3]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n21}), .a ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_B_3_}), .c ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_sel_in_m3_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m2_U2 ( .a ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_sel_in_m2_n8}), .b ({new_AGEMA_signal_307, new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_Z[2]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_239, new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_Y_2_}), .a ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, sbe_n2}), .c ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_sel_in_m2_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m1_U2 ( .a ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_sel_in_m1_n8}), .b ({new_AGEMA_signal_343, new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_Z[1]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_Y_1_}), .a ({new_AGEMA_signal_271, new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_n25}), .c ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_sel_in_m1_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m0_U2 ( .a ({new_AGEMA_signal_367, new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_sel_in_m0_n8}), .b ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_Z[0]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_in_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_319, new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_Y_0_}), .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_n24}), .c ({new_AGEMA_signal_367, new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_sel_in_m0_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U10 ( .a ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_Z[0]}), .b ({new_AGEMA_signal_343, new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_Z[1]}), .c ({new_AGEMA_signal_427, new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_bl}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U9 ( .a ({new_AGEMA_signal_307, new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_Z[2]}), .b ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_Z[3]}), .c ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_bh}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U8 ( .a ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_sb_0_}), .b ({new_AGEMA_signal_391, new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_sb_1_}), .c ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_inv_bb}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U7 ( .a ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_Z[0]}), .b ({new_AGEMA_signal_307, new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_Z[2]}), .c ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_sb_0_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U6 ( .a ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_Z[3]}), .b ({new_AGEMA_signal_343, new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_Z[1]}), .c ({new_AGEMA_signal_391, new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_sb_1_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U5 ( .a ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_Z[4]}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_Z[5]}), .c ({new_AGEMA_signal_395, new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_al}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U4 ( .a ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_Z[6]}), .b ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_Z[7]}), .c ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_ah}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U3 ( .a ({new_AGEMA_signal_403, new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_sa_1_}), .c ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_aa}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U2 ( .a ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_Z[4]}), .b ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_Z[6]}), .c ({new_AGEMA_signal_403, new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_sa_0_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U1 ( .a ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_Z[7]}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_Z[5]}), .c ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_sa_1_}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_236 ( .C ( clk ), .D ( sbe_Z[3] ), .Q ( new_AGEMA_signal_1388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C ( clk ), .D ( new_AGEMA_signal_360 ), .Q ( new_AGEMA_signal_1394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C ( clk ), .D ( new_AGEMA_signal_361 ), .Q ( new_AGEMA_signal_1400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C ( clk ), .D ( new_AGEMA_signal_362 ), .Q ( new_AGEMA_signal_1406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C ( clk ), .D ( new_AGEMA_signal_363 ), .Q ( new_AGEMA_signal_1412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C ( clk ), .D ( sbe_Z[2] ), .Q ( new_AGEMA_signal_1418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C ( clk ), .D ( new_AGEMA_signal_304 ), .Q ( new_AGEMA_signal_1424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C ( clk ), .D ( new_AGEMA_signal_305 ), .Q ( new_AGEMA_signal_1430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C ( clk ), .D ( new_AGEMA_signal_306 ), .Q ( new_AGEMA_signal_1436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C ( clk ), .D ( new_AGEMA_signal_307 ), .Q ( new_AGEMA_signal_1442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C ( clk ), .D ( sbe_inv_bh ), .Q ( new_AGEMA_signal_1448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C ( clk ), .D ( new_AGEMA_signal_384 ), .Q ( new_AGEMA_signal_1454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C ( clk ), .D ( new_AGEMA_signal_385 ), .Q ( new_AGEMA_signal_1460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C ( clk ), .D ( new_AGEMA_signal_386 ), .Q ( new_AGEMA_signal_1466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C ( clk ), .D ( new_AGEMA_signal_387 ), .Q ( new_AGEMA_signal_1472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C ( clk ), .D ( sbe_Z[1] ), .Q ( new_AGEMA_signal_1478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C ( clk ), .D ( new_AGEMA_signal_340 ), .Q ( new_AGEMA_signal_1484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C ( clk ), .D ( new_AGEMA_signal_341 ), .Q ( new_AGEMA_signal_1490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C ( clk ), .D ( new_AGEMA_signal_342 ), .Q ( new_AGEMA_signal_1496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C ( clk ), .D ( new_AGEMA_signal_343 ), .Q ( new_AGEMA_signal_1502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C ( clk ), .D ( sbe_Z[0] ), .Q ( new_AGEMA_signal_1508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C ( clk ), .D ( new_AGEMA_signal_368 ), .Q ( new_AGEMA_signal_1514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C ( clk ), .D ( new_AGEMA_signal_369 ), .Q ( new_AGEMA_signal_1520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C ( clk ), .D ( new_AGEMA_signal_370 ), .Q ( new_AGEMA_signal_1526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C ( clk ), .D ( new_AGEMA_signal_371 ), .Q ( new_AGEMA_signal_1532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C ( clk ), .D ( sbe_inv_bl ), .Q ( new_AGEMA_signal_1538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C ( clk ), .D ( new_AGEMA_signal_424 ), .Q ( new_AGEMA_signal_1544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C ( clk ), .D ( new_AGEMA_signal_425 ), .Q ( new_AGEMA_signal_1550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_404 ( .C ( clk ), .D ( new_AGEMA_signal_426 ), .Q ( new_AGEMA_signal_1556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_410 ( .C ( clk ), .D ( new_AGEMA_signal_427 ), .Q ( new_AGEMA_signal_1562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_416 ( .C ( clk ), .D ( sbe_inv_bb ), .Q ( new_AGEMA_signal_1568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_422 ( .C ( clk ), .D ( new_AGEMA_signal_456 ), .Q ( new_AGEMA_signal_1574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_428 ( .C ( clk ), .D ( new_AGEMA_signal_457 ), .Q ( new_AGEMA_signal_1580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_434 ( .C ( clk ), .D ( new_AGEMA_signal_458 ), .Q ( new_AGEMA_signal_1586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_440 ( .C ( clk ), .D ( new_AGEMA_signal_459 ), .Q ( new_AGEMA_signal_1592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_446 ( .C ( clk ), .D ( sbe_inv_sb_1_ ), .Q ( new_AGEMA_signal_1598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_452 ( .C ( clk ), .D ( new_AGEMA_signal_388 ), .Q ( new_AGEMA_signal_1604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_458 ( .C ( clk ), .D ( new_AGEMA_signal_389 ), .Q ( new_AGEMA_signal_1610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_464 ( .C ( clk ), .D ( new_AGEMA_signal_390 ), .Q ( new_AGEMA_signal_1616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_470 ( .C ( clk ), .D ( new_AGEMA_signal_391 ), .Q ( new_AGEMA_signal_1622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_476 ( .C ( clk ), .D ( sbe_inv_sb_0_ ), .Q ( new_AGEMA_signal_1628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_482 ( .C ( clk ), .D ( new_AGEMA_signal_428 ), .Q ( new_AGEMA_signal_1634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_488 ( .C ( clk ), .D ( new_AGEMA_signal_429 ), .Q ( new_AGEMA_signal_1640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_494 ( .C ( clk ), .D ( new_AGEMA_signal_430 ), .Q ( new_AGEMA_signal_1646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_500 ( .C ( clk ), .D ( new_AGEMA_signal_431 ), .Q ( new_AGEMA_signal_1652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_506 ( .C ( clk ), .D ( sbe_Z[7] ), .Q ( new_AGEMA_signal_1658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_512 ( .C ( clk ), .D ( new_AGEMA_signal_344 ), .Q ( new_AGEMA_signal_1664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_518 ( .C ( clk ), .D ( new_AGEMA_signal_345 ), .Q ( new_AGEMA_signal_1670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_524 ( .C ( clk ), .D ( new_AGEMA_signal_346 ), .Q ( new_AGEMA_signal_1676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_530 ( .C ( clk ), .D ( new_AGEMA_signal_347 ), .Q ( new_AGEMA_signal_1682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_536 ( .C ( clk ), .D ( sbe_Z[6] ), .Q ( new_AGEMA_signal_1688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_542 ( .C ( clk ), .D ( new_AGEMA_signal_348 ), .Q ( new_AGEMA_signal_1694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_548 ( .C ( clk ), .D ( new_AGEMA_signal_349 ), .Q ( new_AGEMA_signal_1700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_554 ( .C ( clk ), .D ( new_AGEMA_signal_350 ), .Q ( new_AGEMA_signal_1706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_560 ( .C ( clk ), .D ( new_AGEMA_signal_351 ), .Q ( new_AGEMA_signal_1712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_566 ( .C ( clk ), .D ( sbe_inv_ah ), .Q ( new_AGEMA_signal_1718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_572 ( .C ( clk ), .D ( new_AGEMA_signal_396 ), .Q ( new_AGEMA_signal_1724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_578 ( .C ( clk ), .D ( new_AGEMA_signal_397 ), .Q ( new_AGEMA_signal_1730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_584 ( .C ( clk ), .D ( new_AGEMA_signal_398 ), .Q ( new_AGEMA_signal_1736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_590 ( .C ( clk ), .D ( new_AGEMA_signal_399 ), .Q ( new_AGEMA_signal_1742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_596 ( .C ( clk ), .D ( sbe_Z[5] ), .Q ( new_AGEMA_signal_1748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_602 ( .C ( clk ), .D ( new_AGEMA_signal_352 ), .Q ( new_AGEMA_signal_1754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_608 ( .C ( clk ), .D ( new_AGEMA_signal_353 ), .Q ( new_AGEMA_signal_1760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_614 ( .C ( clk ), .D ( new_AGEMA_signal_354 ), .Q ( new_AGEMA_signal_1766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_620 ( .C ( clk ), .D ( new_AGEMA_signal_355 ), .Q ( new_AGEMA_signal_1772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_626 ( .C ( clk ), .D ( sbe_Z[4] ), .Q ( new_AGEMA_signal_1778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_632 ( .C ( clk ), .D ( new_AGEMA_signal_356 ), .Q ( new_AGEMA_signal_1784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_638 ( .C ( clk ), .D ( new_AGEMA_signal_357 ), .Q ( new_AGEMA_signal_1790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_644 ( .C ( clk ), .D ( new_AGEMA_signal_358 ), .Q ( new_AGEMA_signal_1796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_650 ( .C ( clk ), .D ( new_AGEMA_signal_359 ), .Q ( new_AGEMA_signal_1802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_656 ( .C ( clk ), .D ( sbe_inv_al ), .Q ( new_AGEMA_signal_1808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_662 ( .C ( clk ), .D ( new_AGEMA_signal_392 ), .Q ( new_AGEMA_signal_1814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_668 ( .C ( clk ), .D ( new_AGEMA_signal_393 ), .Q ( new_AGEMA_signal_1820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_674 ( .C ( clk ), .D ( new_AGEMA_signal_394 ), .Q ( new_AGEMA_signal_1826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_680 ( .C ( clk ), .D ( new_AGEMA_signal_395 ), .Q ( new_AGEMA_signal_1832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_686 ( .C ( clk ), .D ( sbe_inv_aa ), .Q ( new_AGEMA_signal_1838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_692 ( .C ( clk ), .D ( new_AGEMA_signal_432 ), .Q ( new_AGEMA_signal_1844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_698 ( .C ( clk ), .D ( new_AGEMA_signal_433 ), .Q ( new_AGEMA_signal_1850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_704 ( .C ( clk ), .D ( new_AGEMA_signal_434 ), .Q ( new_AGEMA_signal_1856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_710 ( .C ( clk ), .D ( new_AGEMA_signal_435 ), .Q ( new_AGEMA_signal_1862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_716 ( .C ( clk ), .D ( sbe_inv_sa_1_ ), .Q ( new_AGEMA_signal_1868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_722 ( .C ( clk ), .D ( new_AGEMA_signal_404 ), .Q ( new_AGEMA_signal_1874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_728 ( .C ( clk ), .D ( new_AGEMA_signal_405 ), .Q ( new_AGEMA_signal_1880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_734 ( .C ( clk ), .D ( new_AGEMA_signal_406 ), .Q ( new_AGEMA_signal_1886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_740 ( .C ( clk ), .D ( new_AGEMA_signal_407 ), .Q ( new_AGEMA_signal_1892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_746 ( .C ( clk ), .D ( sbe_inv_sa_0_ ), .Q ( new_AGEMA_signal_1898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_752 ( .C ( clk ), .D ( new_AGEMA_signal_400 ), .Q ( new_AGEMA_signal_1904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_758 ( .C ( clk ), .D ( new_AGEMA_signal_401 ), .Q ( new_AGEMA_signal_1910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_764 ( .C ( clk ), .D ( new_AGEMA_signal_402 ), .Q ( new_AGEMA_signal_1916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_770 ( .C ( clk ), .D ( new_AGEMA_signal_403 ), .Q ( new_AGEMA_signal_1922 ) ) ;

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U34 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_n21}), .b ({new_AGEMA_signal_463, new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_inv_n20}), .c ({new_AGEMA_signal_499, new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_inv_c[3]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U33 ( .a ({new_AGEMA_signal_439, new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_n19}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_n18}), .c ({new_AGEMA_signal_463, new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_inv_n20}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U32 ( .a ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_Z[7]}), .b ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_Z[3]}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_n18}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U31 ( .a ({new_AGEMA_signal_403, new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_439, new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_n19}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U30 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_inv_n17}), .b ({new_AGEMA_signal_415, new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_n16}), .c ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_n21}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U29 ( .a ({new_AGEMA_signal_467, new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_n15}), .b ({new_AGEMA_signal_443, new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_n14}), .c ({new_AGEMA_signal_487, new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_inv_c[2]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U28 ( .a ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_n13}), .b ({new_AGEMA_signal_379, new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_n12}), .c ({new_AGEMA_signal_443, new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_n14}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U27 ( .a ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_Z[6]}), .b ({new_AGEMA_signal_307, new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_Z[2]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_379, new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_n12}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U26 ( .a ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_sa_1_}), .b ({new_AGEMA_signal_391, new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_sb_1_}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_n13}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U25 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_n11}), .b ({new_AGEMA_signal_415, new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_n16}), .c ({new_AGEMA_signal_467, new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_n15}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U24 ( .a ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_ah}), .b ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_bh}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_415, new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_n16}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U23 ( .a ({new_AGEMA_signal_491, new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_inv_n10}), .b ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_inv_n9}), .c ({new_AGEMA_signal_503, new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_inv_c[1]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U22 ( .a ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_n8}), .b ({new_AGEMA_signal_383, new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_n7}), .c ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_inv_n9}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U21 ( .a ({new_AGEMA_signal_343, new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_Z[1]}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_Z[5]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_383, new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_n7}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U20 ( .a ({new_AGEMA_signal_395, new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_al}), .b ({new_AGEMA_signal_427, new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_n8}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U19 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_inv_n17}), .b ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_n11}), .c ({new_AGEMA_signal_491, new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_inv_n10}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U18 ( .a ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_aa}), .b ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_inv_bb}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_475, new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_inv_n17}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U17 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_n11}), .b ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_n6}), .c ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_inv_c[0]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U16 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_n5}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_inv_n4}), .c ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_n6}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U15 ( .a ({new_AGEMA_signal_419, new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_n3}), .b ({new_AGEMA_signal_451, new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_n2}), .c ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_inv_n4}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U14 ( .a ({new_AGEMA_signal_395, new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_al}), .b ({new_AGEMA_signal_427, new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_451, new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_n2}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U13 ( .a ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_Z[4]}), .b ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_Z[0]}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_419, new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_n3}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U12 ( .a ({new_AGEMA_signal_391, new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_sb_1_}), .b ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_sa_1_}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_n5}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U11 ( .a ({new_AGEMA_signal_403, new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_n11}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U2 ( .a ({new_AGEMA_signal_487, new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_inv_c[2]}), .b ({new_AGEMA_signal_499, new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_inv_c[3]}), .c ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_inv_dinv_sa}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U1 ( .a ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_inv_c[0]}), .b ({new_AGEMA_signal_503, new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_inv_c[1]}), .c ({new_AGEMA_signal_523, new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_inv_dinv_sb}) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C ( clk ), .D ( new_AGEMA_signal_1388 ), .Q ( new_AGEMA_signal_1389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C ( clk ), .D ( new_AGEMA_signal_1394 ), .Q ( new_AGEMA_signal_1395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C ( clk ), .D ( new_AGEMA_signal_1400 ), .Q ( new_AGEMA_signal_1401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C ( clk ), .D ( new_AGEMA_signal_1406 ), .Q ( new_AGEMA_signal_1407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C ( clk ), .D ( new_AGEMA_signal_1412 ), .Q ( new_AGEMA_signal_1413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C ( clk ), .D ( new_AGEMA_signal_1418 ), .Q ( new_AGEMA_signal_1419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C ( clk ), .D ( new_AGEMA_signal_1424 ), .Q ( new_AGEMA_signal_1425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C ( clk ), .D ( new_AGEMA_signal_1430 ), .Q ( new_AGEMA_signal_1431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C ( clk ), .D ( new_AGEMA_signal_1436 ), .Q ( new_AGEMA_signal_1437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C ( clk ), .D ( new_AGEMA_signal_1442 ), .Q ( new_AGEMA_signal_1443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C ( clk ), .D ( new_AGEMA_signal_1448 ), .Q ( new_AGEMA_signal_1449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C ( clk ), .D ( new_AGEMA_signal_1454 ), .Q ( new_AGEMA_signal_1455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C ( clk ), .D ( new_AGEMA_signal_1460 ), .Q ( new_AGEMA_signal_1461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C ( clk ), .D ( new_AGEMA_signal_1466 ), .Q ( new_AGEMA_signal_1467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C ( clk ), .D ( new_AGEMA_signal_1472 ), .Q ( new_AGEMA_signal_1473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C ( clk ), .D ( new_AGEMA_signal_1478 ), .Q ( new_AGEMA_signal_1479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C ( clk ), .D ( new_AGEMA_signal_1484 ), .Q ( new_AGEMA_signal_1485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C ( clk ), .D ( new_AGEMA_signal_1490 ), .Q ( new_AGEMA_signal_1491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C ( clk ), .D ( new_AGEMA_signal_1496 ), .Q ( new_AGEMA_signal_1497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C ( clk ), .D ( new_AGEMA_signal_1502 ), .Q ( new_AGEMA_signal_1503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C ( clk ), .D ( new_AGEMA_signal_1508 ), .Q ( new_AGEMA_signal_1509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C ( clk ), .D ( new_AGEMA_signal_1514 ), .Q ( new_AGEMA_signal_1515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C ( clk ), .D ( new_AGEMA_signal_1520 ), .Q ( new_AGEMA_signal_1521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C ( clk ), .D ( new_AGEMA_signal_1526 ), .Q ( new_AGEMA_signal_1527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C ( clk ), .D ( new_AGEMA_signal_1532 ), .Q ( new_AGEMA_signal_1533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C ( clk ), .D ( new_AGEMA_signal_1538 ), .Q ( new_AGEMA_signal_1539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C ( clk ), .D ( new_AGEMA_signal_1544 ), .Q ( new_AGEMA_signal_1545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C ( clk ), .D ( new_AGEMA_signal_1550 ), .Q ( new_AGEMA_signal_1551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_405 ( .C ( clk ), .D ( new_AGEMA_signal_1556 ), .Q ( new_AGEMA_signal_1557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_411 ( .C ( clk ), .D ( new_AGEMA_signal_1562 ), .Q ( new_AGEMA_signal_1563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_417 ( .C ( clk ), .D ( new_AGEMA_signal_1568 ), .Q ( new_AGEMA_signal_1569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_423 ( .C ( clk ), .D ( new_AGEMA_signal_1574 ), .Q ( new_AGEMA_signal_1575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_429 ( .C ( clk ), .D ( new_AGEMA_signal_1580 ), .Q ( new_AGEMA_signal_1581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_435 ( .C ( clk ), .D ( new_AGEMA_signal_1586 ), .Q ( new_AGEMA_signal_1587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_441 ( .C ( clk ), .D ( new_AGEMA_signal_1592 ), .Q ( new_AGEMA_signal_1593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_447 ( .C ( clk ), .D ( new_AGEMA_signal_1598 ), .Q ( new_AGEMA_signal_1599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_453 ( .C ( clk ), .D ( new_AGEMA_signal_1604 ), .Q ( new_AGEMA_signal_1605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_459 ( .C ( clk ), .D ( new_AGEMA_signal_1610 ), .Q ( new_AGEMA_signal_1611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_465 ( .C ( clk ), .D ( new_AGEMA_signal_1616 ), .Q ( new_AGEMA_signal_1617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_471 ( .C ( clk ), .D ( new_AGEMA_signal_1622 ), .Q ( new_AGEMA_signal_1623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_477 ( .C ( clk ), .D ( new_AGEMA_signal_1628 ), .Q ( new_AGEMA_signal_1629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_483 ( .C ( clk ), .D ( new_AGEMA_signal_1634 ), .Q ( new_AGEMA_signal_1635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_489 ( .C ( clk ), .D ( new_AGEMA_signal_1640 ), .Q ( new_AGEMA_signal_1641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_495 ( .C ( clk ), .D ( new_AGEMA_signal_1646 ), .Q ( new_AGEMA_signal_1647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_501 ( .C ( clk ), .D ( new_AGEMA_signal_1652 ), .Q ( new_AGEMA_signal_1653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_507 ( .C ( clk ), .D ( new_AGEMA_signal_1658 ), .Q ( new_AGEMA_signal_1659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_513 ( .C ( clk ), .D ( new_AGEMA_signal_1664 ), .Q ( new_AGEMA_signal_1665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_519 ( .C ( clk ), .D ( new_AGEMA_signal_1670 ), .Q ( new_AGEMA_signal_1671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_525 ( .C ( clk ), .D ( new_AGEMA_signal_1676 ), .Q ( new_AGEMA_signal_1677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_531 ( .C ( clk ), .D ( new_AGEMA_signal_1682 ), .Q ( new_AGEMA_signal_1683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_537 ( .C ( clk ), .D ( new_AGEMA_signal_1688 ), .Q ( new_AGEMA_signal_1689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_543 ( .C ( clk ), .D ( new_AGEMA_signal_1694 ), .Q ( new_AGEMA_signal_1695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_549 ( .C ( clk ), .D ( new_AGEMA_signal_1700 ), .Q ( new_AGEMA_signal_1701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_555 ( .C ( clk ), .D ( new_AGEMA_signal_1706 ), .Q ( new_AGEMA_signal_1707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_561 ( .C ( clk ), .D ( new_AGEMA_signal_1712 ), .Q ( new_AGEMA_signal_1713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_567 ( .C ( clk ), .D ( new_AGEMA_signal_1718 ), .Q ( new_AGEMA_signal_1719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_573 ( .C ( clk ), .D ( new_AGEMA_signal_1724 ), .Q ( new_AGEMA_signal_1725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_579 ( .C ( clk ), .D ( new_AGEMA_signal_1730 ), .Q ( new_AGEMA_signal_1731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_585 ( .C ( clk ), .D ( new_AGEMA_signal_1736 ), .Q ( new_AGEMA_signal_1737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_591 ( .C ( clk ), .D ( new_AGEMA_signal_1742 ), .Q ( new_AGEMA_signal_1743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_597 ( .C ( clk ), .D ( new_AGEMA_signal_1748 ), .Q ( new_AGEMA_signal_1749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_603 ( .C ( clk ), .D ( new_AGEMA_signal_1754 ), .Q ( new_AGEMA_signal_1755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_609 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_1761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_615 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_1767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_621 ( .C ( clk ), .D ( new_AGEMA_signal_1772 ), .Q ( new_AGEMA_signal_1773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_627 ( .C ( clk ), .D ( new_AGEMA_signal_1778 ), .Q ( new_AGEMA_signal_1779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_633 ( .C ( clk ), .D ( new_AGEMA_signal_1784 ), .Q ( new_AGEMA_signal_1785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_639 ( .C ( clk ), .D ( new_AGEMA_signal_1790 ), .Q ( new_AGEMA_signal_1791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_645 ( .C ( clk ), .D ( new_AGEMA_signal_1796 ), .Q ( new_AGEMA_signal_1797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_651 ( .C ( clk ), .D ( new_AGEMA_signal_1802 ), .Q ( new_AGEMA_signal_1803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_657 ( .C ( clk ), .D ( new_AGEMA_signal_1808 ), .Q ( new_AGEMA_signal_1809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_663 ( .C ( clk ), .D ( new_AGEMA_signal_1814 ), .Q ( new_AGEMA_signal_1815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_669 ( .C ( clk ), .D ( new_AGEMA_signal_1820 ), .Q ( new_AGEMA_signal_1821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_675 ( .C ( clk ), .D ( new_AGEMA_signal_1826 ), .Q ( new_AGEMA_signal_1827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_681 ( .C ( clk ), .D ( new_AGEMA_signal_1832 ), .Q ( new_AGEMA_signal_1833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_687 ( .C ( clk ), .D ( new_AGEMA_signal_1838 ), .Q ( new_AGEMA_signal_1839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_693 ( .C ( clk ), .D ( new_AGEMA_signal_1844 ), .Q ( new_AGEMA_signal_1845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_699 ( .C ( clk ), .D ( new_AGEMA_signal_1850 ), .Q ( new_AGEMA_signal_1851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_705 ( .C ( clk ), .D ( new_AGEMA_signal_1856 ), .Q ( new_AGEMA_signal_1857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_711 ( .C ( clk ), .D ( new_AGEMA_signal_1862 ), .Q ( new_AGEMA_signal_1863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_717 ( .C ( clk ), .D ( new_AGEMA_signal_1868 ), .Q ( new_AGEMA_signal_1869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_723 ( .C ( clk ), .D ( new_AGEMA_signal_1874 ), .Q ( new_AGEMA_signal_1875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_729 ( .C ( clk ), .D ( new_AGEMA_signal_1880 ), .Q ( new_AGEMA_signal_1881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_735 ( .C ( clk ), .D ( new_AGEMA_signal_1886 ), .Q ( new_AGEMA_signal_1887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_741 ( .C ( clk ), .D ( new_AGEMA_signal_1892 ), .Q ( new_AGEMA_signal_1893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_747 ( .C ( clk ), .D ( new_AGEMA_signal_1898 ), .Q ( new_AGEMA_signal_1899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_753 ( .C ( clk ), .D ( new_AGEMA_signal_1904 ), .Q ( new_AGEMA_signal_1905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_759 ( .C ( clk ), .D ( new_AGEMA_signal_1910 ), .Q ( new_AGEMA_signal_1911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_765 ( .C ( clk ), .D ( new_AGEMA_signal_1916 ), .Q ( new_AGEMA_signal_1917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_771 ( .C ( clk ), .D ( new_AGEMA_signal_1922 ), .Q ( new_AGEMA_signal_1923 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( sbe_inv_c[1] ), .Q ( new_AGEMA_signal_1328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( new_AGEMA_signal_500 ), .Q ( new_AGEMA_signal_1330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( new_AGEMA_signal_501 ), .Q ( new_AGEMA_signal_1332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( new_AGEMA_signal_502 ), .Q ( new_AGEMA_signal_1334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( new_AGEMA_signal_503 ), .Q ( new_AGEMA_signal_1336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( sbe_inv_c[0] ), .Q ( new_AGEMA_signal_1338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( new_AGEMA_signal_504 ), .Q ( new_AGEMA_signal_1340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_505 ), .Q ( new_AGEMA_signal_1342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C ( clk ), .D ( new_AGEMA_signal_506 ), .Q ( new_AGEMA_signal_1344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C ( clk ), .D ( new_AGEMA_signal_507 ), .Q ( new_AGEMA_signal_1346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C ( clk ), .D ( sbe_inv_dinv_sb ), .Q ( new_AGEMA_signal_1348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C ( clk ), .D ( new_AGEMA_signal_520 ), .Q ( new_AGEMA_signal_1350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C ( clk ), .D ( new_AGEMA_signal_521 ), .Q ( new_AGEMA_signal_1352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C ( clk ), .D ( new_AGEMA_signal_522 ), .Q ( new_AGEMA_signal_1354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C ( clk ), .D ( new_AGEMA_signal_523 ), .Q ( new_AGEMA_signal_1356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C ( clk ), .D ( sbe_inv_c[3] ), .Q ( new_AGEMA_signal_1358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C ( clk ), .D ( new_AGEMA_signal_496 ), .Q ( new_AGEMA_signal_1360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C ( clk ), .D ( new_AGEMA_signal_497 ), .Q ( new_AGEMA_signal_1362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C ( clk ), .D ( new_AGEMA_signal_498 ), .Q ( new_AGEMA_signal_1364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C ( clk ), .D ( new_AGEMA_signal_499 ), .Q ( new_AGEMA_signal_1366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C ( clk ), .D ( sbe_inv_c[2] ), .Q ( new_AGEMA_signal_1368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C ( clk ), .D ( new_AGEMA_signal_484 ), .Q ( new_AGEMA_signal_1370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C ( clk ), .D ( new_AGEMA_signal_485 ), .Q ( new_AGEMA_signal_1372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C ( clk ), .D ( new_AGEMA_signal_486 ), .Q ( new_AGEMA_signal_1374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C ( clk ), .D ( new_AGEMA_signal_487 ), .Q ( new_AGEMA_signal_1376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C ( clk ), .D ( sbe_inv_dinv_sa ), .Q ( new_AGEMA_signal_1378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C ( clk ), .D ( new_AGEMA_signal_516 ), .Q ( new_AGEMA_signal_1380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C ( clk ), .D ( new_AGEMA_signal_517 ), .Q ( new_AGEMA_signal_1382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C ( clk ), .D ( new_AGEMA_signal_518 ), .Q ( new_AGEMA_signal_1384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C ( clk ), .D ( new_AGEMA_signal_519 ), .Q ( new_AGEMA_signal_1386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C ( clk ), .D ( new_AGEMA_signal_1389 ), .Q ( new_AGEMA_signal_1390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C ( clk ), .D ( new_AGEMA_signal_1395 ), .Q ( new_AGEMA_signal_1396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C ( clk ), .D ( new_AGEMA_signal_1401 ), .Q ( new_AGEMA_signal_1402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C ( clk ), .D ( new_AGEMA_signal_1407 ), .Q ( new_AGEMA_signal_1408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C ( clk ), .D ( new_AGEMA_signal_1413 ), .Q ( new_AGEMA_signal_1414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C ( clk ), .D ( new_AGEMA_signal_1419 ), .Q ( new_AGEMA_signal_1420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C ( clk ), .D ( new_AGEMA_signal_1425 ), .Q ( new_AGEMA_signal_1426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C ( clk ), .D ( new_AGEMA_signal_1431 ), .Q ( new_AGEMA_signal_1432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C ( clk ), .D ( new_AGEMA_signal_1437 ), .Q ( new_AGEMA_signal_1438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C ( clk ), .D ( new_AGEMA_signal_1443 ), .Q ( new_AGEMA_signal_1444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C ( clk ), .D ( new_AGEMA_signal_1449 ), .Q ( new_AGEMA_signal_1450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C ( clk ), .D ( new_AGEMA_signal_1455 ), .Q ( new_AGEMA_signal_1456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C ( clk ), .D ( new_AGEMA_signal_1461 ), .Q ( new_AGEMA_signal_1462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C ( clk ), .D ( new_AGEMA_signal_1467 ), .Q ( new_AGEMA_signal_1468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C ( clk ), .D ( new_AGEMA_signal_1473 ), .Q ( new_AGEMA_signal_1474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C ( clk ), .D ( new_AGEMA_signal_1479 ), .Q ( new_AGEMA_signal_1480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C ( clk ), .D ( new_AGEMA_signal_1485 ), .Q ( new_AGEMA_signal_1486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C ( clk ), .D ( new_AGEMA_signal_1491 ), .Q ( new_AGEMA_signal_1492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C ( clk ), .D ( new_AGEMA_signal_1497 ), .Q ( new_AGEMA_signal_1498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C ( clk ), .D ( new_AGEMA_signal_1503 ), .Q ( new_AGEMA_signal_1504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C ( clk ), .D ( new_AGEMA_signal_1509 ), .Q ( new_AGEMA_signal_1510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C ( clk ), .D ( new_AGEMA_signal_1515 ), .Q ( new_AGEMA_signal_1516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C ( clk ), .D ( new_AGEMA_signal_1521 ), .Q ( new_AGEMA_signal_1522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C ( clk ), .D ( new_AGEMA_signal_1527 ), .Q ( new_AGEMA_signal_1528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C ( clk ), .D ( new_AGEMA_signal_1533 ), .Q ( new_AGEMA_signal_1534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C ( clk ), .D ( new_AGEMA_signal_1539 ), .Q ( new_AGEMA_signal_1540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C ( clk ), .D ( new_AGEMA_signal_1545 ), .Q ( new_AGEMA_signal_1546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_400 ( .C ( clk ), .D ( new_AGEMA_signal_1551 ), .Q ( new_AGEMA_signal_1552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_406 ( .C ( clk ), .D ( new_AGEMA_signal_1557 ), .Q ( new_AGEMA_signal_1558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_412 ( .C ( clk ), .D ( new_AGEMA_signal_1563 ), .Q ( new_AGEMA_signal_1564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_418 ( .C ( clk ), .D ( new_AGEMA_signal_1569 ), .Q ( new_AGEMA_signal_1570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_424 ( .C ( clk ), .D ( new_AGEMA_signal_1575 ), .Q ( new_AGEMA_signal_1576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_430 ( .C ( clk ), .D ( new_AGEMA_signal_1581 ), .Q ( new_AGEMA_signal_1582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_436 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_1588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_442 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_1594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_448 ( .C ( clk ), .D ( new_AGEMA_signal_1599 ), .Q ( new_AGEMA_signal_1600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_454 ( .C ( clk ), .D ( new_AGEMA_signal_1605 ), .Q ( new_AGEMA_signal_1606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_460 ( .C ( clk ), .D ( new_AGEMA_signal_1611 ), .Q ( new_AGEMA_signal_1612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_466 ( .C ( clk ), .D ( new_AGEMA_signal_1617 ), .Q ( new_AGEMA_signal_1618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_472 ( .C ( clk ), .D ( new_AGEMA_signal_1623 ), .Q ( new_AGEMA_signal_1624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_478 ( .C ( clk ), .D ( new_AGEMA_signal_1629 ), .Q ( new_AGEMA_signal_1630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_484 ( .C ( clk ), .D ( new_AGEMA_signal_1635 ), .Q ( new_AGEMA_signal_1636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_490 ( .C ( clk ), .D ( new_AGEMA_signal_1641 ), .Q ( new_AGEMA_signal_1642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_496 ( .C ( clk ), .D ( new_AGEMA_signal_1647 ), .Q ( new_AGEMA_signal_1648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_502 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_1654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_508 ( .C ( clk ), .D ( new_AGEMA_signal_1659 ), .Q ( new_AGEMA_signal_1660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_514 ( .C ( clk ), .D ( new_AGEMA_signal_1665 ), .Q ( new_AGEMA_signal_1666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_520 ( .C ( clk ), .D ( new_AGEMA_signal_1671 ), .Q ( new_AGEMA_signal_1672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_526 ( .C ( clk ), .D ( new_AGEMA_signal_1677 ), .Q ( new_AGEMA_signal_1678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_532 ( .C ( clk ), .D ( new_AGEMA_signal_1683 ), .Q ( new_AGEMA_signal_1684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_538 ( .C ( clk ), .D ( new_AGEMA_signal_1689 ), .Q ( new_AGEMA_signal_1690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_544 ( .C ( clk ), .D ( new_AGEMA_signal_1695 ), .Q ( new_AGEMA_signal_1696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_550 ( .C ( clk ), .D ( new_AGEMA_signal_1701 ), .Q ( new_AGEMA_signal_1702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_556 ( .C ( clk ), .D ( new_AGEMA_signal_1707 ), .Q ( new_AGEMA_signal_1708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_562 ( .C ( clk ), .D ( new_AGEMA_signal_1713 ), .Q ( new_AGEMA_signal_1714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_568 ( .C ( clk ), .D ( new_AGEMA_signal_1719 ), .Q ( new_AGEMA_signal_1720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_574 ( .C ( clk ), .D ( new_AGEMA_signal_1725 ), .Q ( new_AGEMA_signal_1726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_580 ( .C ( clk ), .D ( new_AGEMA_signal_1731 ), .Q ( new_AGEMA_signal_1732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_586 ( .C ( clk ), .D ( new_AGEMA_signal_1737 ), .Q ( new_AGEMA_signal_1738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_592 ( .C ( clk ), .D ( new_AGEMA_signal_1743 ), .Q ( new_AGEMA_signal_1744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_598 ( .C ( clk ), .D ( new_AGEMA_signal_1749 ), .Q ( new_AGEMA_signal_1750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_604 ( .C ( clk ), .D ( new_AGEMA_signal_1755 ), .Q ( new_AGEMA_signal_1756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_610 ( .C ( clk ), .D ( new_AGEMA_signal_1761 ), .Q ( new_AGEMA_signal_1762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_616 ( .C ( clk ), .D ( new_AGEMA_signal_1767 ), .Q ( new_AGEMA_signal_1768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_622 ( .C ( clk ), .D ( new_AGEMA_signal_1773 ), .Q ( new_AGEMA_signal_1774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_628 ( .C ( clk ), .D ( new_AGEMA_signal_1779 ), .Q ( new_AGEMA_signal_1780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_634 ( .C ( clk ), .D ( new_AGEMA_signal_1785 ), .Q ( new_AGEMA_signal_1786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_640 ( .C ( clk ), .D ( new_AGEMA_signal_1791 ), .Q ( new_AGEMA_signal_1792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_646 ( .C ( clk ), .D ( new_AGEMA_signal_1797 ), .Q ( new_AGEMA_signal_1798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_652 ( .C ( clk ), .D ( new_AGEMA_signal_1803 ), .Q ( new_AGEMA_signal_1804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_658 ( .C ( clk ), .D ( new_AGEMA_signal_1809 ), .Q ( new_AGEMA_signal_1810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_664 ( .C ( clk ), .D ( new_AGEMA_signal_1815 ), .Q ( new_AGEMA_signal_1816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_670 ( .C ( clk ), .D ( new_AGEMA_signal_1821 ), .Q ( new_AGEMA_signal_1822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_676 ( .C ( clk ), .D ( new_AGEMA_signal_1827 ), .Q ( new_AGEMA_signal_1828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_682 ( .C ( clk ), .D ( new_AGEMA_signal_1833 ), .Q ( new_AGEMA_signal_1834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_688 ( .C ( clk ), .D ( new_AGEMA_signal_1839 ), .Q ( new_AGEMA_signal_1840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_694 ( .C ( clk ), .D ( new_AGEMA_signal_1845 ), .Q ( new_AGEMA_signal_1846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_700 ( .C ( clk ), .D ( new_AGEMA_signal_1851 ), .Q ( new_AGEMA_signal_1852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_706 ( .C ( clk ), .D ( new_AGEMA_signal_1857 ), .Q ( new_AGEMA_signal_1858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_712 ( .C ( clk ), .D ( new_AGEMA_signal_1863 ), .Q ( new_AGEMA_signal_1864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_718 ( .C ( clk ), .D ( new_AGEMA_signal_1869 ), .Q ( new_AGEMA_signal_1870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_724 ( .C ( clk ), .D ( new_AGEMA_signal_1875 ), .Q ( new_AGEMA_signal_1876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_730 ( .C ( clk ), .D ( new_AGEMA_signal_1881 ), .Q ( new_AGEMA_signal_1882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_736 ( .C ( clk ), .D ( new_AGEMA_signal_1887 ), .Q ( new_AGEMA_signal_1888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_742 ( .C ( clk ), .D ( new_AGEMA_signal_1893 ), .Q ( new_AGEMA_signal_1894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_748 ( .C ( clk ), .D ( new_AGEMA_signal_1899 ), .Q ( new_AGEMA_signal_1900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_754 ( .C ( clk ), .D ( new_AGEMA_signal_1905 ), .Q ( new_AGEMA_signal_1906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_760 ( .C ( clk ), .D ( new_AGEMA_signal_1911 ), .Q ( new_AGEMA_signal_1912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_766 ( .C ( clk ), .D ( new_AGEMA_signal_1917 ), .Q ( new_AGEMA_signal_1918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_772 ( .C ( clk ), .D ( new_AGEMA_signal_1923 ), .Q ( new_AGEMA_signal_1924 ) ) ;

    /* cells in depth 4 */
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U9 ( .a ({new_AGEMA_signal_535, new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, sbe_inv_dinv_d_1_}), .c ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_dinv_sd}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U8 ( .a ({new_AGEMA_signal_511, new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_inv_dinv_n4}), .b ({new_AGEMA_signal_527, new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, sbe_inv_dinv_n3}), .c ({new_AGEMA_signal_535, new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_inv_dinv_d_0_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U7 ( .a ({new_AGEMA_signal_523, new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_527, new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, sbe_inv_dinv_n3}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U6 ( .a ({new_AGEMA_signal_503, new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_inv_c[1]}), .b ({new_AGEMA_signal_499, new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_inv_c[3]}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({new_AGEMA_signal_511, new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_inv_dinv_n4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U5 ( .a ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_inv_dinv_n2}), .b ({new_AGEMA_signal_515, new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, sbe_inv_dinv_n1}), .c ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, sbe_inv_dinv_d_1_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U4 ( .a ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_inv_c[0]}), .b ({new_AGEMA_signal_487, new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_inv_c[2]}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_515, new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, sbe_inv_dinv_n1}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_U3 ( .a ({new_AGEMA_signal_523, new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_inv_dinv_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_1328 ), .Q ( new_AGEMA_signal_1329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_1330 ), .Q ( new_AGEMA_signal_1331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_1332 ), .Q ( new_AGEMA_signal_1333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_1334 ), .Q ( new_AGEMA_signal_1335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_1336 ), .Q ( new_AGEMA_signal_1337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_1338 ), .Q ( new_AGEMA_signal_1339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_1340 ), .Q ( new_AGEMA_signal_1341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C ( clk ), .D ( new_AGEMA_signal_1342 ), .Q ( new_AGEMA_signal_1343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C ( clk ), .D ( new_AGEMA_signal_1344 ), .Q ( new_AGEMA_signal_1345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C ( clk ), .D ( new_AGEMA_signal_1346 ), .Q ( new_AGEMA_signal_1347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C ( clk ), .D ( new_AGEMA_signal_1348 ), .Q ( new_AGEMA_signal_1349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C ( clk ), .D ( new_AGEMA_signal_1350 ), .Q ( new_AGEMA_signal_1351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C ( clk ), .D ( new_AGEMA_signal_1352 ), .Q ( new_AGEMA_signal_1353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_1355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C ( clk ), .D ( new_AGEMA_signal_1356 ), .Q ( new_AGEMA_signal_1357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C ( clk ), .D ( new_AGEMA_signal_1358 ), .Q ( new_AGEMA_signal_1359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C ( clk ), .D ( new_AGEMA_signal_1360 ), .Q ( new_AGEMA_signal_1361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C ( clk ), .D ( new_AGEMA_signal_1362 ), .Q ( new_AGEMA_signal_1363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C ( clk ), .D ( new_AGEMA_signal_1364 ), .Q ( new_AGEMA_signal_1365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C ( clk ), .D ( new_AGEMA_signal_1366 ), .Q ( new_AGEMA_signal_1367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_1369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C ( clk ), .D ( new_AGEMA_signal_1370 ), .Q ( new_AGEMA_signal_1371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_1373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C ( clk ), .D ( new_AGEMA_signal_1374 ), .Q ( new_AGEMA_signal_1375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C ( clk ), .D ( new_AGEMA_signal_1376 ), .Q ( new_AGEMA_signal_1377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C ( clk ), .D ( new_AGEMA_signal_1378 ), .Q ( new_AGEMA_signal_1379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C ( clk ), .D ( new_AGEMA_signal_1380 ), .Q ( new_AGEMA_signal_1381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C ( clk ), .D ( new_AGEMA_signal_1382 ), .Q ( new_AGEMA_signal_1383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C ( clk ), .D ( new_AGEMA_signal_1384 ), .Q ( new_AGEMA_signal_1385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C ( clk ), .D ( new_AGEMA_signal_1386 ), .Q ( new_AGEMA_signal_1387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_1391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C ( clk ), .D ( new_AGEMA_signal_1396 ), .Q ( new_AGEMA_signal_1397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C ( clk ), .D ( new_AGEMA_signal_1402 ), .Q ( new_AGEMA_signal_1403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C ( clk ), .D ( new_AGEMA_signal_1408 ), .Q ( new_AGEMA_signal_1409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C ( clk ), .D ( new_AGEMA_signal_1414 ), .Q ( new_AGEMA_signal_1415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C ( clk ), .D ( new_AGEMA_signal_1420 ), .Q ( new_AGEMA_signal_1421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C ( clk ), .D ( new_AGEMA_signal_1426 ), .Q ( new_AGEMA_signal_1427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C ( clk ), .D ( new_AGEMA_signal_1432 ), .Q ( new_AGEMA_signal_1433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_1439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C ( clk ), .D ( new_AGEMA_signal_1444 ), .Q ( new_AGEMA_signal_1445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C ( clk ), .D ( new_AGEMA_signal_1450 ), .Q ( new_AGEMA_signal_1451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_1457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C ( clk ), .D ( new_AGEMA_signal_1462 ), .Q ( new_AGEMA_signal_1463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C ( clk ), .D ( new_AGEMA_signal_1468 ), .Q ( new_AGEMA_signal_1469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C ( clk ), .D ( new_AGEMA_signal_1474 ), .Q ( new_AGEMA_signal_1475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C ( clk ), .D ( new_AGEMA_signal_1480 ), .Q ( new_AGEMA_signal_1481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C ( clk ), .D ( new_AGEMA_signal_1486 ), .Q ( new_AGEMA_signal_1487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C ( clk ), .D ( new_AGEMA_signal_1492 ), .Q ( new_AGEMA_signal_1493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C ( clk ), .D ( new_AGEMA_signal_1498 ), .Q ( new_AGEMA_signal_1499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C ( clk ), .D ( new_AGEMA_signal_1504 ), .Q ( new_AGEMA_signal_1505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C ( clk ), .D ( new_AGEMA_signal_1510 ), .Q ( new_AGEMA_signal_1511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_1517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C ( clk ), .D ( new_AGEMA_signal_1522 ), .Q ( new_AGEMA_signal_1523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C ( clk ), .D ( new_AGEMA_signal_1528 ), .Q ( new_AGEMA_signal_1529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C ( clk ), .D ( new_AGEMA_signal_1534 ), .Q ( new_AGEMA_signal_1535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C ( clk ), .D ( new_AGEMA_signal_1540 ), .Q ( new_AGEMA_signal_1541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C ( clk ), .D ( new_AGEMA_signal_1546 ), .Q ( new_AGEMA_signal_1547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_401 ( .C ( clk ), .D ( new_AGEMA_signal_1552 ), .Q ( new_AGEMA_signal_1553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_407 ( .C ( clk ), .D ( new_AGEMA_signal_1558 ), .Q ( new_AGEMA_signal_1559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_413 ( .C ( clk ), .D ( new_AGEMA_signal_1564 ), .Q ( new_AGEMA_signal_1565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_419 ( .C ( clk ), .D ( new_AGEMA_signal_1570 ), .Q ( new_AGEMA_signal_1571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_425 ( .C ( clk ), .D ( new_AGEMA_signal_1576 ), .Q ( new_AGEMA_signal_1577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_431 ( .C ( clk ), .D ( new_AGEMA_signal_1582 ), .Q ( new_AGEMA_signal_1583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_437 ( .C ( clk ), .D ( new_AGEMA_signal_1588 ), .Q ( new_AGEMA_signal_1589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_443 ( .C ( clk ), .D ( new_AGEMA_signal_1594 ), .Q ( new_AGEMA_signal_1595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_449 ( .C ( clk ), .D ( new_AGEMA_signal_1600 ), .Q ( new_AGEMA_signal_1601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_455 ( .C ( clk ), .D ( new_AGEMA_signal_1606 ), .Q ( new_AGEMA_signal_1607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_461 ( .C ( clk ), .D ( new_AGEMA_signal_1612 ), .Q ( new_AGEMA_signal_1613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_467 ( .C ( clk ), .D ( new_AGEMA_signal_1618 ), .Q ( new_AGEMA_signal_1619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_473 ( .C ( clk ), .D ( new_AGEMA_signal_1624 ), .Q ( new_AGEMA_signal_1625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_479 ( .C ( clk ), .D ( new_AGEMA_signal_1630 ), .Q ( new_AGEMA_signal_1631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_485 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_1637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_491 ( .C ( clk ), .D ( new_AGEMA_signal_1642 ), .Q ( new_AGEMA_signal_1643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_497 ( .C ( clk ), .D ( new_AGEMA_signal_1648 ), .Q ( new_AGEMA_signal_1649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_503 ( .C ( clk ), .D ( new_AGEMA_signal_1654 ), .Q ( new_AGEMA_signal_1655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_509 ( .C ( clk ), .D ( new_AGEMA_signal_1660 ), .Q ( new_AGEMA_signal_1661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_515 ( .C ( clk ), .D ( new_AGEMA_signal_1666 ), .Q ( new_AGEMA_signal_1667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_521 ( .C ( clk ), .D ( new_AGEMA_signal_1672 ), .Q ( new_AGEMA_signal_1673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_527 ( .C ( clk ), .D ( new_AGEMA_signal_1678 ), .Q ( new_AGEMA_signal_1679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_533 ( .C ( clk ), .D ( new_AGEMA_signal_1684 ), .Q ( new_AGEMA_signal_1685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_539 ( .C ( clk ), .D ( new_AGEMA_signal_1690 ), .Q ( new_AGEMA_signal_1691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_545 ( .C ( clk ), .D ( new_AGEMA_signal_1696 ), .Q ( new_AGEMA_signal_1697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_551 ( .C ( clk ), .D ( new_AGEMA_signal_1702 ), .Q ( new_AGEMA_signal_1703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_557 ( .C ( clk ), .D ( new_AGEMA_signal_1708 ), .Q ( new_AGEMA_signal_1709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_563 ( .C ( clk ), .D ( new_AGEMA_signal_1714 ), .Q ( new_AGEMA_signal_1715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_569 ( .C ( clk ), .D ( new_AGEMA_signal_1720 ), .Q ( new_AGEMA_signal_1721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_575 ( .C ( clk ), .D ( new_AGEMA_signal_1726 ), .Q ( new_AGEMA_signal_1727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_581 ( .C ( clk ), .D ( new_AGEMA_signal_1732 ), .Q ( new_AGEMA_signal_1733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_587 ( .C ( clk ), .D ( new_AGEMA_signal_1738 ), .Q ( new_AGEMA_signal_1739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_593 ( .C ( clk ), .D ( new_AGEMA_signal_1744 ), .Q ( new_AGEMA_signal_1745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_599 ( .C ( clk ), .D ( new_AGEMA_signal_1750 ), .Q ( new_AGEMA_signal_1751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_605 ( .C ( clk ), .D ( new_AGEMA_signal_1756 ), .Q ( new_AGEMA_signal_1757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_611 ( .C ( clk ), .D ( new_AGEMA_signal_1762 ), .Q ( new_AGEMA_signal_1763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_617 ( .C ( clk ), .D ( new_AGEMA_signal_1768 ), .Q ( new_AGEMA_signal_1769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_623 ( .C ( clk ), .D ( new_AGEMA_signal_1774 ), .Q ( new_AGEMA_signal_1775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_629 ( .C ( clk ), .D ( new_AGEMA_signal_1780 ), .Q ( new_AGEMA_signal_1781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_635 ( .C ( clk ), .D ( new_AGEMA_signal_1786 ), .Q ( new_AGEMA_signal_1787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_641 ( .C ( clk ), .D ( new_AGEMA_signal_1792 ), .Q ( new_AGEMA_signal_1793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_647 ( .C ( clk ), .D ( new_AGEMA_signal_1798 ), .Q ( new_AGEMA_signal_1799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_653 ( .C ( clk ), .D ( new_AGEMA_signal_1804 ), .Q ( new_AGEMA_signal_1805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_659 ( .C ( clk ), .D ( new_AGEMA_signal_1810 ), .Q ( new_AGEMA_signal_1811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_665 ( .C ( clk ), .D ( new_AGEMA_signal_1816 ), .Q ( new_AGEMA_signal_1817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_671 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_1823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_677 ( .C ( clk ), .D ( new_AGEMA_signal_1828 ), .Q ( new_AGEMA_signal_1829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_683 ( .C ( clk ), .D ( new_AGEMA_signal_1834 ), .Q ( new_AGEMA_signal_1835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_689 ( .C ( clk ), .D ( new_AGEMA_signal_1840 ), .Q ( new_AGEMA_signal_1841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_695 ( .C ( clk ), .D ( new_AGEMA_signal_1846 ), .Q ( new_AGEMA_signal_1847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_701 ( .C ( clk ), .D ( new_AGEMA_signal_1852 ), .Q ( new_AGEMA_signal_1853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_707 ( .C ( clk ), .D ( new_AGEMA_signal_1858 ), .Q ( new_AGEMA_signal_1859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_713 ( .C ( clk ), .D ( new_AGEMA_signal_1864 ), .Q ( new_AGEMA_signal_1865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_719 ( .C ( clk ), .D ( new_AGEMA_signal_1870 ), .Q ( new_AGEMA_signal_1871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_725 ( .C ( clk ), .D ( new_AGEMA_signal_1876 ), .Q ( new_AGEMA_signal_1877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_731 ( .C ( clk ), .D ( new_AGEMA_signal_1882 ), .Q ( new_AGEMA_signal_1883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_737 ( .C ( clk ), .D ( new_AGEMA_signal_1888 ), .Q ( new_AGEMA_signal_1889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_743 ( .C ( clk ), .D ( new_AGEMA_signal_1894 ), .Q ( new_AGEMA_signal_1895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_749 ( .C ( clk ), .D ( new_AGEMA_signal_1900 ), .Q ( new_AGEMA_signal_1901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_755 ( .C ( clk ), .D ( new_AGEMA_signal_1906 ), .Q ( new_AGEMA_signal_1907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_761 ( .C ( clk ), .D ( new_AGEMA_signal_1912 ), .Q ( new_AGEMA_signal_1913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_767 ( .C ( clk ), .D ( new_AGEMA_signal_1918 ), .Q ( new_AGEMA_signal_1919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_773 ( .C ( clk ), .D ( new_AGEMA_signal_1924 ), .Q ( new_AGEMA_signal_1925 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_240 ( .C ( clk ), .D ( new_AGEMA_signal_1391 ), .Q ( new_AGEMA_signal_1392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C ( clk ), .D ( new_AGEMA_signal_1397 ), .Q ( new_AGEMA_signal_1398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C ( clk ), .D ( new_AGEMA_signal_1403 ), .Q ( new_AGEMA_signal_1404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C ( clk ), .D ( new_AGEMA_signal_1409 ), .Q ( new_AGEMA_signal_1410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C ( clk ), .D ( new_AGEMA_signal_1415 ), .Q ( new_AGEMA_signal_1416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C ( clk ), .D ( new_AGEMA_signal_1421 ), .Q ( new_AGEMA_signal_1422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C ( clk ), .D ( new_AGEMA_signal_1427 ), .Q ( new_AGEMA_signal_1428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C ( clk ), .D ( new_AGEMA_signal_1433 ), .Q ( new_AGEMA_signal_1434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C ( clk ), .D ( new_AGEMA_signal_1439 ), .Q ( new_AGEMA_signal_1440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C ( clk ), .D ( new_AGEMA_signal_1445 ), .Q ( new_AGEMA_signal_1446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C ( clk ), .D ( new_AGEMA_signal_1451 ), .Q ( new_AGEMA_signal_1452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C ( clk ), .D ( new_AGEMA_signal_1457 ), .Q ( new_AGEMA_signal_1458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C ( clk ), .D ( new_AGEMA_signal_1463 ), .Q ( new_AGEMA_signal_1464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C ( clk ), .D ( new_AGEMA_signal_1469 ), .Q ( new_AGEMA_signal_1470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C ( clk ), .D ( new_AGEMA_signal_1475 ), .Q ( new_AGEMA_signal_1476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C ( clk ), .D ( new_AGEMA_signal_1481 ), .Q ( new_AGEMA_signal_1482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C ( clk ), .D ( new_AGEMA_signal_1487 ), .Q ( new_AGEMA_signal_1488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C ( clk ), .D ( new_AGEMA_signal_1493 ), .Q ( new_AGEMA_signal_1494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C ( clk ), .D ( new_AGEMA_signal_1499 ), .Q ( new_AGEMA_signal_1500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C ( clk ), .D ( new_AGEMA_signal_1505 ), .Q ( new_AGEMA_signal_1506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C ( clk ), .D ( new_AGEMA_signal_1511 ), .Q ( new_AGEMA_signal_1512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C ( clk ), .D ( new_AGEMA_signal_1517 ), .Q ( new_AGEMA_signal_1518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C ( clk ), .D ( new_AGEMA_signal_1523 ), .Q ( new_AGEMA_signal_1524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C ( clk ), .D ( new_AGEMA_signal_1529 ), .Q ( new_AGEMA_signal_1530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C ( clk ), .D ( new_AGEMA_signal_1535 ), .Q ( new_AGEMA_signal_1536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C ( clk ), .D ( new_AGEMA_signal_1541 ), .Q ( new_AGEMA_signal_1542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C ( clk ), .D ( new_AGEMA_signal_1547 ), .Q ( new_AGEMA_signal_1548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_402 ( .C ( clk ), .D ( new_AGEMA_signal_1553 ), .Q ( new_AGEMA_signal_1554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_408 ( .C ( clk ), .D ( new_AGEMA_signal_1559 ), .Q ( new_AGEMA_signal_1560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_414 ( .C ( clk ), .D ( new_AGEMA_signal_1565 ), .Q ( new_AGEMA_signal_1566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_420 ( .C ( clk ), .D ( new_AGEMA_signal_1571 ), .Q ( new_AGEMA_signal_1572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_426 ( .C ( clk ), .D ( new_AGEMA_signal_1577 ), .Q ( new_AGEMA_signal_1578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_432 ( .C ( clk ), .D ( new_AGEMA_signal_1583 ), .Q ( new_AGEMA_signal_1584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_438 ( .C ( clk ), .D ( new_AGEMA_signal_1589 ), .Q ( new_AGEMA_signal_1590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_444 ( .C ( clk ), .D ( new_AGEMA_signal_1595 ), .Q ( new_AGEMA_signal_1596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_450 ( .C ( clk ), .D ( new_AGEMA_signal_1601 ), .Q ( new_AGEMA_signal_1602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_456 ( .C ( clk ), .D ( new_AGEMA_signal_1607 ), .Q ( new_AGEMA_signal_1608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_462 ( .C ( clk ), .D ( new_AGEMA_signal_1613 ), .Q ( new_AGEMA_signal_1614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_468 ( .C ( clk ), .D ( new_AGEMA_signal_1619 ), .Q ( new_AGEMA_signal_1620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_474 ( .C ( clk ), .D ( new_AGEMA_signal_1625 ), .Q ( new_AGEMA_signal_1626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_480 ( .C ( clk ), .D ( new_AGEMA_signal_1631 ), .Q ( new_AGEMA_signal_1632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_486 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_1638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_492 ( .C ( clk ), .D ( new_AGEMA_signal_1643 ), .Q ( new_AGEMA_signal_1644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_498 ( .C ( clk ), .D ( new_AGEMA_signal_1649 ), .Q ( new_AGEMA_signal_1650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_504 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_1656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_510 ( .C ( clk ), .D ( new_AGEMA_signal_1661 ), .Q ( new_AGEMA_signal_1662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_516 ( .C ( clk ), .D ( new_AGEMA_signal_1667 ), .Q ( new_AGEMA_signal_1668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_522 ( .C ( clk ), .D ( new_AGEMA_signal_1673 ), .Q ( new_AGEMA_signal_1674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_528 ( .C ( clk ), .D ( new_AGEMA_signal_1679 ), .Q ( new_AGEMA_signal_1680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_534 ( .C ( clk ), .D ( new_AGEMA_signal_1685 ), .Q ( new_AGEMA_signal_1686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_540 ( .C ( clk ), .D ( new_AGEMA_signal_1691 ), .Q ( new_AGEMA_signal_1692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_546 ( .C ( clk ), .D ( new_AGEMA_signal_1697 ), .Q ( new_AGEMA_signal_1698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_552 ( .C ( clk ), .D ( new_AGEMA_signal_1703 ), .Q ( new_AGEMA_signal_1704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_558 ( .C ( clk ), .D ( new_AGEMA_signal_1709 ), .Q ( new_AGEMA_signal_1710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_564 ( .C ( clk ), .D ( new_AGEMA_signal_1715 ), .Q ( new_AGEMA_signal_1716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_570 ( .C ( clk ), .D ( new_AGEMA_signal_1721 ), .Q ( new_AGEMA_signal_1722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_576 ( .C ( clk ), .D ( new_AGEMA_signal_1727 ), .Q ( new_AGEMA_signal_1728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_582 ( .C ( clk ), .D ( new_AGEMA_signal_1733 ), .Q ( new_AGEMA_signal_1734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_588 ( .C ( clk ), .D ( new_AGEMA_signal_1739 ), .Q ( new_AGEMA_signal_1740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_594 ( .C ( clk ), .D ( new_AGEMA_signal_1745 ), .Q ( new_AGEMA_signal_1746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_600 ( .C ( clk ), .D ( new_AGEMA_signal_1751 ), .Q ( new_AGEMA_signal_1752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_606 ( .C ( clk ), .D ( new_AGEMA_signal_1757 ), .Q ( new_AGEMA_signal_1758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_612 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_1764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_618 ( .C ( clk ), .D ( new_AGEMA_signal_1769 ), .Q ( new_AGEMA_signal_1770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_624 ( .C ( clk ), .D ( new_AGEMA_signal_1775 ), .Q ( new_AGEMA_signal_1776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_630 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_1782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_636 ( .C ( clk ), .D ( new_AGEMA_signal_1787 ), .Q ( new_AGEMA_signal_1788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_642 ( .C ( clk ), .D ( new_AGEMA_signal_1793 ), .Q ( new_AGEMA_signal_1794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_648 ( .C ( clk ), .D ( new_AGEMA_signal_1799 ), .Q ( new_AGEMA_signal_1800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_654 ( .C ( clk ), .D ( new_AGEMA_signal_1805 ), .Q ( new_AGEMA_signal_1806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_660 ( .C ( clk ), .D ( new_AGEMA_signal_1811 ), .Q ( new_AGEMA_signal_1812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_666 ( .C ( clk ), .D ( new_AGEMA_signal_1817 ), .Q ( new_AGEMA_signal_1818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_672 ( .C ( clk ), .D ( new_AGEMA_signal_1823 ), .Q ( new_AGEMA_signal_1824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_678 ( .C ( clk ), .D ( new_AGEMA_signal_1829 ), .Q ( new_AGEMA_signal_1830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_684 ( .C ( clk ), .D ( new_AGEMA_signal_1835 ), .Q ( new_AGEMA_signal_1836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_690 ( .C ( clk ), .D ( new_AGEMA_signal_1841 ), .Q ( new_AGEMA_signal_1842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_696 ( .C ( clk ), .D ( new_AGEMA_signal_1847 ), .Q ( new_AGEMA_signal_1848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_702 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_1854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_708 ( .C ( clk ), .D ( new_AGEMA_signal_1859 ), .Q ( new_AGEMA_signal_1860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_714 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_1866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_720 ( .C ( clk ), .D ( new_AGEMA_signal_1871 ), .Q ( new_AGEMA_signal_1872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_726 ( .C ( clk ), .D ( new_AGEMA_signal_1877 ), .Q ( new_AGEMA_signal_1878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_732 ( .C ( clk ), .D ( new_AGEMA_signal_1883 ), .Q ( new_AGEMA_signal_1884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_738 ( .C ( clk ), .D ( new_AGEMA_signal_1889 ), .Q ( new_AGEMA_signal_1890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_744 ( .C ( clk ), .D ( new_AGEMA_signal_1895 ), .Q ( new_AGEMA_signal_1896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_750 ( .C ( clk ), .D ( new_AGEMA_signal_1901 ), .Q ( new_AGEMA_signal_1902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_756 ( .C ( clk ), .D ( new_AGEMA_signal_1907 ), .Q ( new_AGEMA_signal_1908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_762 ( .C ( clk ), .D ( new_AGEMA_signal_1913 ), .Q ( new_AGEMA_signal_1914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_768 ( .C ( clk ), .D ( new_AGEMA_signal_1919 ), .Q ( new_AGEMA_signal_1920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_774 ( .C ( clk ), .D ( new_AGEMA_signal_1925 ), .Q ( new_AGEMA_signal_1926 ) ) ;

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U39 ( .a ({new_AGEMA_signal_583, new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, sbe_inv_d_0_}), .b ({new_AGEMA_signal_579, new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_d_1_}), .c ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, sbe_inv_dl}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U38 ( .a ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, sbe_inv_d_2_}), .b ({new_AGEMA_signal_571, new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, sbe_inv_d_3_}), .c ({new_AGEMA_signal_591, new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_inv_dh}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U37 ( .a ({new_AGEMA_signal_595, new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, sbe_inv_sd_1_}), .c ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, sbe_inv_dd}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U36 ( .a ({new_AGEMA_signal_583, new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, sbe_inv_d_0_}), .b ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, sbe_inv_d_2_}), .c ({new_AGEMA_signal_595, new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, sbe_inv_sd_0_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_U35 ( .a ({new_AGEMA_signal_579, new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_d_1_}), .b ({new_AGEMA_signal_571, new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, sbe_inv_d_3_}), .c ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, sbe_inv_sd_1_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_pmul_U5 ( .a ({new_AGEMA_signal_563, new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_547, new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, sbe_inv_dinv_pmul_n8}), .c ({new_AGEMA_signal_571, new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, sbe_inv_d_3_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_pmul_U4 ( .a ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1335, new_AGEMA_signal_1333, new_AGEMA_signal_1331, new_AGEMA_signal_1329}), .clk ( clk ), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_547, new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, sbe_inv_dinv_pmul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_pmul_U3 ( .a ({new_AGEMA_signal_563, new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_551, new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, sbe_inv_dinv_pmul_n7}), .c ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, sbe_inv_d_2_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_pmul_U2 ( .a ({new_AGEMA_signal_535, new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1345, new_AGEMA_signal_1343, new_AGEMA_signal_1341, new_AGEMA_signal_1339}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({new_AGEMA_signal_551, new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, sbe_inv_dinv_pmul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_pmul_U1 ( .a ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1355, new_AGEMA_signal_1353, new_AGEMA_signal_1351, new_AGEMA_signal_1349}), .clk ( clk ), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_563, new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, sbe_inv_dinv_pmul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_qmul_U5 ( .a ({new_AGEMA_signal_567, new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, sbe_inv_dinv_qmul_n8}), .c ({new_AGEMA_signal_579, new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_d_1_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_qmul_U4 ( .a ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1365, new_AGEMA_signal_1363, new_AGEMA_signal_1361, new_AGEMA_signal_1359}), .clk ( clk ), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, sbe_inv_dinv_qmul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_qmul_U3 ( .a ({new_AGEMA_signal_567, new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_559, new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, sbe_inv_dinv_qmul_n7}), .c ({new_AGEMA_signal_583, new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, sbe_inv_d_0_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_qmul_U2 ( .a ({new_AGEMA_signal_535, new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1375, new_AGEMA_signal_1373, new_AGEMA_signal_1371, new_AGEMA_signal_1369}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_559, new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, sbe_inv_dinv_qmul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_dinv_qmul_U1 ( .a ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1385, new_AGEMA_signal_1383, new_AGEMA_signal_1381, new_AGEMA_signal_1379}), .clk ( clk ), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_567, new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_dinv_qmul_n9}) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C ( clk ), .D ( new_AGEMA_signal_1392 ), .Q ( new_AGEMA_signal_1393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C ( clk ), .D ( new_AGEMA_signal_1398 ), .Q ( new_AGEMA_signal_1399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C ( clk ), .D ( new_AGEMA_signal_1404 ), .Q ( new_AGEMA_signal_1405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C ( clk ), .D ( new_AGEMA_signal_1410 ), .Q ( new_AGEMA_signal_1411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C ( clk ), .D ( new_AGEMA_signal_1416 ), .Q ( new_AGEMA_signal_1417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C ( clk ), .D ( new_AGEMA_signal_1422 ), .Q ( new_AGEMA_signal_1423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C ( clk ), .D ( new_AGEMA_signal_1428 ), .Q ( new_AGEMA_signal_1429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C ( clk ), .D ( new_AGEMA_signal_1434 ), .Q ( new_AGEMA_signal_1435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C ( clk ), .D ( new_AGEMA_signal_1440 ), .Q ( new_AGEMA_signal_1441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_1447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C ( clk ), .D ( new_AGEMA_signal_1452 ), .Q ( new_AGEMA_signal_1453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C ( clk ), .D ( new_AGEMA_signal_1458 ), .Q ( new_AGEMA_signal_1459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C ( clk ), .D ( new_AGEMA_signal_1464 ), .Q ( new_AGEMA_signal_1465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C ( clk ), .D ( new_AGEMA_signal_1470 ), .Q ( new_AGEMA_signal_1471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C ( clk ), .D ( new_AGEMA_signal_1476 ), .Q ( new_AGEMA_signal_1477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_1483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C ( clk ), .D ( new_AGEMA_signal_1488 ), .Q ( new_AGEMA_signal_1489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C ( clk ), .D ( new_AGEMA_signal_1494 ), .Q ( new_AGEMA_signal_1495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C ( clk ), .D ( new_AGEMA_signal_1500 ), .Q ( new_AGEMA_signal_1501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C ( clk ), .D ( new_AGEMA_signal_1506 ), .Q ( new_AGEMA_signal_1507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C ( clk ), .D ( new_AGEMA_signal_1512 ), .Q ( new_AGEMA_signal_1513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C ( clk ), .D ( new_AGEMA_signal_1518 ), .Q ( new_AGEMA_signal_1519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C ( clk ), .D ( new_AGEMA_signal_1524 ), .Q ( new_AGEMA_signal_1525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C ( clk ), .D ( new_AGEMA_signal_1530 ), .Q ( new_AGEMA_signal_1531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C ( clk ), .D ( new_AGEMA_signal_1536 ), .Q ( new_AGEMA_signal_1537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C ( clk ), .D ( new_AGEMA_signal_1542 ), .Q ( new_AGEMA_signal_1543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C ( clk ), .D ( new_AGEMA_signal_1548 ), .Q ( new_AGEMA_signal_1549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_403 ( .C ( clk ), .D ( new_AGEMA_signal_1554 ), .Q ( new_AGEMA_signal_1555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_409 ( .C ( clk ), .D ( new_AGEMA_signal_1560 ), .Q ( new_AGEMA_signal_1561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_415 ( .C ( clk ), .D ( new_AGEMA_signal_1566 ), .Q ( new_AGEMA_signal_1567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_421 ( .C ( clk ), .D ( new_AGEMA_signal_1572 ), .Q ( new_AGEMA_signal_1573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_427 ( .C ( clk ), .D ( new_AGEMA_signal_1578 ), .Q ( new_AGEMA_signal_1579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_433 ( .C ( clk ), .D ( new_AGEMA_signal_1584 ), .Q ( new_AGEMA_signal_1585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_439 ( .C ( clk ), .D ( new_AGEMA_signal_1590 ), .Q ( new_AGEMA_signal_1591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_445 ( .C ( clk ), .D ( new_AGEMA_signal_1596 ), .Q ( new_AGEMA_signal_1597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_451 ( .C ( clk ), .D ( new_AGEMA_signal_1602 ), .Q ( new_AGEMA_signal_1603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_457 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_1609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_463 ( .C ( clk ), .D ( new_AGEMA_signal_1614 ), .Q ( new_AGEMA_signal_1615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_469 ( .C ( clk ), .D ( new_AGEMA_signal_1620 ), .Q ( new_AGEMA_signal_1621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_475 ( .C ( clk ), .D ( new_AGEMA_signal_1626 ), .Q ( new_AGEMA_signal_1627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_481 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_1633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_487 ( .C ( clk ), .D ( new_AGEMA_signal_1638 ), .Q ( new_AGEMA_signal_1639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_493 ( .C ( clk ), .D ( new_AGEMA_signal_1644 ), .Q ( new_AGEMA_signal_1645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_499 ( .C ( clk ), .D ( new_AGEMA_signal_1650 ), .Q ( new_AGEMA_signal_1651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_505 ( .C ( clk ), .D ( new_AGEMA_signal_1656 ), .Q ( new_AGEMA_signal_1657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_511 ( .C ( clk ), .D ( new_AGEMA_signal_1662 ), .Q ( new_AGEMA_signal_1663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_517 ( .C ( clk ), .D ( new_AGEMA_signal_1668 ), .Q ( new_AGEMA_signal_1669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_523 ( .C ( clk ), .D ( new_AGEMA_signal_1674 ), .Q ( new_AGEMA_signal_1675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_529 ( .C ( clk ), .D ( new_AGEMA_signal_1680 ), .Q ( new_AGEMA_signal_1681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_535 ( .C ( clk ), .D ( new_AGEMA_signal_1686 ), .Q ( new_AGEMA_signal_1687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_541 ( .C ( clk ), .D ( new_AGEMA_signal_1692 ), .Q ( new_AGEMA_signal_1693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_547 ( .C ( clk ), .D ( new_AGEMA_signal_1698 ), .Q ( new_AGEMA_signal_1699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_553 ( .C ( clk ), .D ( new_AGEMA_signal_1704 ), .Q ( new_AGEMA_signal_1705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_559 ( .C ( clk ), .D ( new_AGEMA_signal_1710 ), .Q ( new_AGEMA_signal_1711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_565 ( .C ( clk ), .D ( new_AGEMA_signal_1716 ), .Q ( new_AGEMA_signal_1717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_571 ( .C ( clk ), .D ( new_AGEMA_signal_1722 ), .Q ( new_AGEMA_signal_1723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_577 ( .C ( clk ), .D ( new_AGEMA_signal_1728 ), .Q ( new_AGEMA_signal_1729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_583 ( .C ( clk ), .D ( new_AGEMA_signal_1734 ), .Q ( new_AGEMA_signal_1735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_589 ( .C ( clk ), .D ( new_AGEMA_signal_1740 ), .Q ( new_AGEMA_signal_1741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_595 ( .C ( clk ), .D ( new_AGEMA_signal_1746 ), .Q ( new_AGEMA_signal_1747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_601 ( .C ( clk ), .D ( new_AGEMA_signal_1752 ), .Q ( new_AGEMA_signal_1753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_607 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_1759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_613 ( .C ( clk ), .D ( new_AGEMA_signal_1764 ), .Q ( new_AGEMA_signal_1765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_619 ( .C ( clk ), .D ( new_AGEMA_signal_1770 ), .Q ( new_AGEMA_signal_1771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_625 ( .C ( clk ), .D ( new_AGEMA_signal_1776 ), .Q ( new_AGEMA_signal_1777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_631 ( .C ( clk ), .D ( new_AGEMA_signal_1782 ), .Q ( new_AGEMA_signal_1783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_637 ( .C ( clk ), .D ( new_AGEMA_signal_1788 ), .Q ( new_AGEMA_signal_1789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_643 ( .C ( clk ), .D ( new_AGEMA_signal_1794 ), .Q ( new_AGEMA_signal_1795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_649 ( .C ( clk ), .D ( new_AGEMA_signal_1800 ), .Q ( new_AGEMA_signal_1801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_655 ( .C ( clk ), .D ( new_AGEMA_signal_1806 ), .Q ( new_AGEMA_signal_1807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_661 ( .C ( clk ), .D ( new_AGEMA_signal_1812 ), .Q ( new_AGEMA_signal_1813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_667 ( .C ( clk ), .D ( new_AGEMA_signal_1818 ), .Q ( new_AGEMA_signal_1819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_673 ( .C ( clk ), .D ( new_AGEMA_signal_1824 ), .Q ( new_AGEMA_signal_1825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_679 ( .C ( clk ), .D ( new_AGEMA_signal_1830 ), .Q ( new_AGEMA_signal_1831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_685 ( .C ( clk ), .D ( new_AGEMA_signal_1836 ), .Q ( new_AGEMA_signal_1837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_691 ( .C ( clk ), .D ( new_AGEMA_signal_1842 ), .Q ( new_AGEMA_signal_1843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_697 ( .C ( clk ), .D ( new_AGEMA_signal_1848 ), .Q ( new_AGEMA_signal_1849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_703 ( .C ( clk ), .D ( new_AGEMA_signal_1854 ), .Q ( new_AGEMA_signal_1855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_709 ( .C ( clk ), .D ( new_AGEMA_signal_1860 ), .Q ( new_AGEMA_signal_1861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_715 ( .C ( clk ), .D ( new_AGEMA_signal_1866 ), .Q ( new_AGEMA_signal_1867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_721 ( .C ( clk ), .D ( new_AGEMA_signal_1872 ), .Q ( new_AGEMA_signal_1873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_727 ( .C ( clk ), .D ( new_AGEMA_signal_1878 ), .Q ( new_AGEMA_signal_1879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_733 ( .C ( clk ), .D ( new_AGEMA_signal_1884 ), .Q ( new_AGEMA_signal_1885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_739 ( .C ( clk ), .D ( new_AGEMA_signal_1890 ), .Q ( new_AGEMA_signal_1891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_745 ( .C ( clk ), .D ( new_AGEMA_signal_1896 ), .Q ( new_AGEMA_signal_1897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_751 ( .C ( clk ), .D ( new_AGEMA_signal_1902 ), .Q ( new_AGEMA_signal_1903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_757 ( .C ( clk ), .D ( new_AGEMA_signal_1908 ), .Q ( new_AGEMA_signal_1909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_763 ( .C ( clk ), .D ( new_AGEMA_signal_1914 ), .Q ( new_AGEMA_signal_1915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_769 ( .C ( clk ), .D ( new_AGEMA_signal_1920 ), .Q ( new_AGEMA_signal_1921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_775 ( .C ( clk ), .D ( new_AGEMA_signal_1926 ), .Q ( new_AGEMA_signal_1927 ) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    not_masked #(.security_order(4), .pipeline(1)) sbe_U40 ( .a ({new_AGEMA_signal_731, new_AGEMA_signal_730, new_AGEMA_signal_729, new_AGEMA_signal_728, sbe_C_2_}), .b ({new_AGEMA_signal_743, new_AGEMA_signal_742, new_AGEMA_signal_741, new_AGEMA_signal_740, sbe_n1}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U34 ( .a ({new_AGEMA_signal_755, new_AGEMA_signal_754, new_AGEMA_signal_753, new_AGEMA_signal_752, sbe_C_7_}), .b ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, new_AGEMA_signal_792, sbe_n17}), .c ({new_AGEMA_signal_815, new_AGEMA_signal_814, new_AGEMA_signal_813, new_AGEMA_signal_812, sbe_n16}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U33 ( .a ({new_AGEMA_signal_723, new_AGEMA_signal_722, new_AGEMA_signal_721, new_AGEMA_signal_720, sbe_C_4_}), .b ({new_AGEMA_signal_771, new_AGEMA_signal_770, new_AGEMA_signal_769, new_AGEMA_signal_768, sbe_n18}), .c ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, new_AGEMA_signal_792, sbe_n17}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U32 ( .a ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, new_AGEMA_signal_756, sbe_C_5_}), .b ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}), .c ({new_AGEMA_signal_771, new_AGEMA_signal_770, new_AGEMA_signal_769, new_AGEMA_signal_768, sbe_n18}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U31 ( .a ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}), .b ({new_AGEMA_signal_723, new_AGEMA_signal_722, new_AGEMA_signal_721, new_AGEMA_signal_720, sbe_C_4_}), .c ({new_AGEMA_signal_775, new_AGEMA_signal_774, new_AGEMA_signal_773, new_AGEMA_signal_772, sbe_n15}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U30 ( .a ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, new_AGEMA_signal_716, sbe_C_6_}), .b ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}), .c ({new_AGEMA_signal_779, new_AGEMA_signal_778, new_AGEMA_signal_777, new_AGEMA_signal_776, sbe_n14}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U21 ( .a ({new_AGEMA_signal_819, new_AGEMA_signal_818, new_AGEMA_signal_817, new_AGEMA_signal_816, sbe_n6}), .b ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}), .c ({new_AGEMA_signal_851, new_AGEMA_signal_850, new_AGEMA_signal_849, new_AGEMA_signal_848, sbe_X[6]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U20 ( .a ({new_AGEMA_signal_731, new_AGEMA_signal_730, new_AGEMA_signal_729, new_AGEMA_signal_728, sbe_C_2_}), .b ({new_AGEMA_signal_819, new_AGEMA_signal_818, new_AGEMA_signal_817, new_AGEMA_signal_816, sbe_n6}), .c ({new_AGEMA_signal_855, new_AGEMA_signal_854, new_AGEMA_signal_853, new_AGEMA_signal_852, sbe_X[5]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U19 ( .a ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, new_AGEMA_signal_744, sbe_D_5_}), .b ({new_AGEMA_signal_799, new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, sbe_n20}), .c ({new_AGEMA_signal_819, new_AGEMA_signal_818, new_AGEMA_signal_817, new_AGEMA_signal_816, sbe_n6}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U18 ( .a ({new_AGEMA_signal_803, new_AGEMA_signal_802, new_AGEMA_signal_801, new_AGEMA_signal_800, sbe_n5}), .b ({new_AGEMA_signal_791, new_AGEMA_signal_790, new_AGEMA_signal_789, new_AGEMA_signal_788, sbe_D_0_}), .c ({new_AGEMA_signal_823, new_AGEMA_signal_822, new_AGEMA_signal_821, new_AGEMA_signal_820, sbe_X[3]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U17 ( .a ({new_AGEMA_signal_799, new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, sbe_n20}), .b ({new_AGEMA_signal_751, new_AGEMA_signal_750, new_AGEMA_signal_749, new_AGEMA_signal_748, sbe_n4}), .c ({new_AGEMA_signal_827, new_AGEMA_signal_826, new_AGEMA_signal_825, new_AGEMA_signal_824, sbe_D_3_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U16 ( .a ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, new_AGEMA_signal_756, sbe_C_5_}), .b ({new_AGEMA_signal_783, new_AGEMA_signal_782, new_AGEMA_signal_781, new_AGEMA_signal_780, sbe_D_6_}), .c ({new_AGEMA_signal_799, new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, sbe_n20}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U15 ( .a ({new_AGEMA_signal_755, new_AGEMA_signal_754, new_AGEMA_signal_753, new_AGEMA_signal_752, sbe_C_7_}), .b ({new_AGEMA_signal_763, new_AGEMA_signal_762, new_AGEMA_signal_761, new_AGEMA_signal_760, sbe_C_3_}), .c ({new_AGEMA_signal_783, new_AGEMA_signal_782, new_AGEMA_signal_781, new_AGEMA_signal_780, sbe_D_6_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U14 ( .a ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, new_AGEMA_signal_744, sbe_D_5_}), .b ({new_AGEMA_signal_803, new_AGEMA_signal_802, new_AGEMA_signal_801, new_AGEMA_signal_800, sbe_n5}), .c ({new_AGEMA_signal_831, new_AGEMA_signal_830, new_AGEMA_signal_829, new_AGEMA_signal_828, sbe_D_2_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U13 ( .a ({new_AGEMA_signal_731, new_AGEMA_signal_730, new_AGEMA_signal_729, new_AGEMA_signal_728, sbe_C_2_}), .b ({new_AGEMA_signal_787, new_AGEMA_signal_786, new_AGEMA_signal_785, new_AGEMA_signal_784, sbe_n19}), .c ({new_AGEMA_signal_803, new_AGEMA_signal_802, new_AGEMA_signal_801, new_AGEMA_signal_800, sbe_n5}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U12 ( .a ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, new_AGEMA_signal_756, sbe_C_5_}), .b ({new_AGEMA_signal_763, new_AGEMA_signal_762, new_AGEMA_signal_761, new_AGEMA_signal_760, sbe_C_3_}), .c ({new_AGEMA_signal_787, new_AGEMA_signal_786, new_AGEMA_signal_785, new_AGEMA_signal_784, sbe_n19}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U11 ( .a ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, new_AGEMA_signal_716, sbe_C_6_}), .b ({new_AGEMA_signal_735, new_AGEMA_signal_734, new_AGEMA_signal_733, new_AGEMA_signal_732, sbe_C_0_}), .c ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, new_AGEMA_signal_744, sbe_D_5_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U10 ( .a ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}), .b ({new_AGEMA_signal_751, new_AGEMA_signal_750, new_AGEMA_signal_749, new_AGEMA_signal_748, sbe_n4}), .c ({new_AGEMA_signal_791, new_AGEMA_signal_790, new_AGEMA_signal_789, new_AGEMA_signal_788, sbe_D_0_}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) sbe_U9 ( .a ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, new_AGEMA_signal_716, sbe_C_6_}), .b ({new_AGEMA_signal_723, new_AGEMA_signal_722, new_AGEMA_signal_721, new_AGEMA_signal_720, sbe_C_4_}), .c ({new_AGEMA_signal_751, new_AGEMA_signal_750, new_AGEMA_signal_749, new_AGEMA_signal_748, sbe_n4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_U4 ( .a ({new_AGEMA_signal_727, new_AGEMA_signal_726, new_AGEMA_signal_725, new_AGEMA_signal_724, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_671, new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, sbe_inv_pmul_ph[1]}), .c ({new_AGEMA_signal_755, new_AGEMA_signal_754, new_AGEMA_signal_753, new_AGEMA_signal_752, sbe_C_7_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_U3 ( .a ({new_AGEMA_signal_691, new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_675, new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, sbe_inv_pmul_ph[0]}), .c ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, new_AGEMA_signal_716, sbe_C_6_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_U2 ( .a ({new_AGEMA_signal_727, new_AGEMA_signal_726, new_AGEMA_signal_725, new_AGEMA_signal_724, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_679, new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, sbe_inv_pmul_pl[1]}), .c ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, new_AGEMA_signal_756, sbe_C_5_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_U1 ( .a ({new_AGEMA_signal_691, new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_683, new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, sbe_inv_pmul_pl[0]}), .c ({new_AGEMA_signal_723, new_AGEMA_signal_722, new_AGEMA_signal_721, new_AGEMA_signal_720, sbe_C_4_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_himul_U5 ( .a ({new_AGEMA_signal_639, new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_603, new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, sbe_inv_pmul_himul_n8}), .c ({new_AGEMA_signal_671, new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, sbe_inv_pmul_ph[1]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_himul_U4 ( .a ({new_AGEMA_signal_571, new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, sbe_inv_d_3_}), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1411, new_AGEMA_signal_1405, new_AGEMA_signal_1399, new_AGEMA_signal_1393}), .clk ( clk ), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_603, new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, sbe_inv_pmul_himul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_himul_U3 ( .a ({new_AGEMA_signal_639, new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_607, new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, sbe_inv_pmul_himul_n7}), .c ({new_AGEMA_signal_675, new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, sbe_inv_pmul_ph[0]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_himul_U2 ( .a ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, sbe_inv_d_2_}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1441, new_AGEMA_signal_1435, new_AGEMA_signal_1429, new_AGEMA_signal_1423}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({new_AGEMA_signal_607, new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, sbe_inv_pmul_himul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_himul_U1 ( .a ({new_AGEMA_signal_591, new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_inv_dh}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1471, new_AGEMA_signal_1465, new_AGEMA_signal_1459, new_AGEMA_signal_1453}), .clk ( clk ), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_639, new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_inv_pmul_himul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_lomul_U5 ( .a ({new_AGEMA_signal_643, new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_611, new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, sbe_inv_pmul_lomul_n8}), .c ({new_AGEMA_signal_679, new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, sbe_inv_pmul_pl[1]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_lomul_U4 ( .a ({new_AGEMA_signal_579, new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_d_1_}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1501, new_AGEMA_signal_1495, new_AGEMA_signal_1489, new_AGEMA_signal_1483}), .clk ( clk ), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({new_AGEMA_signal_611, new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, sbe_inv_pmul_lomul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_lomul_U3 ( .a ({new_AGEMA_signal_643, new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_615, new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, sbe_inv_pmul_lomul_n7}), .c ({new_AGEMA_signal_683, new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, sbe_inv_pmul_pl[0]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_lomul_U2 ( .a ({new_AGEMA_signal_583, new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, sbe_inv_d_0_}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1531, new_AGEMA_signal_1525, new_AGEMA_signal_1519, new_AGEMA_signal_1513}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_615, new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, sbe_inv_pmul_lomul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_lomul_U1 ( .a ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, sbe_inv_dl}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1561, new_AGEMA_signal_1555, new_AGEMA_signal_1549, new_AGEMA_signal_1543}), .clk ( clk ), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_643, new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, sbe_inv_pmul_lomul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_summul_U5 ( .a ({new_AGEMA_signal_651, new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_687, new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, sbe_inv_pmul_summul_n8}), .c ({new_AGEMA_signal_727, new_AGEMA_signal_726, new_AGEMA_signal_725, new_AGEMA_signal_724, sbe_inv_pmul_p_1_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_summul_U4 ( .a ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, sbe_inv_dd}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1591, new_AGEMA_signal_1585, new_AGEMA_signal_1579, new_AGEMA_signal_1573}), .clk ( clk ), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({new_AGEMA_signal_687, new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, sbe_inv_pmul_summul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_summul_U3 ( .a ({new_AGEMA_signal_651, new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, sbe_inv_pmul_summul_n7}), .c ({new_AGEMA_signal_691, new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, sbe_inv_pmul_p_0_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_summul_U2 ( .a ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1621, new_AGEMA_signal_1615, new_AGEMA_signal_1609, new_AGEMA_signal_1603}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, sbe_inv_pmul_summul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_pmul_summul_U1 ( .a ({new_AGEMA_signal_595, new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1651, new_AGEMA_signal_1645, new_AGEMA_signal_1639, new_AGEMA_signal_1633}), .clk ( clk ), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_651, new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_inv_pmul_summul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_U4 ( .a ({new_AGEMA_signal_739, new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_695, new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, sbe_inv_qmul_ph[1]}), .c ({new_AGEMA_signal_763, new_AGEMA_signal_762, new_AGEMA_signal_761, new_AGEMA_signal_760, sbe_C_3_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_U3 ( .a ({new_AGEMA_signal_715, new_AGEMA_signal_714, new_AGEMA_signal_713, new_AGEMA_signal_712, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_699, new_AGEMA_signal_698, new_AGEMA_signal_697, new_AGEMA_signal_696, sbe_inv_qmul_ph[0]}), .c ({new_AGEMA_signal_731, new_AGEMA_signal_730, new_AGEMA_signal_729, new_AGEMA_signal_728, sbe_C_2_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_U2 ( .a ({new_AGEMA_signal_739, new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_703, new_AGEMA_signal_702, new_AGEMA_signal_701, new_AGEMA_signal_700, sbe_inv_qmul_pl[1]}), .c ({new_AGEMA_signal_767, new_AGEMA_signal_766, new_AGEMA_signal_765, new_AGEMA_signal_764, sbe_C_1_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_U1 ( .a ({new_AGEMA_signal_715, new_AGEMA_signal_714, new_AGEMA_signal_713, new_AGEMA_signal_712, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_707, new_AGEMA_signal_706, new_AGEMA_signal_705, new_AGEMA_signal_704, sbe_inv_qmul_pl[0]}), .c ({new_AGEMA_signal_735, new_AGEMA_signal_734, new_AGEMA_signal_733, new_AGEMA_signal_732, sbe_C_0_}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_himul_U5 ( .a ({new_AGEMA_signal_655, new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_619, new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, sbe_inv_qmul_himul_n8}), .c ({new_AGEMA_signal_695, new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, sbe_inv_qmul_ph[1]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_himul_U4 ( .a ({new_AGEMA_signal_571, new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, sbe_inv_d_3_}), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1681, new_AGEMA_signal_1675, new_AGEMA_signal_1669, new_AGEMA_signal_1663}), .clk ( clk ), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({new_AGEMA_signal_619, new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, sbe_inv_qmul_himul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_himul_U3 ( .a ({new_AGEMA_signal_655, new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, sbe_inv_qmul_himul_n7}), .c ({new_AGEMA_signal_699, new_AGEMA_signal_698, new_AGEMA_signal_697, new_AGEMA_signal_696, sbe_inv_qmul_ph[0]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_himul_U2 ( .a ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, sbe_inv_d_2_}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1711, new_AGEMA_signal_1705, new_AGEMA_signal_1699, new_AGEMA_signal_1693}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, sbe_inv_qmul_himul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_himul_U1 ( .a ({new_AGEMA_signal_591, new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_inv_dh}), .b ({new_AGEMA_signal_1747, new_AGEMA_signal_1741, new_AGEMA_signal_1735, new_AGEMA_signal_1729, new_AGEMA_signal_1723}), .clk ( clk ), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_655, new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, sbe_inv_qmul_himul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_lomul_U5 ( .a ({new_AGEMA_signal_659, new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_627, new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, sbe_inv_qmul_lomul_n8}), .c ({new_AGEMA_signal_703, new_AGEMA_signal_702, new_AGEMA_signal_701, new_AGEMA_signal_700, sbe_inv_qmul_pl[1]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_lomul_U4 ( .a ({new_AGEMA_signal_579, new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_d_1_}), .b ({new_AGEMA_signal_1777, new_AGEMA_signal_1771, new_AGEMA_signal_1765, new_AGEMA_signal_1759, new_AGEMA_signal_1753}), .clk ( clk ), .r ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({new_AGEMA_signal_627, new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, sbe_inv_qmul_lomul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_lomul_U3 ( .a ({new_AGEMA_signal_659, new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_631, new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, sbe_inv_qmul_lomul_n7}), .c ({new_AGEMA_signal_707, new_AGEMA_signal_706, new_AGEMA_signal_705, new_AGEMA_signal_704, sbe_inv_qmul_pl[0]}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_lomul_U2 ( .a ({new_AGEMA_signal_583, new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, sbe_inv_d_0_}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1801, new_AGEMA_signal_1795, new_AGEMA_signal_1789, new_AGEMA_signal_1783}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .c ({new_AGEMA_signal_631, new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, sbe_inv_qmul_lomul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_lomul_U1 ( .a ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, sbe_inv_dl}), .b ({new_AGEMA_signal_1837, new_AGEMA_signal_1831, new_AGEMA_signal_1825, new_AGEMA_signal_1819, new_AGEMA_signal_1813}), .clk ( clk ), .r ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_659, new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, sbe_inv_qmul_lomul_n9}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_summul_U5 ( .a ({new_AGEMA_signal_667, new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_711, new_AGEMA_signal_710, new_AGEMA_signal_709, new_AGEMA_signal_708, sbe_inv_qmul_summul_n8}), .c ({new_AGEMA_signal_739, new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, sbe_inv_qmul_p_1_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_summul_U4 ( .a ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, sbe_inv_dd}), .b ({new_AGEMA_signal_1867, new_AGEMA_signal_1861, new_AGEMA_signal_1855, new_AGEMA_signal_1849, new_AGEMA_signal_1843}), .clk ( clk ), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .c ({new_AGEMA_signal_711, new_AGEMA_signal_710, new_AGEMA_signal_709, new_AGEMA_signal_708, sbe_inv_qmul_summul_n8}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_summul_U3 ( .a ({new_AGEMA_signal_667, new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_663, new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, sbe_inv_qmul_summul_n7}), .c ({new_AGEMA_signal_715, new_AGEMA_signal_714, new_AGEMA_signal_713, new_AGEMA_signal_712, sbe_inv_qmul_p_0_}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_summul_U2 ( .a ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1891, new_AGEMA_signal_1885, new_AGEMA_signal_1879, new_AGEMA_signal_1873}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({new_AGEMA_signal_663, new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, sbe_inv_qmul_summul_n7}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) sbe_inv_qmul_summul_U1 ( .a ({new_AGEMA_signal_595, new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1921, new_AGEMA_signal_1915, new_AGEMA_signal_1909, new_AGEMA_signal_1903}), .clk ( clk ), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_667, new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, sbe_inv_qmul_summul_n9}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m7_U2 ( .a ({new_AGEMA_signal_807, new_AGEMA_signal_806, new_AGEMA_signal_805, new_AGEMA_signal_804, sbe_sel_out_m7_n8}), .b ({new_AGEMA_signal_835, new_AGEMA_signal_834, new_AGEMA_signal_833, new_AGEMA_signal_832, O[7]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_775, new_AGEMA_signal_774, new_AGEMA_signal_773, new_AGEMA_signal_772, sbe_n15}), .a ({new_AGEMA_signal_787, new_AGEMA_signal_786, new_AGEMA_signal_785, new_AGEMA_signal_784, sbe_n19}), .c ({new_AGEMA_signal_807, new_AGEMA_signal_806, new_AGEMA_signal_805, new_AGEMA_signal_804, sbe_sel_out_m7_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m6_U2 ( .a ({new_AGEMA_signal_875, new_AGEMA_signal_874, new_AGEMA_signal_873, new_AGEMA_signal_872, sbe_sel_out_m6_n8}), .b ({new_AGEMA_signal_891, new_AGEMA_signal_890, new_AGEMA_signal_889, new_AGEMA_signal_888, O[6]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_851, new_AGEMA_signal_850, new_AGEMA_signal_849, new_AGEMA_signal_848, sbe_X[6]}), .a ({new_AGEMA_signal_783, new_AGEMA_signal_782, new_AGEMA_signal_781, new_AGEMA_signal_780, sbe_D_6_}), .c ({new_AGEMA_signal_875, new_AGEMA_signal_874, new_AGEMA_signal_873, new_AGEMA_signal_872, sbe_sel_out_m6_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m5_U2 ( .a ({new_AGEMA_signal_879, new_AGEMA_signal_878, new_AGEMA_signal_877, new_AGEMA_signal_876, sbe_sel_out_m5_n8}), .b ({new_AGEMA_signal_895, new_AGEMA_signal_894, new_AGEMA_signal_893, new_AGEMA_signal_892, O[5]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_855, new_AGEMA_signal_854, new_AGEMA_signal_853, new_AGEMA_signal_852, sbe_X[5]}), .a ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, new_AGEMA_signal_744, sbe_D_5_}), .c ({new_AGEMA_signal_879, new_AGEMA_signal_878, new_AGEMA_signal_877, new_AGEMA_signal_876, sbe_sel_out_m5_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m4_U2 ( .a ({new_AGEMA_signal_839, new_AGEMA_signal_838, new_AGEMA_signal_837, new_AGEMA_signal_836, sbe_sel_out_m4_n8}), .b ({new_AGEMA_signal_859, new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, O[4]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_779, new_AGEMA_signal_778, new_AGEMA_signal_777, new_AGEMA_signal_776, sbe_n14}), .a ({new_AGEMA_signal_799, new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, sbe_n20}), .c ({new_AGEMA_signal_839, new_AGEMA_signal_838, new_AGEMA_signal_837, new_AGEMA_signal_836, sbe_sel_out_m4_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m3_U2 ( .a ({new_AGEMA_signal_863, new_AGEMA_signal_862, new_AGEMA_signal_861, new_AGEMA_signal_860, sbe_sel_out_m3_n8}), .b ({new_AGEMA_signal_883, new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, O[3]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_823, new_AGEMA_signal_822, new_AGEMA_signal_821, new_AGEMA_signal_820, sbe_X[3]}), .a ({new_AGEMA_signal_827, new_AGEMA_signal_826, new_AGEMA_signal_825, new_AGEMA_signal_824, sbe_D_3_}), .c ({new_AGEMA_signal_863, new_AGEMA_signal_862, new_AGEMA_signal_861, new_AGEMA_signal_860, sbe_sel_out_m3_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m2_U2 ( .a ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, new_AGEMA_signal_864, sbe_sel_out_m2_n8}), .b ({new_AGEMA_signal_887, new_AGEMA_signal_886, new_AGEMA_signal_885, new_AGEMA_signal_884, O[2]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_815, new_AGEMA_signal_814, new_AGEMA_signal_813, new_AGEMA_signal_812, sbe_n16}), .a ({new_AGEMA_signal_831, new_AGEMA_signal_830, new_AGEMA_signal_829, new_AGEMA_signal_828, sbe_D_2_}), .c ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, new_AGEMA_signal_864, sbe_sel_out_m2_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m1_U2 ( .a ({new_AGEMA_signal_843, new_AGEMA_signal_842, new_AGEMA_signal_841, new_AGEMA_signal_840, sbe_sel_out_m1_n8}), .b ({new_AGEMA_signal_871, new_AGEMA_signal_870, new_AGEMA_signal_869, new_AGEMA_signal_868, O[1]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_771, new_AGEMA_signal_770, new_AGEMA_signal_769, new_AGEMA_signal_768, sbe_n18}), .a ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, new_AGEMA_signal_792, sbe_n17}), .c ({new_AGEMA_signal_843, new_AGEMA_signal_842, new_AGEMA_signal_841, new_AGEMA_signal_840, sbe_sel_out_m1_n8}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m0_U2 ( .a ({new_AGEMA_signal_811, new_AGEMA_signal_810, new_AGEMA_signal_809, new_AGEMA_signal_808, sbe_sel_out_m0_n8}), .b ({new_AGEMA_signal_847, new_AGEMA_signal_846, new_AGEMA_signal_845, new_AGEMA_signal_844, O[0]}) ) ;
    mux2_masked #(.security_order(4), .pipeline(1)) sbe_sel_out_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_743, new_AGEMA_signal_742, new_AGEMA_signal_741, new_AGEMA_signal_740, sbe_n1}), .a ({new_AGEMA_signal_791, new_AGEMA_signal_790, new_AGEMA_signal_789, new_AGEMA_signal_788, sbe_D_0_}), .c ({new_AGEMA_signal_811, new_AGEMA_signal_810, new_AGEMA_signal_809, new_AGEMA_signal_808, sbe_sel_out_m0_n8}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_835, new_AGEMA_signal_834, new_AGEMA_signal_833, new_AGEMA_signal_832, O[7]}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_891, new_AGEMA_signal_890, new_AGEMA_signal_889, new_AGEMA_signal_888, O[6]}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_895, new_AGEMA_signal_894, new_AGEMA_signal_893, new_AGEMA_signal_892, O[5]}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_859, new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, O[4]}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_883, new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, O[3]}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_887, new_AGEMA_signal_886, new_AGEMA_signal_885, new_AGEMA_signal_884, O[2]}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_871, new_AGEMA_signal_870, new_AGEMA_signal_869, new_AGEMA_signal_868, O[1]}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_847, new_AGEMA_signal_846, new_AGEMA_signal_845, new_AGEMA_signal_844, O[0]}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
